module SimpleDualPortRam(
  input         clock,
  input         reset,
  input  [8:0]  io_raddr,
  output [63:0] io_rdata,
  input  [8:0]  io_waddr,
  input         io_wen,
  input  [7:0]  io_wstrb,
  input  [63:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] bank_0 [0:511]; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_0_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_0_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_0_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_0_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_0_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_0_MPORT_mask; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_0_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  reg  bank_0_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_0_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_1 [0:511]; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_1_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_1_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_1_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_1_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_1_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_1_MPORT_mask; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_1_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  reg  bank_1_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_1_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_2 [0:511]; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_2_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_2_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_2_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_2_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_2_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_2_MPORT_mask; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_2_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  reg  bank_2_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_2_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_3 [0:511]; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_3_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_3_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_3_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_3_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_3_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_3_MPORT_mask; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_3_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  reg  bank_3_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_3_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_4 [0:511]; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_4_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_4_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_4_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_4_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_4_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_4_MPORT_mask; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_4_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  reg  bank_4_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_4_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_5 [0:511]; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_5_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_5_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_5_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_5_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_5_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_5_MPORT_mask; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_5_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  reg  bank_5_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_5_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_6 [0:511]; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_6_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_6_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_6_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_6_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_6_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_6_MPORT_mask; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_6_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  reg  bank_6_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_6_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_7 [0:511]; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_7_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_7_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_7_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [7:0] bank_7_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
  wire [8:0] bank_7_MPORT_addr; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_7_MPORT_mask; // @[SimpleDualPortRam.scala 71:29]
  wire  bank_7_MPORT_en; // @[SimpleDualPortRam.scala 71:29]
  reg  bank_7_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_7_io_rdata_MPORT_addr_pipe_0;
  wire  _T_2 = |io_wstrb | ~io_wen; // @[SimpleDualPortRam.scala 67:20]
  wire [31:0] io_rdata_lo = {bank_3_io_rdata_MPORT_data,bank_2_io_rdata_MPORT_data,bank_1_io_rdata_MPORT_data,
    bank_0_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 73:44]
  wire [31:0] io_rdata_hi = {bank_7_io_rdata_MPORT_data,bank_6_io_rdata_MPORT_data,bank_5_io_rdata_MPORT_data,
    bank_4_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 73:44]
  assign bank_0_io_rdata_MPORT_en = bank_0_io_rdata_MPORT_en_pipe_0;
  assign bank_0_io_rdata_MPORT_addr = bank_0_io_rdata_MPORT_addr_pipe_0;
  assign bank_0_io_rdata_MPORT_data = bank_0[bank_0_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 71:29]
  assign bank_0_MPORT_data = io_wdata[7:0];
  assign bank_0_MPORT_addr = io_waddr;
  assign bank_0_MPORT_mask = io_wstrb[0];
  assign bank_0_MPORT_en = io_wen;
  assign bank_1_io_rdata_MPORT_en = bank_1_io_rdata_MPORT_en_pipe_0;
  assign bank_1_io_rdata_MPORT_addr = bank_1_io_rdata_MPORT_addr_pipe_0;
  assign bank_1_io_rdata_MPORT_data = bank_1[bank_1_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 71:29]
  assign bank_1_MPORT_data = io_wdata[15:8];
  assign bank_1_MPORT_addr = io_waddr;
  assign bank_1_MPORT_mask = io_wstrb[1];
  assign bank_1_MPORT_en = io_wen;
  assign bank_2_io_rdata_MPORT_en = bank_2_io_rdata_MPORT_en_pipe_0;
  assign bank_2_io_rdata_MPORT_addr = bank_2_io_rdata_MPORT_addr_pipe_0;
  assign bank_2_io_rdata_MPORT_data = bank_2[bank_2_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 71:29]
  assign bank_2_MPORT_data = io_wdata[23:16];
  assign bank_2_MPORT_addr = io_waddr;
  assign bank_2_MPORT_mask = io_wstrb[2];
  assign bank_2_MPORT_en = io_wen;
  assign bank_3_io_rdata_MPORT_en = bank_3_io_rdata_MPORT_en_pipe_0;
  assign bank_3_io_rdata_MPORT_addr = bank_3_io_rdata_MPORT_addr_pipe_0;
  assign bank_3_io_rdata_MPORT_data = bank_3[bank_3_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 71:29]
  assign bank_3_MPORT_data = io_wdata[31:24];
  assign bank_3_MPORT_addr = io_waddr;
  assign bank_3_MPORT_mask = io_wstrb[3];
  assign bank_3_MPORT_en = io_wen;
  assign bank_4_io_rdata_MPORT_en = bank_4_io_rdata_MPORT_en_pipe_0;
  assign bank_4_io_rdata_MPORT_addr = bank_4_io_rdata_MPORT_addr_pipe_0;
  assign bank_4_io_rdata_MPORT_data = bank_4[bank_4_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 71:29]
  assign bank_4_MPORT_data = io_wdata[39:32];
  assign bank_4_MPORT_addr = io_waddr;
  assign bank_4_MPORT_mask = io_wstrb[4];
  assign bank_4_MPORT_en = io_wen;
  assign bank_5_io_rdata_MPORT_en = bank_5_io_rdata_MPORT_en_pipe_0;
  assign bank_5_io_rdata_MPORT_addr = bank_5_io_rdata_MPORT_addr_pipe_0;
  assign bank_5_io_rdata_MPORT_data = bank_5[bank_5_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 71:29]
  assign bank_5_MPORT_data = io_wdata[47:40];
  assign bank_5_MPORT_addr = io_waddr;
  assign bank_5_MPORT_mask = io_wstrb[5];
  assign bank_5_MPORT_en = io_wen;
  assign bank_6_io_rdata_MPORT_en = bank_6_io_rdata_MPORT_en_pipe_0;
  assign bank_6_io_rdata_MPORT_addr = bank_6_io_rdata_MPORT_addr_pipe_0;
  assign bank_6_io_rdata_MPORT_data = bank_6[bank_6_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 71:29]
  assign bank_6_MPORT_data = io_wdata[55:48];
  assign bank_6_MPORT_addr = io_waddr;
  assign bank_6_MPORT_mask = io_wstrb[6];
  assign bank_6_MPORT_en = io_wen;
  assign bank_7_io_rdata_MPORT_en = bank_7_io_rdata_MPORT_en_pipe_0;
  assign bank_7_io_rdata_MPORT_addr = bank_7_io_rdata_MPORT_addr_pipe_0;
  assign bank_7_io_rdata_MPORT_data = bank_7[bank_7_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 71:29]
  assign bank_7_MPORT_data = io_wdata[63:56];
  assign bank_7_MPORT_addr = io_waddr;
  assign bank_7_MPORT_mask = io_wstrb[7];
  assign bank_7_MPORT_en = io_wen;
  assign io_rdata = {io_rdata_hi,io_rdata_lo}; // @[SimpleDualPortRam.scala 73:44]
  always @(posedge clock) begin
    if (bank_0_MPORT_en & bank_0_MPORT_mask) begin
      bank_0[bank_0_MPORT_addr] <= bank_0_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
    end
    bank_0_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_0_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_1_MPORT_en & bank_1_MPORT_mask) begin
      bank_1[bank_1_MPORT_addr] <= bank_1_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
    end
    bank_1_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_1_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_2_MPORT_en & bank_2_MPORT_mask) begin
      bank_2[bank_2_MPORT_addr] <= bank_2_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
    end
    bank_2_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_2_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_3_MPORT_en & bank_3_MPORT_mask) begin
      bank_3[bank_3_MPORT_addr] <= bank_3_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
    end
    bank_3_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_3_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_4_MPORT_en & bank_4_MPORT_mask) begin
      bank_4[bank_4_MPORT_addr] <= bank_4_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
    end
    bank_4_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_4_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_5_MPORT_en & bank_5_MPORT_mask) begin
      bank_5[bank_5_MPORT_addr] <= bank_5_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
    end
    bank_5_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_5_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_6_MPORT_en & bank_6_MPORT_mask) begin
      bank_6[bank_6_MPORT_addr] <= bank_6_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
    end
    bank_6_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_6_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_7_MPORT_en & bank_7_MPORT_mask) begin
      bank_7[bank_7_MPORT_addr] <= bank_7_MPORT_data; // @[SimpleDualPortRam.scala 71:29]
    end
    bank_7_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_7_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed: when write port enable is high, write vector cannot be all 0\n    at SimpleDualPortRam.scala:66 assert(\n"
            ); // @[SimpleDualPortRam.scala 66:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fatal; // @[SimpleDualPortRam.scala 66:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_0[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_1[initvar] = _RAND_3[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_2[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_3[initvar] = _RAND_9[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_4[initvar] = _RAND_12[7:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_5[initvar] = _RAND_15[7:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_6[initvar] = _RAND_18[7:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_7[initvar] = _RAND_21[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bank_0_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bank_0_io_rdata_MPORT_addr_pipe_0 = _RAND_2[8:0];
  _RAND_4 = {1{`RANDOM}};
  bank_1_io_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  bank_1_io_rdata_MPORT_addr_pipe_0 = _RAND_5[8:0];
  _RAND_7 = {1{`RANDOM}};
  bank_2_io_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  bank_2_io_rdata_MPORT_addr_pipe_0 = _RAND_8[8:0];
  _RAND_10 = {1{`RANDOM}};
  bank_3_io_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  bank_3_io_rdata_MPORT_addr_pipe_0 = _RAND_11[8:0];
  _RAND_13 = {1{`RANDOM}};
  bank_4_io_rdata_MPORT_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  bank_4_io_rdata_MPORT_addr_pipe_0 = _RAND_14[8:0];
  _RAND_16 = {1{`RANDOM}};
  bank_5_io_rdata_MPORT_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  bank_5_io_rdata_MPORT_addr_pipe_0 = _RAND_17[8:0];
  _RAND_19 = {1{`RANDOM}};
  bank_6_io_rdata_MPORT_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  bank_6_io_rdata_MPORT_addr_pipe_0 = _RAND_20[8:0];
  _RAND_22 = {1{`RANDOM}};
  bank_7_io_rdata_MPORT_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  bank_7_io_rdata_MPORT_addr_pipe_0 = _RAND_23[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Bank(
  input         clock,
  input         reset,
  input  [8:0]  io_way_0_r_addr,
  output [63:0] io_way_0_r_data,
  input  [8:0]  io_way_0_w_addr,
  input  [7:0]  io_way_0_w_en,
  input  [63:0] io_way_0_w_data,
  input  [8:0]  io_way_1_r_addr,
  output [63:0] io_way_1_r_data,
  input  [8:0]  io_way_1_w_addr,
  input  [7:0]  io_way_1_w_en,
  input  [63:0] io_way_1_w_data
);
  wire  bank0_clock; // @[Bank.scala 26:22]
  wire  bank0_reset; // @[Bank.scala 26:22]
  wire [8:0] bank0_io_raddr; // @[Bank.scala 26:22]
  wire [63:0] bank0_io_rdata; // @[Bank.scala 26:22]
  wire [8:0] bank0_io_waddr; // @[Bank.scala 26:22]
  wire  bank0_io_wen; // @[Bank.scala 26:22]
  wire [7:0] bank0_io_wstrb; // @[Bank.scala 26:22]
  wire [63:0] bank0_io_wdata; // @[Bank.scala 26:22]
  wire  bank1_clock; // @[Bank.scala 26:22]
  wire  bank1_reset; // @[Bank.scala 26:22]
  wire [8:0] bank1_io_raddr; // @[Bank.scala 26:22]
  wire [63:0] bank1_io_rdata; // @[Bank.scala 26:22]
  wire [8:0] bank1_io_waddr; // @[Bank.scala 26:22]
  wire  bank1_io_wen; // @[Bank.scala 26:22]
  wire [7:0] bank1_io_wstrb; // @[Bank.scala 26:22]
  wire [63:0] bank1_io_wdata; // @[Bank.scala 26:22]
  SimpleDualPortRam bank0 ( // @[Bank.scala 26:22]
    .clock(bank0_clock),
    .reset(bank0_reset),
    .io_raddr(bank0_io_raddr),
    .io_rdata(bank0_io_rdata),
    .io_waddr(bank0_io_waddr),
    .io_wen(bank0_io_wen),
    .io_wstrb(bank0_io_wstrb),
    .io_wdata(bank0_io_wdata)
  );
  SimpleDualPortRam bank1 ( // @[Bank.scala 26:22]
    .clock(bank1_clock),
    .reset(bank1_reset),
    .io_raddr(bank1_io_raddr),
    .io_rdata(bank1_io_rdata),
    .io_waddr(bank1_io_waddr),
    .io_wen(bank1_io_wen),
    .io_wstrb(bank1_io_wstrb),
    .io_wdata(bank1_io_wdata)
  );
  assign io_way_0_r_data = bank0_io_rdata; // @[Bank.scala 32:22]
  assign io_way_1_r_data = bank1_io_rdata; // @[Bank.scala 32:22]
  assign bank0_clock = clock;
  assign bank0_reset = reset;
  assign bank0_io_raddr = io_way_0_r_addr; // @[Bank.scala 31:22]
  assign bank0_io_waddr = io_way_0_w_addr; // @[Bank.scala 36:19]
  assign bank0_io_wen = |io_way_0_w_en; // @[Bank.scala 35:37]
  assign bank0_io_wstrb = io_way_0_w_en; // @[Bank.scala 38:19]
  assign bank0_io_wdata = io_way_0_w_data; // @[Bank.scala 37:19]
  assign bank1_clock = clock;
  assign bank1_reset = reset;
  assign bank1_io_raddr = io_way_1_r_addr; // @[Bank.scala 31:22]
  assign bank1_io_waddr = io_way_1_w_addr; // @[Bank.scala 36:19]
  assign bank1_io_wen = |io_way_1_w_en; // @[Bank.scala 35:37]
  assign bank1_io_wstrb = io_way_1_w_en; // @[Bank.scala 38:19]
  assign bank1_io_wdata = io_way_1_w_data; // @[Bank.scala 37:19]
endmodule
module SimpleDualPortRam_2(
  input         clock,
  input         reset,
  input  [8:0]  io_raddr,
  output [19:0] io_rdata,
  input  [8:0]  io_waddr,
  input         io_wen,
  input         io_wstrb,
  input  [19:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] bank [0:511]; // @[SimpleDualPortRam.scala 81:29]
  wire  bank_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 81:29]
  wire [8:0] bank_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 81:29]
  wire [19:0] bank_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 81:29]
  wire [19:0] bank_MPORT_data; // @[SimpleDualPortRam.scala 81:29]
  wire [8:0] bank_MPORT_addr; // @[SimpleDualPortRam.scala 81:29]
  wire  bank_MPORT_mask; // @[SimpleDualPortRam.scala 81:29]
  wire  bank_MPORT_en; // @[SimpleDualPortRam.scala 81:29]
  reg  bank_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_io_rdata_MPORT_addr_pipe_0;
  wire  _T_2 = |io_wstrb | ~io_wen; // @[SimpleDualPortRam.scala 67:20]
  wire [31:0] _GEN_7 = {{12'd0}, bank_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 83:20 84:18 86:18]
  assign bank_io_rdata_MPORT_en = bank_io_rdata_MPORT_en_pipe_0;
  assign bank_io_rdata_MPORT_addr = bank_io_rdata_MPORT_addr_pipe_0;
  assign bank_io_rdata_MPORT_data = bank[bank_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 81:29]
  assign bank_MPORT_data = io_wdata;
  assign bank_MPORT_addr = io_waddr;
  assign bank_MPORT_mask = 1'h1;
  assign bank_MPORT_en = io_wen;
  assign io_rdata = _GEN_7[19:0];
  always @(posedge clock) begin
    if (bank_MPORT_en & bank_MPORT_mask) begin
      bank[bank_MPORT_addr] <= bank_MPORT_data; // @[SimpleDualPortRam.scala 81:29]
    end
    bank_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed: when write port enable is high, write vector cannot be all 0\n    at SimpleDualPortRam.scala:66 assert(\n"
            ); // @[SimpleDualPortRam.scala 66:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fatal; // @[SimpleDualPortRam.scala 66:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bank_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bank_io_rdata_MPORT_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Tag(
  input         clock,
  input         reset,
  input  [8:0]  io_way_0_r_addr,
  output [16:0] io_way_0_r_data,
  input  [8:0]  io_way_0_w_addr,
  input         io_way_0_w_en,
  input  [16:0] io_way_0_w_data,
  input  [8:0]  io_way_1_r_addr,
  output [16:0] io_way_1_r_data,
  input  [8:0]  io_way_1_w_addr,
  input         io_way_1_w_en,
  input  [16:0] io_way_1_w_data
);
  wire  tag_0_clock; // @[Tag.scala 23:21]
  wire  tag_0_reset; // @[Tag.scala 23:21]
  wire [8:0] tag_0_io_raddr; // @[Tag.scala 23:21]
  wire [19:0] tag_0_io_rdata; // @[Tag.scala 23:21]
  wire [8:0] tag_0_io_waddr; // @[Tag.scala 23:21]
  wire  tag_0_io_wen; // @[Tag.scala 23:21]
  wire  tag_0_io_wstrb; // @[Tag.scala 23:21]
  wire [19:0] tag_0_io_wdata; // @[Tag.scala 23:21]
  wire  tag_1_clock; // @[Tag.scala 23:21]
  wire  tag_1_reset; // @[Tag.scala 23:21]
  wire [8:0] tag_1_io_raddr; // @[Tag.scala 23:21]
  wire [19:0] tag_1_io_rdata; // @[Tag.scala 23:21]
  wire [8:0] tag_1_io_waddr; // @[Tag.scala 23:21]
  wire  tag_1_io_wen; // @[Tag.scala 23:21]
  wire  tag_1_io_wstrb; // @[Tag.scala 23:21]
  wire [19:0] tag_1_io_wdata; // @[Tag.scala 23:21]
  SimpleDualPortRam_2 tag_0 ( // @[Tag.scala 23:21]
    .clock(tag_0_clock),
    .reset(tag_0_reset),
    .io_raddr(tag_0_io_raddr),
    .io_rdata(tag_0_io_rdata),
    .io_waddr(tag_0_io_waddr),
    .io_wen(tag_0_io_wen),
    .io_wstrb(tag_0_io_wstrb),
    .io_wdata(tag_0_io_wdata)
  );
  SimpleDualPortRam_2 tag_1 ( // @[Tag.scala 23:21]
    .clock(tag_1_clock),
    .reset(tag_1_reset),
    .io_raddr(tag_1_io_raddr),
    .io_rdata(tag_1_io_rdata),
    .io_waddr(tag_1_io_waddr),
    .io_wen(tag_1_io_wen),
    .io_wstrb(tag_1_io_wstrb),
    .io_wdata(tag_1_io_wdata)
  );
  assign io_way_0_r_data = tag_0_io_rdata[16:0]; // @[Tag.scala 29:22]
  assign io_way_1_r_data = tag_1_io_rdata[16:0]; // @[Tag.scala 29:22]
  assign tag_0_clock = clock;
  assign tag_0_reset = reset;
  assign tag_0_io_raddr = io_way_0_r_addr; // @[Tag.scala 28:22]
  assign tag_0_io_waddr = io_way_0_w_addr; // @[Tag.scala 31:18]
  assign tag_0_io_wen = io_way_0_w_en; // @[Tag.scala 32:18]
  assign tag_0_io_wstrb = io_way_0_w_en; // @[Tag.scala 34:18]
  assign tag_0_io_wdata = {{3'd0}, io_way_0_w_data}; // @[Tag.scala 33:18]
  assign tag_1_clock = clock;
  assign tag_1_reset = reset;
  assign tag_1_io_raddr = io_way_1_r_addr; // @[Tag.scala 28:22]
  assign tag_1_io_waddr = io_way_1_w_addr; // @[Tag.scala 31:18]
  assign tag_1_io_wen = io_way_1_w_en; // @[Tag.scala 32:18]
  assign tag_1_io_wstrb = io_way_1_w_en; // @[Tag.scala 34:18]
  assign tag_1_io_wdata = {{3'd0}, io_way_1_w_data}; // @[Tag.scala 33:18]
endmodule
module ICache(
  input         clock,
  input         reset,
  input         io_cpu_req,
  input  [31:0] io_cpu_addr_0,
  input  [31:0] io_cpu_addr_1,
  output [31:0] io_cpu_inst_0,
  output [31:0] io_cpu_inst_1,
  output        io_cpu_inst_valid_0,
  output        io_cpu_inst_valid_1,
  input         io_cpu_cpu_stall,
  output        io_cpu_icache_stall,
  output        io_cpu_tlb1_refill,
  output        io_cpu_tlb1_invalid,
  output [18:0] io_cpu_tlb2_vpn,
  input         io_cpu_tlb2_found,
  input         io_cpu_tlb2_entry_G,
  input         io_cpu_tlb2_entry_V0,
  input         io_cpu_tlb2_entry_V1,
  input         io_cpu_tlb2_entry_D0,
  input         io_cpu_tlb2_entry_D1,
  input         io_cpu_tlb2_entry_C0,
  input         io_cpu_tlb2_entry_C1,
  input  [19:0] io_cpu_tlb2_entry_PFN0,
  input  [19:0] io_cpu_tlb2_entry_PFN1,
  input  [18:0] io_cpu_tlb2_entry_VPN2,
  input  [7:0]  io_cpu_tlb2_entry_ASID,
  input         io_cpu_fence_value,
  input  [31:0] io_cpu_fence_addr,
  input         io_cpu_fence_tlb,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output [7:0]  io_axi_ar_bits_len,
  output [2:0]  io_axi_ar_bits_size,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [31:0] io_axi_r_bits_data,
  input         io_axi_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
`endif // RANDOMIZE_REG_INIT
  wire  bank_ram_clock; // @[ICache.scala 112:24]
  wire  bank_ram_reset; // @[ICache.scala 112:24]
  wire [8:0] bank_ram_io_way_0_r_addr; // @[ICache.scala 112:24]
  wire [63:0] bank_ram_io_way_0_r_data; // @[ICache.scala 112:24]
  wire [8:0] bank_ram_io_way_0_w_addr; // @[ICache.scala 112:24]
  wire [7:0] bank_ram_io_way_0_w_en; // @[ICache.scala 112:24]
  wire [63:0] bank_ram_io_way_0_w_data; // @[ICache.scala 112:24]
  wire [8:0] bank_ram_io_way_1_r_addr; // @[ICache.scala 112:24]
  wire [63:0] bank_ram_io_way_1_r_data; // @[ICache.scala 112:24]
  wire [8:0] bank_ram_io_way_1_w_addr; // @[ICache.scala 112:24]
  wire [7:0] bank_ram_io_way_1_w_en; // @[ICache.scala 112:24]
  wire [63:0] bank_ram_io_way_1_w_data; // @[ICache.scala 112:24]
  wire  tag_ram_clock; // @[ICache.scala 125:23]
  wire  tag_ram_reset; // @[ICache.scala 125:23]
  wire [8:0] tag_ram_io_way_0_r_addr; // @[ICache.scala 125:23]
  wire [16:0] tag_ram_io_way_0_r_data; // @[ICache.scala 125:23]
  wire [8:0] tag_ram_io_way_0_w_addr; // @[ICache.scala 125:23]
  wire  tag_ram_io_way_0_w_en; // @[ICache.scala 125:23]
  wire [16:0] tag_ram_io_way_0_w_data; // @[ICache.scala 125:23]
  wire [8:0] tag_ram_io_way_1_r_addr; // @[ICache.scala 125:23]
  wire [16:0] tag_ram_io_way_1_r_data; // @[ICache.scala 125:23]
  wire [8:0] tag_ram_io_way_1_w_addr; // @[ICache.scala 125:23]
  wire  tag_ram_io_way_1_w_en; // @[ICache.scala 125:23]
  wire [16:0] tag_ram_io_way_1_w_data; // @[ICache.scala 125:23]
  reg  meta_0_valid_0; // @[ICache.scala 34:21]
  reg  meta_0_valid_1; // @[ICache.scala 34:21]
  reg  meta_0_lru; // @[ICache.scala 34:21]
  reg  meta_1_valid_0; // @[ICache.scala 34:21]
  reg  meta_1_valid_1; // @[ICache.scala 34:21]
  reg  meta_1_lru; // @[ICache.scala 34:21]
  reg  meta_2_valid_0; // @[ICache.scala 34:21]
  reg  meta_2_valid_1; // @[ICache.scala 34:21]
  reg  meta_2_lru; // @[ICache.scala 34:21]
  reg  meta_3_valid_0; // @[ICache.scala 34:21]
  reg  meta_3_valid_1; // @[ICache.scala 34:21]
  reg  meta_3_lru; // @[ICache.scala 34:21]
  reg  meta_4_valid_0; // @[ICache.scala 34:21]
  reg  meta_4_valid_1; // @[ICache.scala 34:21]
  reg  meta_4_lru; // @[ICache.scala 34:21]
  reg  meta_5_valid_0; // @[ICache.scala 34:21]
  reg  meta_5_valid_1; // @[ICache.scala 34:21]
  reg  meta_5_lru; // @[ICache.scala 34:21]
  reg  meta_6_valid_0; // @[ICache.scala 34:21]
  reg  meta_6_valid_1; // @[ICache.scala 34:21]
  reg  meta_6_lru; // @[ICache.scala 34:21]
  reg  meta_7_valid_0; // @[ICache.scala 34:21]
  reg  meta_7_valid_1; // @[ICache.scala 34:21]
  reg  meta_7_lru; // @[ICache.scala 34:21]
  reg  meta_8_valid_0; // @[ICache.scala 34:21]
  reg  meta_8_valid_1; // @[ICache.scala 34:21]
  reg  meta_8_lru; // @[ICache.scala 34:21]
  reg  meta_9_valid_0; // @[ICache.scala 34:21]
  reg  meta_9_valid_1; // @[ICache.scala 34:21]
  reg  meta_9_lru; // @[ICache.scala 34:21]
  reg  meta_10_valid_0; // @[ICache.scala 34:21]
  reg  meta_10_valid_1; // @[ICache.scala 34:21]
  reg  meta_10_lru; // @[ICache.scala 34:21]
  reg  meta_11_valid_0; // @[ICache.scala 34:21]
  reg  meta_11_valid_1; // @[ICache.scala 34:21]
  reg  meta_11_lru; // @[ICache.scala 34:21]
  reg  meta_12_valid_0; // @[ICache.scala 34:21]
  reg  meta_12_valid_1; // @[ICache.scala 34:21]
  reg  meta_12_lru; // @[ICache.scala 34:21]
  reg  meta_13_valid_0; // @[ICache.scala 34:21]
  reg  meta_13_valid_1; // @[ICache.scala 34:21]
  reg  meta_13_lru; // @[ICache.scala 34:21]
  reg  meta_14_valid_0; // @[ICache.scala 34:21]
  reg  meta_14_valid_1; // @[ICache.scala 34:21]
  reg  meta_14_lru; // @[ICache.scala 34:21]
  reg  meta_15_valid_0; // @[ICache.scala 34:21]
  reg  meta_15_valid_1; // @[ICache.scala 34:21]
  reg  meta_15_lru; // @[ICache.scala 34:21]
  reg  meta_16_valid_0; // @[ICache.scala 34:21]
  reg  meta_16_valid_1; // @[ICache.scala 34:21]
  reg  meta_16_lru; // @[ICache.scala 34:21]
  reg  meta_17_valid_0; // @[ICache.scala 34:21]
  reg  meta_17_valid_1; // @[ICache.scala 34:21]
  reg  meta_17_lru; // @[ICache.scala 34:21]
  reg  meta_18_valid_0; // @[ICache.scala 34:21]
  reg  meta_18_valid_1; // @[ICache.scala 34:21]
  reg  meta_18_lru; // @[ICache.scala 34:21]
  reg  meta_19_valid_0; // @[ICache.scala 34:21]
  reg  meta_19_valid_1; // @[ICache.scala 34:21]
  reg  meta_19_lru; // @[ICache.scala 34:21]
  reg  meta_20_valid_0; // @[ICache.scala 34:21]
  reg  meta_20_valid_1; // @[ICache.scala 34:21]
  reg  meta_20_lru; // @[ICache.scala 34:21]
  reg  meta_21_valid_0; // @[ICache.scala 34:21]
  reg  meta_21_valid_1; // @[ICache.scala 34:21]
  reg  meta_21_lru; // @[ICache.scala 34:21]
  reg  meta_22_valid_0; // @[ICache.scala 34:21]
  reg  meta_22_valid_1; // @[ICache.scala 34:21]
  reg  meta_22_lru; // @[ICache.scala 34:21]
  reg  meta_23_valid_0; // @[ICache.scala 34:21]
  reg  meta_23_valid_1; // @[ICache.scala 34:21]
  reg  meta_23_lru; // @[ICache.scala 34:21]
  reg  meta_24_valid_0; // @[ICache.scala 34:21]
  reg  meta_24_valid_1; // @[ICache.scala 34:21]
  reg  meta_24_lru; // @[ICache.scala 34:21]
  reg  meta_25_valid_0; // @[ICache.scala 34:21]
  reg  meta_25_valid_1; // @[ICache.scala 34:21]
  reg  meta_25_lru; // @[ICache.scala 34:21]
  reg  meta_26_valid_0; // @[ICache.scala 34:21]
  reg  meta_26_valid_1; // @[ICache.scala 34:21]
  reg  meta_26_lru; // @[ICache.scala 34:21]
  reg  meta_27_valid_0; // @[ICache.scala 34:21]
  reg  meta_27_valid_1; // @[ICache.scala 34:21]
  reg  meta_27_lru; // @[ICache.scala 34:21]
  reg  meta_28_valid_0; // @[ICache.scala 34:21]
  reg  meta_28_valid_1; // @[ICache.scala 34:21]
  reg  meta_28_lru; // @[ICache.scala 34:21]
  reg  meta_29_valid_0; // @[ICache.scala 34:21]
  reg  meta_29_valid_1; // @[ICache.scala 34:21]
  reg  meta_29_lru; // @[ICache.scala 34:21]
  reg  meta_30_valid_0; // @[ICache.scala 34:21]
  reg  meta_30_valid_1; // @[ICache.scala 34:21]
  reg  meta_30_lru; // @[ICache.scala 34:21]
  reg  meta_31_valid_0; // @[ICache.scala 34:21]
  reg  meta_31_valid_1; // @[ICache.scala 34:21]
  reg  meta_31_lru; // @[ICache.scala 34:21]
  reg  meta_32_valid_0; // @[ICache.scala 34:21]
  reg  meta_32_valid_1; // @[ICache.scala 34:21]
  reg  meta_32_lru; // @[ICache.scala 34:21]
  reg  meta_33_valid_0; // @[ICache.scala 34:21]
  reg  meta_33_valid_1; // @[ICache.scala 34:21]
  reg  meta_33_lru; // @[ICache.scala 34:21]
  reg  meta_34_valid_0; // @[ICache.scala 34:21]
  reg  meta_34_valid_1; // @[ICache.scala 34:21]
  reg  meta_34_lru; // @[ICache.scala 34:21]
  reg  meta_35_valid_0; // @[ICache.scala 34:21]
  reg  meta_35_valid_1; // @[ICache.scala 34:21]
  reg  meta_35_lru; // @[ICache.scala 34:21]
  reg  meta_36_valid_0; // @[ICache.scala 34:21]
  reg  meta_36_valid_1; // @[ICache.scala 34:21]
  reg  meta_36_lru; // @[ICache.scala 34:21]
  reg  meta_37_valid_0; // @[ICache.scala 34:21]
  reg  meta_37_valid_1; // @[ICache.scala 34:21]
  reg  meta_37_lru; // @[ICache.scala 34:21]
  reg  meta_38_valid_0; // @[ICache.scala 34:21]
  reg  meta_38_valid_1; // @[ICache.scala 34:21]
  reg  meta_38_lru; // @[ICache.scala 34:21]
  reg  meta_39_valid_0; // @[ICache.scala 34:21]
  reg  meta_39_valid_1; // @[ICache.scala 34:21]
  reg  meta_39_lru; // @[ICache.scala 34:21]
  reg  meta_40_valid_0; // @[ICache.scala 34:21]
  reg  meta_40_valid_1; // @[ICache.scala 34:21]
  reg  meta_40_lru; // @[ICache.scala 34:21]
  reg  meta_41_valid_0; // @[ICache.scala 34:21]
  reg  meta_41_valid_1; // @[ICache.scala 34:21]
  reg  meta_41_lru; // @[ICache.scala 34:21]
  reg  meta_42_valid_0; // @[ICache.scala 34:21]
  reg  meta_42_valid_1; // @[ICache.scala 34:21]
  reg  meta_42_lru; // @[ICache.scala 34:21]
  reg  meta_43_valid_0; // @[ICache.scala 34:21]
  reg  meta_43_valid_1; // @[ICache.scala 34:21]
  reg  meta_43_lru; // @[ICache.scala 34:21]
  reg  meta_44_valid_0; // @[ICache.scala 34:21]
  reg  meta_44_valid_1; // @[ICache.scala 34:21]
  reg  meta_44_lru; // @[ICache.scala 34:21]
  reg  meta_45_valid_0; // @[ICache.scala 34:21]
  reg  meta_45_valid_1; // @[ICache.scala 34:21]
  reg  meta_45_lru; // @[ICache.scala 34:21]
  reg  meta_46_valid_0; // @[ICache.scala 34:21]
  reg  meta_46_valid_1; // @[ICache.scala 34:21]
  reg  meta_46_lru; // @[ICache.scala 34:21]
  reg  meta_47_valid_0; // @[ICache.scala 34:21]
  reg  meta_47_valid_1; // @[ICache.scala 34:21]
  reg  meta_47_lru; // @[ICache.scala 34:21]
  reg  meta_48_valid_0; // @[ICache.scala 34:21]
  reg  meta_48_valid_1; // @[ICache.scala 34:21]
  reg  meta_48_lru; // @[ICache.scala 34:21]
  reg  meta_49_valid_0; // @[ICache.scala 34:21]
  reg  meta_49_valid_1; // @[ICache.scala 34:21]
  reg  meta_49_lru; // @[ICache.scala 34:21]
  reg  meta_50_valid_0; // @[ICache.scala 34:21]
  reg  meta_50_valid_1; // @[ICache.scala 34:21]
  reg  meta_50_lru; // @[ICache.scala 34:21]
  reg  meta_51_valid_0; // @[ICache.scala 34:21]
  reg  meta_51_valid_1; // @[ICache.scala 34:21]
  reg  meta_51_lru; // @[ICache.scala 34:21]
  reg  meta_52_valid_0; // @[ICache.scala 34:21]
  reg  meta_52_valid_1; // @[ICache.scala 34:21]
  reg  meta_52_lru; // @[ICache.scala 34:21]
  reg  meta_53_valid_0; // @[ICache.scala 34:21]
  reg  meta_53_valid_1; // @[ICache.scala 34:21]
  reg  meta_53_lru; // @[ICache.scala 34:21]
  reg  meta_54_valid_0; // @[ICache.scala 34:21]
  reg  meta_54_valid_1; // @[ICache.scala 34:21]
  reg  meta_54_lru; // @[ICache.scala 34:21]
  reg  meta_55_valid_0; // @[ICache.scala 34:21]
  reg  meta_55_valid_1; // @[ICache.scala 34:21]
  reg  meta_55_lru; // @[ICache.scala 34:21]
  reg  meta_56_valid_0; // @[ICache.scala 34:21]
  reg  meta_56_valid_1; // @[ICache.scala 34:21]
  reg  meta_56_lru; // @[ICache.scala 34:21]
  reg  meta_57_valid_0; // @[ICache.scala 34:21]
  reg  meta_57_valid_1; // @[ICache.scala 34:21]
  reg  meta_57_lru; // @[ICache.scala 34:21]
  reg  meta_58_valid_0; // @[ICache.scala 34:21]
  reg  meta_58_valid_1; // @[ICache.scala 34:21]
  reg  meta_58_lru; // @[ICache.scala 34:21]
  reg  meta_59_valid_0; // @[ICache.scala 34:21]
  reg  meta_59_valid_1; // @[ICache.scala 34:21]
  reg  meta_59_lru; // @[ICache.scala 34:21]
  reg  meta_60_valid_0; // @[ICache.scala 34:21]
  reg  meta_60_valid_1; // @[ICache.scala 34:21]
  reg  meta_60_lru; // @[ICache.scala 34:21]
  reg  meta_61_valid_0; // @[ICache.scala 34:21]
  reg  meta_61_valid_1; // @[ICache.scala 34:21]
  reg  meta_61_lru; // @[ICache.scala 34:21]
  reg  meta_62_valid_0; // @[ICache.scala 34:21]
  reg  meta_62_valid_1; // @[ICache.scala 34:21]
  reg  meta_62_lru; // @[ICache.scala 34:21]
  reg  meta_63_valid_0; // @[ICache.scala 34:21]
  reg  meta_63_valid_1; // @[ICache.scala 34:21]
  reg  meta_63_lru; // @[ICache.scala 34:21]
  reg  meta_64_valid_0; // @[ICache.scala 34:21]
  reg  meta_64_valid_1; // @[ICache.scala 34:21]
  reg  meta_64_lru; // @[ICache.scala 34:21]
  reg  meta_65_valid_0; // @[ICache.scala 34:21]
  reg  meta_65_valid_1; // @[ICache.scala 34:21]
  reg  meta_65_lru; // @[ICache.scala 34:21]
  reg  meta_66_valid_0; // @[ICache.scala 34:21]
  reg  meta_66_valid_1; // @[ICache.scala 34:21]
  reg  meta_66_lru; // @[ICache.scala 34:21]
  reg  meta_67_valid_0; // @[ICache.scala 34:21]
  reg  meta_67_valid_1; // @[ICache.scala 34:21]
  reg  meta_67_lru; // @[ICache.scala 34:21]
  reg  meta_68_valid_0; // @[ICache.scala 34:21]
  reg  meta_68_valid_1; // @[ICache.scala 34:21]
  reg  meta_68_lru; // @[ICache.scala 34:21]
  reg  meta_69_valid_0; // @[ICache.scala 34:21]
  reg  meta_69_valid_1; // @[ICache.scala 34:21]
  reg  meta_69_lru; // @[ICache.scala 34:21]
  reg  meta_70_valid_0; // @[ICache.scala 34:21]
  reg  meta_70_valid_1; // @[ICache.scala 34:21]
  reg  meta_70_lru; // @[ICache.scala 34:21]
  reg  meta_71_valid_0; // @[ICache.scala 34:21]
  reg  meta_71_valid_1; // @[ICache.scala 34:21]
  reg  meta_71_lru; // @[ICache.scala 34:21]
  reg  meta_72_valid_0; // @[ICache.scala 34:21]
  reg  meta_72_valid_1; // @[ICache.scala 34:21]
  reg  meta_72_lru; // @[ICache.scala 34:21]
  reg  meta_73_valid_0; // @[ICache.scala 34:21]
  reg  meta_73_valid_1; // @[ICache.scala 34:21]
  reg  meta_73_lru; // @[ICache.scala 34:21]
  reg  meta_74_valid_0; // @[ICache.scala 34:21]
  reg  meta_74_valid_1; // @[ICache.scala 34:21]
  reg  meta_74_lru; // @[ICache.scala 34:21]
  reg  meta_75_valid_0; // @[ICache.scala 34:21]
  reg  meta_75_valid_1; // @[ICache.scala 34:21]
  reg  meta_75_lru; // @[ICache.scala 34:21]
  reg  meta_76_valid_0; // @[ICache.scala 34:21]
  reg  meta_76_valid_1; // @[ICache.scala 34:21]
  reg  meta_76_lru; // @[ICache.scala 34:21]
  reg  meta_77_valid_0; // @[ICache.scala 34:21]
  reg  meta_77_valid_1; // @[ICache.scala 34:21]
  reg  meta_77_lru; // @[ICache.scala 34:21]
  reg  meta_78_valid_0; // @[ICache.scala 34:21]
  reg  meta_78_valid_1; // @[ICache.scala 34:21]
  reg  meta_78_lru; // @[ICache.scala 34:21]
  reg  meta_79_valid_0; // @[ICache.scala 34:21]
  reg  meta_79_valid_1; // @[ICache.scala 34:21]
  reg  meta_79_lru; // @[ICache.scala 34:21]
  reg  meta_80_valid_0; // @[ICache.scala 34:21]
  reg  meta_80_valid_1; // @[ICache.scala 34:21]
  reg  meta_80_lru; // @[ICache.scala 34:21]
  reg  meta_81_valid_0; // @[ICache.scala 34:21]
  reg  meta_81_valid_1; // @[ICache.scala 34:21]
  reg  meta_81_lru; // @[ICache.scala 34:21]
  reg  meta_82_valid_0; // @[ICache.scala 34:21]
  reg  meta_82_valid_1; // @[ICache.scala 34:21]
  reg  meta_82_lru; // @[ICache.scala 34:21]
  reg  meta_83_valid_0; // @[ICache.scala 34:21]
  reg  meta_83_valid_1; // @[ICache.scala 34:21]
  reg  meta_83_lru; // @[ICache.scala 34:21]
  reg  meta_84_valid_0; // @[ICache.scala 34:21]
  reg  meta_84_valid_1; // @[ICache.scala 34:21]
  reg  meta_84_lru; // @[ICache.scala 34:21]
  reg  meta_85_valid_0; // @[ICache.scala 34:21]
  reg  meta_85_valid_1; // @[ICache.scala 34:21]
  reg  meta_85_lru; // @[ICache.scala 34:21]
  reg  meta_86_valid_0; // @[ICache.scala 34:21]
  reg  meta_86_valid_1; // @[ICache.scala 34:21]
  reg  meta_86_lru; // @[ICache.scala 34:21]
  reg  meta_87_valid_0; // @[ICache.scala 34:21]
  reg  meta_87_valid_1; // @[ICache.scala 34:21]
  reg  meta_87_lru; // @[ICache.scala 34:21]
  reg  meta_88_valid_0; // @[ICache.scala 34:21]
  reg  meta_88_valid_1; // @[ICache.scala 34:21]
  reg  meta_88_lru; // @[ICache.scala 34:21]
  reg  meta_89_valid_0; // @[ICache.scala 34:21]
  reg  meta_89_valid_1; // @[ICache.scala 34:21]
  reg  meta_89_lru; // @[ICache.scala 34:21]
  reg  meta_90_valid_0; // @[ICache.scala 34:21]
  reg  meta_90_valid_1; // @[ICache.scala 34:21]
  reg  meta_90_lru; // @[ICache.scala 34:21]
  reg  meta_91_valid_0; // @[ICache.scala 34:21]
  reg  meta_91_valid_1; // @[ICache.scala 34:21]
  reg  meta_91_lru; // @[ICache.scala 34:21]
  reg  meta_92_valid_0; // @[ICache.scala 34:21]
  reg  meta_92_valid_1; // @[ICache.scala 34:21]
  reg  meta_92_lru; // @[ICache.scala 34:21]
  reg  meta_93_valid_0; // @[ICache.scala 34:21]
  reg  meta_93_valid_1; // @[ICache.scala 34:21]
  reg  meta_93_lru; // @[ICache.scala 34:21]
  reg  meta_94_valid_0; // @[ICache.scala 34:21]
  reg  meta_94_valid_1; // @[ICache.scala 34:21]
  reg  meta_94_lru; // @[ICache.scala 34:21]
  reg  meta_95_valid_0; // @[ICache.scala 34:21]
  reg  meta_95_valid_1; // @[ICache.scala 34:21]
  reg  meta_95_lru; // @[ICache.scala 34:21]
  reg  meta_96_valid_0; // @[ICache.scala 34:21]
  reg  meta_96_valid_1; // @[ICache.scala 34:21]
  reg  meta_96_lru; // @[ICache.scala 34:21]
  reg  meta_97_valid_0; // @[ICache.scala 34:21]
  reg  meta_97_valid_1; // @[ICache.scala 34:21]
  reg  meta_97_lru; // @[ICache.scala 34:21]
  reg  meta_98_valid_0; // @[ICache.scala 34:21]
  reg  meta_98_valid_1; // @[ICache.scala 34:21]
  reg  meta_98_lru; // @[ICache.scala 34:21]
  reg  meta_99_valid_0; // @[ICache.scala 34:21]
  reg  meta_99_valid_1; // @[ICache.scala 34:21]
  reg  meta_99_lru; // @[ICache.scala 34:21]
  reg  meta_100_valid_0; // @[ICache.scala 34:21]
  reg  meta_100_valid_1; // @[ICache.scala 34:21]
  reg  meta_100_lru; // @[ICache.scala 34:21]
  reg  meta_101_valid_0; // @[ICache.scala 34:21]
  reg  meta_101_valid_1; // @[ICache.scala 34:21]
  reg  meta_101_lru; // @[ICache.scala 34:21]
  reg  meta_102_valid_0; // @[ICache.scala 34:21]
  reg  meta_102_valid_1; // @[ICache.scala 34:21]
  reg  meta_102_lru; // @[ICache.scala 34:21]
  reg  meta_103_valid_0; // @[ICache.scala 34:21]
  reg  meta_103_valid_1; // @[ICache.scala 34:21]
  reg  meta_103_lru; // @[ICache.scala 34:21]
  reg  meta_104_valid_0; // @[ICache.scala 34:21]
  reg  meta_104_valid_1; // @[ICache.scala 34:21]
  reg  meta_104_lru; // @[ICache.scala 34:21]
  reg  meta_105_valid_0; // @[ICache.scala 34:21]
  reg  meta_105_valid_1; // @[ICache.scala 34:21]
  reg  meta_105_lru; // @[ICache.scala 34:21]
  reg  meta_106_valid_0; // @[ICache.scala 34:21]
  reg  meta_106_valid_1; // @[ICache.scala 34:21]
  reg  meta_106_lru; // @[ICache.scala 34:21]
  reg  meta_107_valid_0; // @[ICache.scala 34:21]
  reg  meta_107_valid_1; // @[ICache.scala 34:21]
  reg  meta_107_lru; // @[ICache.scala 34:21]
  reg  meta_108_valid_0; // @[ICache.scala 34:21]
  reg  meta_108_valid_1; // @[ICache.scala 34:21]
  reg  meta_108_lru; // @[ICache.scala 34:21]
  reg  meta_109_valid_0; // @[ICache.scala 34:21]
  reg  meta_109_valid_1; // @[ICache.scala 34:21]
  reg  meta_109_lru; // @[ICache.scala 34:21]
  reg  meta_110_valid_0; // @[ICache.scala 34:21]
  reg  meta_110_valid_1; // @[ICache.scala 34:21]
  reg  meta_110_lru; // @[ICache.scala 34:21]
  reg  meta_111_valid_0; // @[ICache.scala 34:21]
  reg  meta_111_valid_1; // @[ICache.scala 34:21]
  reg  meta_111_lru; // @[ICache.scala 34:21]
  reg  meta_112_valid_0; // @[ICache.scala 34:21]
  reg  meta_112_valid_1; // @[ICache.scala 34:21]
  reg  meta_112_lru; // @[ICache.scala 34:21]
  reg  meta_113_valid_0; // @[ICache.scala 34:21]
  reg  meta_113_valid_1; // @[ICache.scala 34:21]
  reg  meta_113_lru; // @[ICache.scala 34:21]
  reg  meta_114_valid_0; // @[ICache.scala 34:21]
  reg  meta_114_valid_1; // @[ICache.scala 34:21]
  reg  meta_114_lru; // @[ICache.scala 34:21]
  reg  meta_115_valid_0; // @[ICache.scala 34:21]
  reg  meta_115_valid_1; // @[ICache.scala 34:21]
  reg  meta_115_lru; // @[ICache.scala 34:21]
  reg  meta_116_valid_0; // @[ICache.scala 34:21]
  reg  meta_116_valid_1; // @[ICache.scala 34:21]
  reg  meta_116_lru; // @[ICache.scala 34:21]
  reg  meta_117_valid_0; // @[ICache.scala 34:21]
  reg  meta_117_valid_1; // @[ICache.scala 34:21]
  reg  meta_117_lru; // @[ICache.scala 34:21]
  reg  meta_118_valid_0; // @[ICache.scala 34:21]
  reg  meta_118_valid_1; // @[ICache.scala 34:21]
  reg  meta_118_lru; // @[ICache.scala 34:21]
  reg  meta_119_valid_0; // @[ICache.scala 34:21]
  reg  meta_119_valid_1; // @[ICache.scala 34:21]
  reg  meta_119_lru; // @[ICache.scala 34:21]
  reg  meta_120_valid_0; // @[ICache.scala 34:21]
  reg  meta_120_valid_1; // @[ICache.scala 34:21]
  reg  meta_120_lru; // @[ICache.scala 34:21]
  reg  meta_121_valid_0; // @[ICache.scala 34:21]
  reg  meta_121_valid_1; // @[ICache.scala 34:21]
  reg  meta_121_lru; // @[ICache.scala 34:21]
  reg  meta_122_valid_0; // @[ICache.scala 34:21]
  reg  meta_122_valid_1; // @[ICache.scala 34:21]
  reg  meta_122_lru; // @[ICache.scala 34:21]
  reg  meta_123_valid_0; // @[ICache.scala 34:21]
  reg  meta_123_valid_1; // @[ICache.scala 34:21]
  reg  meta_123_lru; // @[ICache.scala 34:21]
  reg  meta_124_valid_0; // @[ICache.scala 34:21]
  reg  meta_124_valid_1; // @[ICache.scala 34:21]
  reg  meta_124_lru; // @[ICache.scala 34:21]
  reg  meta_125_valid_0; // @[ICache.scala 34:21]
  reg  meta_125_valid_1; // @[ICache.scala 34:21]
  reg  meta_125_lru; // @[ICache.scala 34:21]
  reg  meta_126_valid_0; // @[ICache.scala 34:21]
  reg  meta_126_valid_1; // @[ICache.scala 34:21]
  reg  meta_126_lru; // @[ICache.scala 34:21]
  reg  meta_127_valid_0; // @[ICache.scala 34:21]
  reg  meta_127_valid_1; // @[ICache.scala 34:21]
  reg  meta_127_lru; // @[ICache.scala 34:21]
  reg  meta_128_valid_0; // @[ICache.scala 34:21]
  reg  meta_128_valid_1; // @[ICache.scala 34:21]
  reg  meta_128_lru; // @[ICache.scala 34:21]
  reg  meta_129_valid_0; // @[ICache.scala 34:21]
  reg  meta_129_valid_1; // @[ICache.scala 34:21]
  reg  meta_129_lru; // @[ICache.scala 34:21]
  reg  meta_130_valid_0; // @[ICache.scala 34:21]
  reg  meta_130_valid_1; // @[ICache.scala 34:21]
  reg  meta_130_lru; // @[ICache.scala 34:21]
  reg  meta_131_valid_0; // @[ICache.scala 34:21]
  reg  meta_131_valid_1; // @[ICache.scala 34:21]
  reg  meta_131_lru; // @[ICache.scala 34:21]
  reg  meta_132_valid_0; // @[ICache.scala 34:21]
  reg  meta_132_valid_1; // @[ICache.scala 34:21]
  reg  meta_132_lru; // @[ICache.scala 34:21]
  reg  meta_133_valid_0; // @[ICache.scala 34:21]
  reg  meta_133_valid_1; // @[ICache.scala 34:21]
  reg  meta_133_lru; // @[ICache.scala 34:21]
  reg  meta_134_valid_0; // @[ICache.scala 34:21]
  reg  meta_134_valid_1; // @[ICache.scala 34:21]
  reg  meta_134_lru; // @[ICache.scala 34:21]
  reg  meta_135_valid_0; // @[ICache.scala 34:21]
  reg  meta_135_valid_1; // @[ICache.scala 34:21]
  reg  meta_135_lru; // @[ICache.scala 34:21]
  reg  meta_136_valid_0; // @[ICache.scala 34:21]
  reg  meta_136_valid_1; // @[ICache.scala 34:21]
  reg  meta_136_lru; // @[ICache.scala 34:21]
  reg  meta_137_valid_0; // @[ICache.scala 34:21]
  reg  meta_137_valid_1; // @[ICache.scala 34:21]
  reg  meta_137_lru; // @[ICache.scala 34:21]
  reg  meta_138_valid_0; // @[ICache.scala 34:21]
  reg  meta_138_valid_1; // @[ICache.scala 34:21]
  reg  meta_138_lru; // @[ICache.scala 34:21]
  reg  meta_139_valid_0; // @[ICache.scala 34:21]
  reg  meta_139_valid_1; // @[ICache.scala 34:21]
  reg  meta_139_lru; // @[ICache.scala 34:21]
  reg  meta_140_valid_0; // @[ICache.scala 34:21]
  reg  meta_140_valid_1; // @[ICache.scala 34:21]
  reg  meta_140_lru; // @[ICache.scala 34:21]
  reg  meta_141_valid_0; // @[ICache.scala 34:21]
  reg  meta_141_valid_1; // @[ICache.scala 34:21]
  reg  meta_141_lru; // @[ICache.scala 34:21]
  reg  meta_142_valid_0; // @[ICache.scala 34:21]
  reg  meta_142_valid_1; // @[ICache.scala 34:21]
  reg  meta_142_lru; // @[ICache.scala 34:21]
  reg  meta_143_valid_0; // @[ICache.scala 34:21]
  reg  meta_143_valid_1; // @[ICache.scala 34:21]
  reg  meta_143_lru; // @[ICache.scala 34:21]
  reg  meta_144_valid_0; // @[ICache.scala 34:21]
  reg  meta_144_valid_1; // @[ICache.scala 34:21]
  reg  meta_144_lru; // @[ICache.scala 34:21]
  reg  meta_145_valid_0; // @[ICache.scala 34:21]
  reg  meta_145_valid_1; // @[ICache.scala 34:21]
  reg  meta_145_lru; // @[ICache.scala 34:21]
  reg  meta_146_valid_0; // @[ICache.scala 34:21]
  reg  meta_146_valid_1; // @[ICache.scala 34:21]
  reg  meta_146_lru; // @[ICache.scala 34:21]
  reg  meta_147_valid_0; // @[ICache.scala 34:21]
  reg  meta_147_valid_1; // @[ICache.scala 34:21]
  reg  meta_147_lru; // @[ICache.scala 34:21]
  reg  meta_148_valid_0; // @[ICache.scala 34:21]
  reg  meta_148_valid_1; // @[ICache.scala 34:21]
  reg  meta_148_lru; // @[ICache.scala 34:21]
  reg  meta_149_valid_0; // @[ICache.scala 34:21]
  reg  meta_149_valid_1; // @[ICache.scala 34:21]
  reg  meta_149_lru; // @[ICache.scala 34:21]
  reg  meta_150_valid_0; // @[ICache.scala 34:21]
  reg  meta_150_valid_1; // @[ICache.scala 34:21]
  reg  meta_150_lru; // @[ICache.scala 34:21]
  reg  meta_151_valid_0; // @[ICache.scala 34:21]
  reg  meta_151_valid_1; // @[ICache.scala 34:21]
  reg  meta_151_lru; // @[ICache.scala 34:21]
  reg  meta_152_valid_0; // @[ICache.scala 34:21]
  reg  meta_152_valid_1; // @[ICache.scala 34:21]
  reg  meta_152_lru; // @[ICache.scala 34:21]
  reg  meta_153_valid_0; // @[ICache.scala 34:21]
  reg  meta_153_valid_1; // @[ICache.scala 34:21]
  reg  meta_153_lru; // @[ICache.scala 34:21]
  reg  meta_154_valid_0; // @[ICache.scala 34:21]
  reg  meta_154_valid_1; // @[ICache.scala 34:21]
  reg  meta_154_lru; // @[ICache.scala 34:21]
  reg  meta_155_valid_0; // @[ICache.scala 34:21]
  reg  meta_155_valid_1; // @[ICache.scala 34:21]
  reg  meta_155_lru; // @[ICache.scala 34:21]
  reg  meta_156_valid_0; // @[ICache.scala 34:21]
  reg  meta_156_valid_1; // @[ICache.scala 34:21]
  reg  meta_156_lru; // @[ICache.scala 34:21]
  reg  meta_157_valid_0; // @[ICache.scala 34:21]
  reg  meta_157_valid_1; // @[ICache.scala 34:21]
  reg  meta_157_lru; // @[ICache.scala 34:21]
  reg  meta_158_valid_0; // @[ICache.scala 34:21]
  reg  meta_158_valid_1; // @[ICache.scala 34:21]
  reg  meta_158_lru; // @[ICache.scala 34:21]
  reg  meta_159_valid_0; // @[ICache.scala 34:21]
  reg  meta_159_valid_1; // @[ICache.scala 34:21]
  reg  meta_159_lru; // @[ICache.scala 34:21]
  reg  meta_160_valid_0; // @[ICache.scala 34:21]
  reg  meta_160_valid_1; // @[ICache.scala 34:21]
  reg  meta_160_lru; // @[ICache.scala 34:21]
  reg  meta_161_valid_0; // @[ICache.scala 34:21]
  reg  meta_161_valid_1; // @[ICache.scala 34:21]
  reg  meta_161_lru; // @[ICache.scala 34:21]
  reg  meta_162_valid_0; // @[ICache.scala 34:21]
  reg  meta_162_valid_1; // @[ICache.scala 34:21]
  reg  meta_162_lru; // @[ICache.scala 34:21]
  reg  meta_163_valid_0; // @[ICache.scala 34:21]
  reg  meta_163_valid_1; // @[ICache.scala 34:21]
  reg  meta_163_lru; // @[ICache.scala 34:21]
  reg  meta_164_valid_0; // @[ICache.scala 34:21]
  reg  meta_164_valid_1; // @[ICache.scala 34:21]
  reg  meta_164_lru; // @[ICache.scala 34:21]
  reg  meta_165_valid_0; // @[ICache.scala 34:21]
  reg  meta_165_valid_1; // @[ICache.scala 34:21]
  reg  meta_165_lru; // @[ICache.scala 34:21]
  reg  meta_166_valid_0; // @[ICache.scala 34:21]
  reg  meta_166_valid_1; // @[ICache.scala 34:21]
  reg  meta_166_lru; // @[ICache.scala 34:21]
  reg  meta_167_valid_0; // @[ICache.scala 34:21]
  reg  meta_167_valid_1; // @[ICache.scala 34:21]
  reg  meta_167_lru; // @[ICache.scala 34:21]
  reg  meta_168_valid_0; // @[ICache.scala 34:21]
  reg  meta_168_valid_1; // @[ICache.scala 34:21]
  reg  meta_168_lru; // @[ICache.scala 34:21]
  reg  meta_169_valid_0; // @[ICache.scala 34:21]
  reg  meta_169_valid_1; // @[ICache.scala 34:21]
  reg  meta_169_lru; // @[ICache.scala 34:21]
  reg  meta_170_valid_0; // @[ICache.scala 34:21]
  reg  meta_170_valid_1; // @[ICache.scala 34:21]
  reg  meta_170_lru; // @[ICache.scala 34:21]
  reg  meta_171_valid_0; // @[ICache.scala 34:21]
  reg  meta_171_valid_1; // @[ICache.scala 34:21]
  reg  meta_171_lru; // @[ICache.scala 34:21]
  reg  meta_172_valid_0; // @[ICache.scala 34:21]
  reg  meta_172_valid_1; // @[ICache.scala 34:21]
  reg  meta_172_lru; // @[ICache.scala 34:21]
  reg  meta_173_valid_0; // @[ICache.scala 34:21]
  reg  meta_173_valid_1; // @[ICache.scala 34:21]
  reg  meta_173_lru; // @[ICache.scala 34:21]
  reg  meta_174_valid_0; // @[ICache.scala 34:21]
  reg  meta_174_valid_1; // @[ICache.scala 34:21]
  reg  meta_174_lru; // @[ICache.scala 34:21]
  reg  meta_175_valid_0; // @[ICache.scala 34:21]
  reg  meta_175_valid_1; // @[ICache.scala 34:21]
  reg  meta_175_lru; // @[ICache.scala 34:21]
  reg  meta_176_valid_0; // @[ICache.scala 34:21]
  reg  meta_176_valid_1; // @[ICache.scala 34:21]
  reg  meta_176_lru; // @[ICache.scala 34:21]
  reg  meta_177_valid_0; // @[ICache.scala 34:21]
  reg  meta_177_valid_1; // @[ICache.scala 34:21]
  reg  meta_177_lru; // @[ICache.scala 34:21]
  reg  meta_178_valid_0; // @[ICache.scala 34:21]
  reg  meta_178_valid_1; // @[ICache.scala 34:21]
  reg  meta_178_lru; // @[ICache.scala 34:21]
  reg  meta_179_valid_0; // @[ICache.scala 34:21]
  reg  meta_179_valid_1; // @[ICache.scala 34:21]
  reg  meta_179_lru; // @[ICache.scala 34:21]
  reg  meta_180_valid_0; // @[ICache.scala 34:21]
  reg  meta_180_valid_1; // @[ICache.scala 34:21]
  reg  meta_180_lru; // @[ICache.scala 34:21]
  reg  meta_181_valid_0; // @[ICache.scala 34:21]
  reg  meta_181_valid_1; // @[ICache.scala 34:21]
  reg  meta_181_lru; // @[ICache.scala 34:21]
  reg  meta_182_valid_0; // @[ICache.scala 34:21]
  reg  meta_182_valid_1; // @[ICache.scala 34:21]
  reg  meta_182_lru; // @[ICache.scala 34:21]
  reg  meta_183_valid_0; // @[ICache.scala 34:21]
  reg  meta_183_valid_1; // @[ICache.scala 34:21]
  reg  meta_183_lru; // @[ICache.scala 34:21]
  reg  meta_184_valid_0; // @[ICache.scala 34:21]
  reg  meta_184_valid_1; // @[ICache.scala 34:21]
  reg  meta_184_lru; // @[ICache.scala 34:21]
  reg  meta_185_valid_0; // @[ICache.scala 34:21]
  reg  meta_185_valid_1; // @[ICache.scala 34:21]
  reg  meta_185_lru; // @[ICache.scala 34:21]
  reg  meta_186_valid_0; // @[ICache.scala 34:21]
  reg  meta_186_valid_1; // @[ICache.scala 34:21]
  reg  meta_186_lru; // @[ICache.scala 34:21]
  reg  meta_187_valid_0; // @[ICache.scala 34:21]
  reg  meta_187_valid_1; // @[ICache.scala 34:21]
  reg  meta_187_lru; // @[ICache.scala 34:21]
  reg  meta_188_valid_0; // @[ICache.scala 34:21]
  reg  meta_188_valid_1; // @[ICache.scala 34:21]
  reg  meta_188_lru; // @[ICache.scala 34:21]
  reg  meta_189_valid_0; // @[ICache.scala 34:21]
  reg  meta_189_valid_1; // @[ICache.scala 34:21]
  reg  meta_189_lru; // @[ICache.scala 34:21]
  reg  meta_190_valid_0; // @[ICache.scala 34:21]
  reg  meta_190_valid_1; // @[ICache.scala 34:21]
  reg  meta_190_lru; // @[ICache.scala 34:21]
  reg  meta_191_valid_0; // @[ICache.scala 34:21]
  reg  meta_191_valid_1; // @[ICache.scala 34:21]
  reg  meta_191_lru; // @[ICache.scala 34:21]
  reg  meta_192_valid_0; // @[ICache.scala 34:21]
  reg  meta_192_valid_1; // @[ICache.scala 34:21]
  reg  meta_192_lru; // @[ICache.scala 34:21]
  reg  meta_193_valid_0; // @[ICache.scala 34:21]
  reg  meta_193_valid_1; // @[ICache.scala 34:21]
  reg  meta_193_lru; // @[ICache.scala 34:21]
  reg  meta_194_valid_0; // @[ICache.scala 34:21]
  reg  meta_194_valid_1; // @[ICache.scala 34:21]
  reg  meta_194_lru; // @[ICache.scala 34:21]
  reg  meta_195_valid_0; // @[ICache.scala 34:21]
  reg  meta_195_valid_1; // @[ICache.scala 34:21]
  reg  meta_195_lru; // @[ICache.scala 34:21]
  reg  meta_196_valid_0; // @[ICache.scala 34:21]
  reg  meta_196_valid_1; // @[ICache.scala 34:21]
  reg  meta_196_lru; // @[ICache.scala 34:21]
  reg  meta_197_valid_0; // @[ICache.scala 34:21]
  reg  meta_197_valid_1; // @[ICache.scala 34:21]
  reg  meta_197_lru; // @[ICache.scala 34:21]
  reg  meta_198_valid_0; // @[ICache.scala 34:21]
  reg  meta_198_valid_1; // @[ICache.scala 34:21]
  reg  meta_198_lru; // @[ICache.scala 34:21]
  reg  meta_199_valid_0; // @[ICache.scala 34:21]
  reg  meta_199_valid_1; // @[ICache.scala 34:21]
  reg  meta_199_lru; // @[ICache.scala 34:21]
  reg  meta_200_valid_0; // @[ICache.scala 34:21]
  reg  meta_200_valid_1; // @[ICache.scala 34:21]
  reg  meta_200_lru; // @[ICache.scala 34:21]
  reg  meta_201_valid_0; // @[ICache.scala 34:21]
  reg  meta_201_valid_1; // @[ICache.scala 34:21]
  reg  meta_201_lru; // @[ICache.scala 34:21]
  reg  meta_202_valid_0; // @[ICache.scala 34:21]
  reg  meta_202_valid_1; // @[ICache.scala 34:21]
  reg  meta_202_lru; // @[ICache.scala 34:21]
  reg  meta_203_valid_0; // @[ICache.scala 34:21]
  reg  meta_203_valid_1; // @[ICache.scala 34:21]
  reg  meta_203_lru; // @[ICache.scala 34:21]
  reg  meta_204_valid_0; // @[ICache.scala 34:21]
  reg  meta_204_valid_1; // @[ICache.scala 34:21]
  reg  meta_204_lru; // @[ICache.scala 34:21]
  reg  meta_205_valid_0; // @[ICache.scala 34:21]
  reg  meta_205_valid_1; // @[ICache.scala 34:21]
  reg  meta_205_lru; // @[ICache.scala 34:21]
  reg  meta_206_valid_0; // @[ICache.scala 34:21]
  reg  meta_206_valid_1; // @[ICache.scala 34:21]
  reg  meta_206_lru; // @[ICache.scala 34:21]
  reg  meta_207_valid_0; // @[ICache.scala 34:21]
  reg  meta_207_valid_1; // @[ICache.scala 34:21]
  reg  meta_207_lru; // @[ICache.scala 34:21]
  reg  meta_208_valid_0; // @[ICache.scala 34:21]
  reg  meta_208_valid_1; // @[ICache.scala 34:21]
  reg  meta_208_lru; // @[ICache.scala 34:21]
  reg  meta_209_valid_0; // @[ICache.scala 34:21]
  reg  meta_209_valid_1; // @[ICache.scala 34:21]
  reg  meta_209_lru; // @[ICache.scala 34:21]
  reg  meta_210_valid_0; // @[ICache.scala 34:21]
  reg  meta_210_valid_1; // @[ICache.scala 34:21]
  reg  meta_210_lru; // @[ICache.scala 34:21]
  reg  meta_211_valid_0; // @[ICache.scala 34:21]
  reg  meta_211_valid_1; // @[ICache.scala 34:21]
  reg  meta_211_lru; // @[ICache.scala 34:21]
  reg  meta_212_valid_0; // @[ICache.scala 34:21]
  reg  meta_212_valid_1; // @[ICache.scala 34:21]
  reg  meta_212_lru; // @[ICache.scala 34:21]
  reg  meta_213_valid_0; // @[ICache.scala 34:21]
  reg  meta_213_valid_1; // @[ICache.scala 34:21]
  reg  meta_213_lru; // @[ICache.scala 34:21]
  reg  meta_214_valid_0; // @[ICache.scala 34:21]
  reg  meta_214_valid_1; // @[ICache.scala 34:21]
  reg  meta_214_lru; // @[ICache.scala 34:21]
  reg  meta_215_valid_0; // @[ICache.scala 34:21]
  reg  meta_215_valid_1; // @[ICache.scala 34:21]
  reg  meta_215_lru; // @[ICache.scala 34:21]
  reg  meta_216_valid_0; // @[ICache.scala 34:21]
  reg  meta_216_valid_1; // @[ICache.scala 34:21]
  reg  meta_216_lru; // @[ICache.scala 34:21]
  reg  meta_217_valid_0; // @[ICache.scala 34:21]
  reg  meta_217_valid_1; // @[ICache.scala 34:21]
  reg  meta_217_lru; // @[ICache.scala 34:21]
  reg  meta_218_valid_0; // @[ICache.scala 34:21]
  reg  meta_218_valid_1; // @[ICache.scala 34:21]
  reg  meta_218_lru; // @[ICache.scala 34:21]
  reg  meta_219_valid_0; // @[ICache.scala 34:21]
  reg  meta_219_valid_1; // @[ICache.scala 34:21]
  reg  meta_219_lru; // @[ICache.scala 34:21]
  reg  meta_220_valid_0; // @[ICache.scala 34:21]
  reg  meta_220_valid_1; // @[ICache.scala 34:21]
  reg  meta_220_lru; // @[ICache.scala 34:21]
  reg  meta_221_valid_0; // @[ICache.scala 34:21]
  reg  meta_221_valid_1; // @[ICache.scala 34:21]
  reg  meta_221_lru; // @[ICache.scala 34:21]
  reg  meta_222_valid_0; // @[ICache.scala 34:21]
  reg  meta_222_valid_1; // @[ICache.scala 34:21]
  reg  meta_222_lru; // @[ICache.scala 34:21]
  reg  meta_223_valid_0; // @[ICache.scala 34:21]
  reg  meta_223_valid_1; // @[ICache.scala 34:21]
  reg  meta_223_lru; // @[ICache.scala 34:21]
  reg  meta_224_valid_0; // @[ICache.scala 34:21]
  reg  meta_224_valid_1; // @[ICache.scala 34:21]
  reg  meta_224_lru; // @[ICache.scala 34:21]
  reg  meta_225_valid_0; // @[ICache.scala 34:21]
  reg  meta_225_valid_1; // @[ICache.scala 34:21]
  reg  meta_225_lru; // @[ICache.scala 34:21]
  reg  meta_226_valid_0; // @[ICache.scala 34:21]
  reg  meta_226_valid_1; // @[ICache.scala 34:21]
  reg  meta_226_lru; // @[ICache.scala 34:21]
  reg  meta_227_valid_0; // @[ICache.scala 34:21]
  reg  meta_227_valid_1; // @[ICache.scala 34:21]
  reg  meta_227_lru; // @[ICache.scala 34:21]
  reg  meta_228_valid_0; // @[ICache.scala 34:21]
  reg  meta_228_valid_1; // @[ICache.scala 34:21]
  reg  meta_228_lru; // @[ICache.scala 34:21]
  reg  meta_229_valid_0; // @[ICache.scala 34:21]
  reg  meta_229_valid_1; // @[ICache.scala 34:21]
  reg  meta_229_lru; // @[ICache.scala 34:21]
  reg  meta_230_valid_0; // @[ICache.scala 34:21]
  reg  meta_230_valid_1; // @[ICache.scala 34:21]
  reg  meta_230_lru; // @[ICache.scala 34:21]
  reg  meta_231_valid_0; // @[ICache.scala 34:21]
  reg  meta_231_valid_1; // @[ICache.scala 34:21]
  reg  meta_231_lru; // @[ICache.scala 34:21]
  reg  meta_232_valid_0; // @[ICache.scala 34:21]
  reg  meta_232_valid_1; // @[ICache.scala 34:21]
  reg  meta_232_lru; // @[ICache.scala 34:21]
  reg  meta_233_valid_0; // @[ICache.scala 34:21]
  reg  meta_233_valid_1; // @[ICache.scala 34:21]
  reg  meta_233_lru; // @[ICache.scala 34:21]
  reg  meta_234_valid_0; // @[ICache.scala 34:21]
  reg  meta_234_valid_1; // @[ICache.scala 34:21]
  reg  meta_234_lru; // @[ICache.scala 34:21]
  reg  meta_235_valid_0; // @[ICache.scala 34:21]
  reg  meta_235_valid_1; // @[ICache.scala 34:21]
  reg  meta_235_lru; // @[ICache.scala 34:21]
  reg  meta_236_valid_0; // @[ICache.scala 34:21]
  reg  meta_236_valid_1; // @[ICache.scala 34:21]
  reg  meta_236_lru; // @[ICache.scala 34:21]
  reg  meta_237_valid_0; // @[ICache.scala 34:21]
  reg  meta_237_valid_1; // @[ICache.scala 34:21]
  reg  meta_237_lru; // @[ICache.scala 34:21]
  reg  meta_238_valid_0; // @[ICache.scala 34:21]
  reg  meta_238_valid_1; // @[ICache.scala 34:21]
  reg  meta_238_lru; // @[ICache.scala 34:21]
  reg  meta_239_valid_0; // @[ICache.scala 34:21]
  reg  meta_239_valid_1; // @[ICache.scala 34:21]
  reg  meta_239_lru; // @[ICache.scala 34:21]
  reg  meta_240_valid_0; // @[ICache.scala 34:21]
  reg  meta_240_valid_1; // @[ICache.scala 34:21]
  reg  meta_240_lru; // @[ICache.scala 34:21]
  reg  meta_241_valid_0; // @[ICache.scala 34:21]
  reg  meta_241_valid_1; // @[ICache.scala 34:21]
  reg  meta_241_lru; // @[ICache.scala 34:21]
  reg  meta_242_valid_0; // @[ICache.scala 34:21]
  reg  meta_242_valid_1; // @[ICache.scala 34:21]
  reg  meta_242_lru; // @[ICache.scala 34:21]
  reg  meta_243_valid_0; // @[ICache.scala 34:21]
  reg  meta_243_valid_1; // @[ICache.scala 34:21]
  reg  meta_243_lru; // @[ICache.scala 34:21]
  reg  meta_244_valid_0; // @[ICache.scala 34:21]
  reg  meta_244_valid_1; // @[ICache.scala 34:21]
  reg  meta_244_lru; // @[ICache.scala 34:21]
  reg  meta_245_valid_0; // @[ICache.scala 34:21]
  reg  meta_245_valid_1; // @[ICache.scala 34:21]
  reg  meta_245_lru; // @[ICache.scala 34:21]
  reg  meta_246_valid_0; // @[ICache.scala 34:21]
  reg  meta_246_valid_1; // @[ICache.scala 34:21]
  reg  meta_246_lru; // @[ICache.scala 34:21]
  reg  meta_247_valid_0; // @[ICache.scala 34:21]
  reg  meta_247_valid_1; // @[ICache.scala 34:21]
  reg  meta_247_lru; // @[ICache.scala 34:21]
  reg  meta_248_valid_0; // @[ICache.scala 34:21]
  reg  meta_248_valid_1; // @[ICache.scala 34:21]
  reg  meta_248_lru; // @[ICache.scala 34:21]
  reg  meta_249_valid_0; // @[ICache.scala 34:21]
  reg  meta_249_valid_1; // @[ICache.scala 34:21]
  reg  meta_249_lru; // @[ICache.scala 34:21]
  reg  meta_250_valid_0; // @[ICache.scala 34:21]
  reg  meta_250_valid_1; // @[ICache.scala 34:21]
  reg  meta_250_lru; // @[ICache.scala 34:21]
  reg  meta_251_valid_0; // @[ICache.scala 34:21]
  reg  meta_251_valid_1; // @[ICache.scala 34:21]
  reg  meta_251_lru; // @[ICache.scala 34:21]
  reg  meta_252_valid_0; // @[ICache.scala 34:21]
  reg  meta_252_valid_1; // @[ICache.scala 34:21]
  reg  meta_252_lru; // @[ICache.scala 34:21]
  reg  meta_253_valid_0; // @[ICache.scala 34:21]
  reg  meta_253_valid_1; // @[ICache.scala 34:21]
  reg  meta_253_lru; // @[ICache.scala 34:21]
  reg  meta_254_valid_0; // @[ICache.scala 34:21]
  reg  meta_254_valid_1; // @[ICache.scala 34:21]
  reg  meta_254_lru; // @[ICache.scala 34:21]
  reg  meta_255_valid_0; // @[ICache.scala 34:21]
  reg  meta_255_valid_1; // @[ICache.scala 34:21]
  reg  meta_255_lru; // @[ICache.scala 34:21]
  reg  meta_256_valid_0; // @[ICache.scala 34:21]
  reg  meta_256_valid_1; // @[ICache.scala 34:21]
  reg  meta_256_lru; // @[ICache.scala 34:21]
  reg  meta_257_valid_0; // @[ICache.scala 34:21]
  reg  meta_257_valid_1; // @[ICache.scala 34:21]
  reg  meta_257_lru; // @[ICache.scala 34:21]
  reg  meta_258_valid_0; // @[ICache.scala 34:21]
  reg  meta_258_valid_1; // @[ICache.scala 34:21]
  reg  meta_258_lru; // @[ICache.scala 34:21]
  reg  meta_259_valid_0; // @[ICache.scala 34:21]
  reg  meta_259_valid_1; // @[ICache.scala 34:21]
  reg  meta_259_lru; // @[ICache.scala 34:21]
  reg  meta_260_valid_0; // @[ICache.scala 34:21]
  reg  meta_260_valid_1; // @[ICache.scala 34:21]
  reg  meta_260_lru; // @[ICache.scala 34:21]
  reg  meta_261_valid_0; // @[ICache.scala 34:21]
  reg  meta_261_valid_1; // @[ICache.scala 34:21]
  reg  meta_261_lru; // @[ICache.scala 34:21]
  reg  meta_262_valid_0; // @[ICache.scala 34:21]
  reg  meta_262_valid_1; // @[ICache.scala 34:21]
  reg  meta_262_lru; // @[ICache.scala 34:21]
  reg  meta_263_valid_0; // @[ICache.scala 34:21]
  reg  meta_263_valid_1; // @[ICache.scala 34:21]
  reg  meta_263_lru; // @[ICache.scala 34:21]
  reg  meta_264_valid_0; // @[ICache.scala 34:21]
  reg  meta_264_valid_1; // @[ICache.scala 34:21]
  reg  meta_264_lru; // @[ICache.scala 34:21]
  reg  meta_265_valid_0; // @[ICache.scala 34:21]
  reg  meta_265_valid_1; // @[ICache.scala 34:21]
  reg  meta_265_lru; // @[ICache.scala 34:21]
  reg  meta_266_valid_0; // @[ICache.scala 34:21]
  reg  meta_266_valid_1; // @[ICache.scala 34:21]
  reg  meta_266_lru; // @[ICache.scala 34:21]
  reg  meta_267_valid_0; // @[ICache.scala 34:21]
  reg  meta_267_valid_1; // @[ICache.scala 34:21]
  reg  meta_267_lru; // @[ICache.scala 34:21]
  reg  meta_268_valid_0; // @[ICache.scala 34:21]
  reg  meta_268_valid_1; // @[ICache.scala 34:21]
  reg  meta_268_lru; // @[ICache.scala 34:21]
  reg  meta_269_valid_0; // @[ICache.scala 34:21]
  reg  meta_269_valid_1; // @[ICache.scala 34:21]
  reg  meta_269_lru; // @[ICache.scala 34:21]
  reg  meta_270_valid_0; // @[ICache.scala 34:21]
  reg  meta_270_valid_1; // @[ICache.scala 34:21]
  reg  meta_270_lru; // @[ICache.scala 34:21]
  reg  meta_271_valid_0; // @[ICache.scala 34:21]
  reg  meta_271_valid_1; // @[ICache.scala 34:21]
  reg  meta_271_lru; // @[ICache.scala 34:21]
  reg  meta_272_valid_0; // @[ICache.scala 34:21]
  reg  meta_272_valid_1; // @[ICache.scala 34:21]
  reg  meta_272_lru; // @[ICache.scala 34:21]
  reg  meta_273_valid_0; // @[ICache.scala 34:21]
  reg  meta_273_valid_1; // @[ICache.scala 34:21]
  reg  meta_273_lru; // @[ICache.scala 34:21]
  reg  meta_274_valid_0; // @[ICache.scala 34:21]
  reg  meta_274_valid_1; // @[ICache.scala 34:21]
  reg  meta_274_lru; // @[ICache.scala 34:21]
  reg  meta_275_valid_0; // @[ICache.scala 34:21]
  reg  meta_275_valid_1; // @[ICache.scala 34:21]
  reg  meta_275_lru; // @[ICache.scala 34:21]
  reg  meta_276_valid_0; // @[ICache.scala 34:21]
  reg  meta_276_valid_1; // @[ICache.scala 34:21]
  reg  meta_276_lru; // @[ICache.scala 34:21]
  reg  meta_277_valid_0; // @[ICache.scala 34:21]
  reg  meta_277_valid_1; // @[ICache.scala 34:21]
  reg  meta_277_lru; // @[ICache.scala 34:21]
  reg  meta_278_valid_0; // @[ICache.scala 34:21]
  reg  meta_278_valid_1; // @[ICache.scala 34:21]
  reg  meta_278_lru; // @[ICache.scala 34:21]
  reg  meta_279_valid_0; // @[ICache.scala 34:21]
  reg  meta_279_valid_1; // @[ICache.scala 34:21]
  reg  meta_279_lru; // @[ICache.scala 34:21]
  reg  meta_280_valid_0; // @[ICache.scala 34:21]
  reg  meta_280_valid_1; // @[ICache.scala 34:21]
  reg  meta_280_lru; // @[ICache.scala 34:21]
  reg  meta_281_valid_0; // @[ICache.scala 34:21]
  reg  meta_281_valid_1; // @[ICache.scala 34:21]
  reg  meta_281_lru; // @[ICache.scala 34:21]
  reg  meta_282_valid_0; // @[ICache.scala 34:21]
  reg  meta_282_valid_1; // @[ICache.scala 34:21]
  reg  meta_282_lru; // @[ICache.scala 34:21]
  reg  meta_283_valid_0; // @[ICache.scala 34:21]
  reg  meta_283_valid_1; // @[ICache.scala 34:21]
  reg  meta_283_lru; // @[ICache.scala 34:21]
  reg  meta_284_valid_0; // @[ICache.scala 34:21]
  reg  meta_284_valid_1; // @[ICache.scala 34:21]
  reg  meta_284_lru; // @[ICache.scala 34:21]
  reg  meta_285_valid_0; // @[ICache.scala 34:21]
  reg  meta_285_valid_1; // @[ICache.scala 34:21]
  reg  meta_285_lru; // @[ICache.scala 34:21]
  reg  meta_286_valid_0; // @[ICache.scala 34:21]
  reg  meta_286_valid_1; // @[ICache.scala 34:21]
  reg  meta_286_lru; // @[ICache.scala 34:21]
  reg  meta_287_valid_0; // @[ICache.scala 34:21]
  reg  meta_287_valid_1; // @[ICache.scala 34:21]
  reg  meta_287_lru; // @[ICache.scala 34:21]
  reg  meta_288_valid_0; // @[ICache.scala 34:21]
  reg  meta_288_valid_1; // @[ICache.scala 34:21]
  reg  meta_288_lru; // @[ICache.scala 34:21]
  reg  meta_289_valid_0; // @[ICache.scala 34:21]
  reg  meta_289_valid_1; // @[ICache.scala 34:21]
  reg  meta_289_lru; // @[ICache.scala 34:21]
  reg  meta_290_valid_0; // @[ICache.scala 34:21]
  reg  meta_290_valid_1; // @[ICache.scala 34:21]
  reg  meta_290_lru; // @[ICache.scala 34:21]
  reg  meta_291_valid_0; // @[ICache.scala 34:21]
  reg  meta_291_valid_1; // @[ICache.scala 34:21]
  reg  meta_291_lru; // @[ICache.scala 34:21]
  reg  meta_292_valid_0; // @[ICache.scala 34:21]
  reg  meta_292_valid_1; // @[ICache.scala 34:21]
  reg  meta_292_lru; // @[ICache.scala 34:21]
  reg  meta_293_valid_0; // @[ICache.scala 34:21]
  reg  meta_293_valid_1; // @[ICache.scala 34:21]
  reg  meta_293_lru; // @[ICache.scala 34:21]
  reg  meta_294_valid_0; // @[ICache.scala 34:21]
  reg  meta_294_valid_1; // @[ICache.scala 34:21]
  reg  meta_294_lru; // @[ICache.scala 34:21]
  reg  meta_295_valid_0; // @[ICache.scala 34:21]
  reg  meta_295_valid_1; // @[ICache.scala 34:21]
  reg  meta_295_lru; // @[ICache.scala 34:21]
  reg  meta_296_valid_0; // @[ICache.scala 34:21]
  reg  meta_296_valid_1; // @[ICache.scala 34:21]
  reg  meta_296_lru; // @[ICache.scala 34:21]
  reg  meta_297_valid_0; // @[ICache.scala 34:21]
  reg  meta_297_valid_1; // @[ICache.scala 34:21]
  reg  meta_297_lru; // @[ICache.scala 34:21]
  reg  meta_298_valid_0; // @[ICache.scala 34:21]
  reg  meta_298_valid_1; // @[ICache.scala 34:21]
  reg  meta_298_lru; // @[ICache.scala 34:21]
  reg  meta_299_valid_0; // @[ICache.scala 34:21]
  reg  meta_299_valid_1; // @[ICache.scala 34:21]
  reg  meta_299_lru; // @[ICache.scala 34:21]
  reg  meta_300_valid_0; // @[ICache.scala 34:21]
  reg  meta_300_valid_1; // @[ICache.scala 34:21]
  reg  meta_300_lru; // @[ICache.scala 34:21]
  reg  meta_301_valid_0; // @[ICache.scala 34:21]
  reg  meta_301_valid_1; // @[ICache.scala 34:21]
  reg  meta_301_lru; // @[ICache.scala 34:21]
  reg  meta_302_valid_0; // @[ICache.scala 34:21]
  reg  meta_302_valid_1; // @[ICache.scala 34:21]
  reg  meta_302_lru; // @[ICache.scala 34:21]
  reg  meta_303_valid_0; // @[ICache.scala 34:21]
  reg  meta_303_valid_1; // @[ICache.scala 34:21]
  reg  meta_303_lru; // @[ICache.scala 34:21]
  reg  meta_304_valid_0; // @[ICache.scala 34:21]
  reg  meta_304_valid_1; // @[ICache.scala 34:21]
  reg  meta_304_lru; // @[ICache.scala 34:21]
  reg  meta_305_valid_0; // @[ICache.scala 34:21]
  reg  meta_305_valid_1; // @[ICache.scala 34:21]
  reg  meta_305_lru; // @[ICache.scala 34:21]
  reg  meta_306_valid_0; // @[ICache.scala 34:21]
  reg  meta_306_valid_1; // @[ICache.scala 34:21]
  reg  meta_306_lru; // @[ICache.scala 34:21]
  reg  meta_307_valid_0; // @[ICache.scala 34:21]
  reg  meta_307_valid_1; // @[ICache.scala 34:21]
  reg  meta_307_lru; // @[ICache.scala 34:21]
  reg  meta_308_valid_0; // @[ICache.scala 34:21]
  reg  meta_308_valid_1; // @[ICache.scala 34:21]
  reg  meta_308_lru; // @[ICache.scala 34:21]
  reg  meta_309_valid_0; // @[ICache.scala 34:21]
  reg  meta_309_valid_1; // @[ICache.scala 34:21]
  reg  meta_309_lru; // @[ICache.scala 34:21]
  reg  meta_310_valid_0; // @[ICache.scala 34:21]
  reg  meta_310_valid_1; // @[ICache.scala 34:21]
  reg  meta_310_lru; // @[ICache.scala 34:21]
  reg  meta_311_valid_0; // @[ICache.scala 34:21]
  reg  meta_311_valid_1; // @[ICache.scala 34:21]
  reg  meta_311_lru; // @[ICache.scala 34:21]
  reg  meta_312_valid_0; // @[ICache.scala 34:21]
  reg  meta_312_valid_1; // @[ICache.scala 34:21]
  reg  meta_312_lru; // @[ICache.scala 34:21]
  reg  meta_313_valid_0; // @[ICache.scala 34:21]
  reg  meta_313_valid_1; // @[ICache.scala 34:21]
  reg  meta_313_lru; // @[ICache.scala 34:21]
  reg  meta_314_valid_0; // @[ICache.scala 34:21]
  reg  meta_314_valid_1; // @[ICache.scala 34:21]
  reg  meta_314_lru; // @[ICache.scala 34:21]
  reg  meta_315_valid_0; // @[ICache.scala 34:21]
  reg  meta_315_valid_1; // @[ICache.scala 34:21]
  reg  meta_315_lru; // @[ICache.scala 34:21]
  reg  meta_316_valid_0; // @[ICache.scala 34:21]
  reg  meta_316_valid_1; // @[ICache.scala 34:21]
  reg  meta_316_lru; // @[ICache.scala 34:21]
  reg  meta_317_valid_0; // @[ICache.scala 34:21]
  reg  meta_317_valid_1; // @[ICache.scala 34:21]
  reg  meta_317_lru; // @[ICache.scala 34:21]
  reg  meta_318_valid_0; // @[ICache.scala 34:21]
  reg  meta_318_valid_1; // @[ICache.scala 34:21]
  reg  meta_318_lru; // @[ICache.scala 34:21]
  reg  meta_319_valid_0; // @[ICache.scala 34:21]
  reg  meta_319_valid_1; // @[ICache.scala 34:21]
  reg  meta_319_lru; // @[ICache.scala 34:21]
  reg  meta_320_valid_0; // @[ICache.scala 34:21]
  reg  meta_320_valid_1; // @[ICache.scala 34:21]
  reg  meta_320_lru; // @[ICache.scala 34:21]
  reg  meta_321_valid_0; // @[ICache.scala 34:21]
  reg  meta_321_valid_1; // @[ICache.scala 34:21]
  reg  meta_321_lru; // @[ICache.scala 34:21]
  reg  meta_322_valid_0; // @[ICache.scala 34:21]
  reg  meta_322_valid_1; // @[ICache.scala 34:21]
  reg  meta_322_lru; // @[ICache.scala 34:21]
  reg  meta_323_valid_0; // @[ICache.scala 34:21]
  reg  meta_323_valid_1; // @[ICache.scala 34:21]
  reg  meta_323_lru; // @[ICache.scala 34:21]
  reg  meta_324_valid_0; // @[ICache.scala 34:21]
  reg  meta_324_valid_1; // @[ICache.scala 34:21]
  reg  meta_324_lru; // @[ICache.scala 34:21]
  reg  meta_325_valid_0; // @[ICache.scala 34:21]
  reg  meta_325_valid_1; // @[ICache.scala 34:21]
  reg  meta_325_lru; // @[ICache.scala 34:21]
  reg  meta_326_valid_0; // @[ICache.scala 34:21]
  reg  meta_326_valid_1; // @[ICache.scala 34:21]
  reg  meta_326_lru; // @[ICache.scala 34:21]
  reg  meta_327_valid_0; // @[ICache.scala 34:21]
  reg  meta_327_valid_1; // @[ICache.scala 34:21]
  reg  meta_327_lru; // @[ICache.scala 34:21]
  reg  meta_328_valid_0; // @[ICache.scala 34:21]
  reg  meta_328_valid_1; // @[ICache.scala 34:21]
  reg  meta_328_lru; // @[ICache.scala 34:21]
  reg  meta_329_valid_0; // @[ICache.scala 34:21]
  reg  meta_329_valid_1; // @[ICache.scala 34:21]
  reg  meta_329_lru; // @[ICache.scala 34:21]
  reg  meta_330_valid_0; // @[ICache.scala 34:21]
  reg  meta_330_valid_1; // @[ICache.scala 34:21]
  reg  meta_330_lru; // @[ICache.scala 34:21]
  reg  meta_331_valid_0; // @[ICache.scala 34:21]
  reg  meta_331_valid_1; // @[ICache.scala 34:21]
  reg  meta_331_lru; // @[ICache.scala 34:21]
  reg  meta_332_valid_0; // @[ICache.scala 34:21]
  reg  meta_332_valid_1; // @[ICache.scala 34:21]
  reg  meta_332_lru; // @[ICache.scala 34:21]
  reg  meta_333_valid_0; // @[ICache.scala 34:21]
  reg  meta_333_valid_1; // @[ICache.scala 34:21]
  reg  meta_333_lru; // @[ICache.scala 34:21]
  reg  meta_334_valid_0; // @[ICache.scala 34:21]
  reg  meta_334_valid_1; // @[ICache.scala 34:21]
  reg  meta_334_lru; // @[ICache.scala 34:21]
  reg  meta_335_valid_0; // @[ICache.scala 34:21]
  reg  meta_335_valid_1; // @[ICache.scala 34:21]
  reg  meta_335_lru; // @[ICache.scala 34:21]
  reg  meta_336_valid_0; // @[ICache.scala 34:21]
  reg  meta_336_valid_1; // @[ICache.scala 34:21]
  reg  meta_336_lru; // @[ICache.scala 34:21]
  reg  meta_337_valid_0; // @[ICache.scala 34:21]
  reg  meta_337_valid_1; // @[ICache.scala 34:21]
  reg  meta_337_lru; // @[ICache.scala 34:21]
  reg  meta_338_valid_0; // @[ICache.scala 34:21]
  reg  meta_338_valid_1; // @[ICache.scala 34:21]
  reg  meta_338_lru; // @[ICache.scala 34:21]
  reg  meta_339_valid_0; // @[ICache.scala 34:21]
  reg  meta_339_valid_1; // @[ICache.scala 34:21]
  reg  meta_339_lru; // @[ICache.scala 34:21]
  reg  meta_340_valid_0; // @[ICache.scala 34:21]
  reg  meta_340_valid_1; // @[ICache.scala 34:21]
  reg  meta_340_lru; // @[ICache.scala 34:21]
  reg  meta_341_valid_0; // @[ICache.scala 34:21]
  reg  meta_341_valid_1; // @[ICache.scala 34:21]
  reg  meta_341_lru; // @[ICache.scala 34:21]
  reg  meta_342_valid_0; // @[ICache.scala 34:21]
  reg  meta_342_valid_1; // @[ICache.scala 34:21]
  reg  meta_342_lru; // @[ICache.scala 34:21]
  reg  meta_343_valid_0; // @[ICache.scala 34:21]
  reg  meta_343_valid_1; // @[ICache.scala 34:21]
  reg  meta_343_lru; // @[ICache.scala 34:21]
  reg  meta_344_valid_0; // @[ICache.scala 34:21]
  reg  meta_344_valid_1; // @[ICache.scala 34:21]
  reg  meta_344_lru; // @[ICache.scala 34:21]
  reg  meta_345_valid_0; // @[ICache.scala 34:21]
  reg  meta_345_valid_1; // @[ICache.scala 34:21]
  reg  meta_345_lru; // @[ICache.scala 34:21]
  reg  meta_346_valid_0; // @[ICache.scala 34:21]
  reg  meta_346_valid_1; // @[ICache.scala 34:21]
  reg  meta_346_lru; // @[ICache.scala 34:21]
  reg  meta_347_valid_0; // @[ICache.scala 34:21]
  reg  meta_347_valid_1; // @[ICache.scala 34:21]
  reg  meta_347_lru; // @[ICache.scala 34:21]
  reg  meta_348_valid_0; // @[ICache.scala 34:21]
  reg  meta_348_valid_1; // @[ICache.scala 34:21]
  reg  meta_348_lru; // @[ICache.scala 34:21]
  reg  meta_349_valid_0; // @[ICache.scala 34:21]
  reg  meta_349_valid_1; // @[ICache.scala 34:21]
  reg  meta_349_lru; // @[ICache.scala 34:21]
  reg  meta_350_valid_0; // @[ICache.scala 34:21]
  reg  meta_350_valid_1; // @[ICache.scala 34:21]
  reg  meta_350_lru; // @[ICache.scala 34:21]
  reg  meta_351_valid_0; // @[ICache.scala 34:21]
  reg  meta_351_valid_1; // @[ICache.scala 34:21]
  reg  meta_351_lru; // @[ICache.scala 34:21]
  reg  meta_352_valid_0; // @[ICache.scala 34:21]
  reg  meta_352_valid_1; // @[ICache.scala 34:21]
  reg  meta_352_lru; // @[ICache.scala 34:21]
  reg  meta_353_valid_0; // @[ICache.scala 34:21]
  reg  meta_353_valid_1; // @[ICache.scala 34:21]
  reg  meta_353_lru; // @[ICache.scala 34:21]
  reg  meta_354_valid_0; // @[ICache.scala 34:21]
  reg  meta_354_valid_1; // @[ICache.scala 34:21]
  reg  meta_354_lru; // @[ICache.scala 34:21]
  reg  meta_355_valid_0; // @[ICache.scala 34:21]
  reg  meta_355_valid_1; // @[ICache.scala 34:21]
  reg  meta_355_lru; // @[ICache.scala 34:21]
  reg  meta_356_valid_0; // @[ICache.scala 34:21]
  reg  meta_356_valid_1; // @[ICache.scala 34:21]
  reg  meta_356_lru; // @[ICache.scala 34:21]
  reg  meta_357_valid_0; // @[ICache.scala 34:21]
  reg  meta_357_valid_1; // @[ICache.scala 34:21]
  reg  meta_357_lru; // @[ICache.scala 34:21]
  reg  meta_358_valid_0; // @[ICache.scala 34:21]
  reg  meta_358_valid_1; // @[ICache.scala 34:21]
  reg  meta_358_lru; // @[ICache.scala 34:21]
  reg  meta_359_valid_0; // @[ICache.scala 34:21]
  reg  meta_359_valid_1; // @[ICache.scala 34:21]
  reg  meta_359_lru; // @[ICache.scala 34:21]
  reg  meta_360_valid_0; // @[ICache.scala 34:21]
  reg  meta_360_valid_1; // @[ICache.scala 34:21]
  reg  meta_360_lru; // @[ICache.scala 34:21]
  reg  meta_361_valid_0; // @[ICache.scala 34:21]
  reg  meta_361_valid_1; // @[ICache.scala 34:21]
  reg  meta_361_lru; // @[ICache.scala 34:21]
  reg  meta_362_valid_0; // @[ICache.scala 34:21]
  reg  meta_362_valid_1; // @[ICache.scala 34:21]
  reg  meta_362_lru; // @[ICache.scala 34:21]
  reg  meta_363_valid_0; // @[ICache.scala 34:21]
  reg  meta_363_valid_1; // @[ICache.scala 34:21]
  reg  meta_363_lru; // @[ICache.scala 34:21]
  reg  meta_364_valid_0; // @[ICache.scala 34:21]
  reg  meta_364_valid_1; // @[ICache.scala 34:21]
  reg  meta_364_lru; // @[ICache.scala 34:21]
  reg  meta_365_valid_0; // @[ICache.scala 34:21]
  reg  meta_365_valid_1; // @[ICache.scala 34:21]
  reg  meta_365_lru; // @[ICache.scala 34:21]
  reg  meta_366_valid_0; // @[ICache.scala 34:21]
  reg  meta_366_valid_1; // @[ICache.scala 34:21]
  reg  meta_366_lru; // @[ICache.scala 34:21]
  reg  meta_367_valid_0; // @[ICache.scala 34:21]
  reg  meta_367_valid_1; // @[ICache.scala 34:21]
  reg  meta_367_lru; // @[ICache.scala 34:21]
  reg  meta_368_valid_0; // @[ICache.scala 34:21]
  reg  meta_368_valid_1; // @[ICache.scala 34:21]
  reg  meta_368_lru; // @[ICache.scala 34:21]
  reg  meta_369_valid_0; // @[ICache.scala 34:21]
  reg  meta_369_valid_1; // @[ICache.scala 34:21]
  reg  meta_369_lru; // @[ICache.scala 34:21]
  reg  meta_370_valid_0; // @[ICache.scala 34:21]
  reg  meta_370_valid_1; // @[ICache.scala 34:21]
  reg  meta_370_lru; // @[ICache.scala 34:21]
  reg  meta_371_valid_0; // @[ICache.scala 34:21]
  reg  meta_371_valid_1; // @[ICache.scala 34:21]
  reg  meta_371_lru; // @[ICache.scala 34:21]
  reg  meta_372_valid_0; // @[ICache.scala 34:21]
  reg  meta_372_valid_1; // @[ICache.scala 34:21]
  reg  meta_372_lru; // @[ICache.scala 34:21]
  reg  meta_373_valid_0; // @[ICache.scala 34:21]
  reg  meta_373_valid_1; // @[ICache.scala 34:21]
  reg  meta_373_lru; // @[ICache.scala 34:21]
  reg  meta_374_valid_0; // @[ICache.scala 34:21]
  reg  meta_374_valid_1; // @[ICache.scala 34:21]
  reg  meta_374_lru; // @[ICache.scala 34:21]
  reg  meta_375_valid_0; // @[ICache.scala 34:21]
  reg  meta_375_valid_1; // @[ICache.scala 34:21]
  reg  meta_375_lru; // @[ICache.scala 34:21]
  reg  meta_376_valid_0; // @[ICache.scala 34:21]
  reg  meta_376_valid_1; // @[ICache.scala 34:21]
  reg  meta_376_lru; // @[ICache.scala 34:21]
  reg  meta_377_valid_0; // @[ICache.scala 34:21]
  reg  meta_377_valid_1; // @[ICache.scala 34:21]
  reg  meta_377_lru; // @[ICache.scala 34:21]
  reg  meta_378_valid_0; // @[ICache.scala 34:21]
  reg  meta_378_valid_1; // @[ICache.scala 34:21]
  reg  meta_378_lru; // @[ICache.scala 34:21]
  reg  meta_379_valid_0; // @[ICache.scala 34:21]
  reg  meta_379_valid_1; // @[ICache.scala 34:21]
  reg  meta_379_lru; // @[ICache.scala 34:21]
  reg  meta_380_valid_0; // @[ICache.scala 34:21]
  reg  meta_380_valid_1; // @[ICache.scala 34:21]
  reg  meta_380_lru; // @[ICache.scala 34:21]
  reg  meta_381_valid_0; // @[ICache.scala 34:21]
  reg  meta_381_valid_1; // @[ICache.scala 34:21]
  reg  meta_381_lru; // @[ICache.scala 34:21]
  reg  meta_382_valid_0; // @[ICache.scala 34:21]
  reg  meta_382_valid_1; // @[ICache.scala 34:21]
  reg  meta_382_lru; // @[ICache.scala 34:21]
  reg  meta_383_valid_0; // @[ICache.scala 34:21]
  reg  meta_383_valid_1; // @[ICache.scala 34:21]
  reg  meta_383_lru; // @[ICache.scala 34:21]
  reg  meta_384_valid_0; // @[ICache.scala 34:21]
  reg  meta_384_valid_1; // @[ICache.scala 34:21]
  reg  meta_384_lru; // @[ICache.scala 34:21]
  reg  meta_385_valid_0; // @[ICache.scala 34:21]
  reg  meta_385_valid_1; // @[ICache.scala 34:21]
  reg  meta_385_lru; // @[ICache.scala 34:21]
  reg  meta_386_valid_0; // @[ICache.scala 34:21]
  reg  meta_386_valid_1; // @[ICache.scala 34:21]
  reg  meta_386_lru; // @[ICache.scala 34:21]
  reg  meta_387_valid_0; // @[ICache.scala 34:21]
  reg  meta_387_valid_1; // @[ICache.scala 34:21]
  reg  meta_387_lru; // @[ICache.scala 34:21]
  reg  meta_388_valid_0; // @[ICache.scala 34:21]
  reg  meta_388_valid_1; // @[ICache.scala 34:21]
  reg  meta_388_lru; // @[ICache.scala 34:21]
  reg  meta_389_valid_0; // @[ICache.scala 34:21]
  reg  meta_389_valid_1; // @[ICache.scala 34:21]
  reg  meta_389_lru; // @[ICache.scala 34:21]
  reg  meta_390_valid_0; // @[ICache.scala 34:21]
  reg  meta_390_valid_1; // @[ICache.scala 34:21]
  reg  meta_390_lru; // @[ICache.scala 34:21]
  reg  meta_391_valid_0; // @[ICache.scala 34:21]
  reg  meta_391_valid_1; // @[ICache.scala 34:21]
  reg  meta_391_lru; // @[ICache.scala 34:21]
  reg  meta_392_valid_0; // @[ICache.scala 34:21]
  reg  meta_392_valid_1; // @[ICache.scala 34:21]
  reg  meta_392_lru; // @[ICache.scala 34:21]
  reg  meta_393_valid_0; // @[ICache.scala 34:21]
  reg  meta_393_valid_1; // @[ICache.scala 34:21]
  reg  meta_393_lru; // @[ICache.scala 34:21]
  reg  meta_394_valid_0; // @[ICache.scala 34:21]
  reg  meta_394_valid_1; // @[ICache.scala 34:21]
  reg  meta_394_lru; // @[ICache.scala 34:21]
  reg  meta_395_valid_0; // @[ICache.scala 34:21]
  reg  meta_395_valid_1; // @[ICache.scala 34:21]
  reg  meta_395_lru; // @[ICache.scala 34:21]
  reg  meta_396_valid_0; // @[ICache.scala 34:21]
  reg  meta_396_valid_1; // @[ICache.scala 34:21]
  reg  meta_396_lru; // @[ICache.scala 34:21]
  reg  meta_397_valid_0; // @[ICache.scala 34:21]
  reg  meta_397_valid_1; // @[ICache.scala 34:21]
  reg  meta_397_lru; // @[ICache.scala 34:21]
  reg  meta_398_valid_0; // @[ICache.scala 34:21]
  reg  meta_398_valid_1; // @[ICache.scala 34:21]
  reg  meta_398_lru; // @[ICache.scala 34:21]
  reg  meta_399_valid_0; // @[ICache.scala 34:21]
  reg  meta_399_valid_1; // @[ICache.scala 34:21]
  reg  meta_399_lru; // @[ICache.scala 34:21]
  reg  meta_400_valid_0; // @[ICache.scala 34:21]
  reg  meta_400_valid_1; // @[ICache.scala 34:21]
  reg  meta_400_lru; // @[ICache.scala 34:21]
  reg  meta_401_valid_0; // @[ICache.scala 34:21]
  reg  meta_401_valid_1; // @[ICache.scala 34:21]
  reg  meta_401_lru; // @[ICache.scala 34:21]
  reg  meta_402_valid_0; // @[ICache.scala 34:21]
  reg  meta_402_valid_1; // @[ICache.scala 34:21]
  reg  meta_402_lru; // @[ICache.scala 34:21]
  reg  meta_403_valid_0; // @[ICache.scala 34:21]
  reg  meta_403_valid_1; // @[ICache.scala 34:21]
  reg  meta_403_lru; // @[ICache.scala 34:21]
  reg  meta_404_valid_0; // @[ICache.scala 34:21]
  reg  meta_404_valid_1; // @[ICache.scala 34:21]
  reg  meta_404_lru; // @[ICache.scala 34:21]
  reg  meta_405_valid_0; // @[ICache.scala 34:21]
  reg  meta_405_valid_1; // @[ICache.scala 34:21]
  reg  meta_405_lru; // @[ICache.scala 34:21]
  reg  meta_406_valid_0; // @[ICache.scala 34:21]
  reg  meta_406_valid_1; // @[ICache.scala 34:21]
  reg  meta_406_lru; // @[ICache.scala 34:21]
  reg  meta_407_valid_0; // @[ICache.scala 34:21]
  reg  meta_407_valid_1; // @[ICache.scala 34:21]
  reg  meta_407_lru; // @[ICache.scala 34:21]
  reg  meta_408_valid_0; // @[ICache.scala 34:21]
  reg  meta_408_valid_1; // @[ICache.scala 34:21]
  reg  meta_408_lru; // @[ICache.scala 34:21]
  reg  meta_409_valid_0; // @[ICache.scala 34:21]
  reg  meta_409_valid_1; // @[ICache.scala 34:21]
  reg  meta_409_lru; // @[ICache.scala 34:21]
  reg  meta_410_valid_0; // @[ICache.scala 34:21]
  reg  meta_410_valid_1; // @[ICache.scala 34:21]
  reg  meta_410_lru; // @[ICache.scala 34:21]
  reg  meta_411_valid_0; // @[ICache.scala 34:21]
  reg  meta_411_valid_1; // @[ICache.scala 34:21]
  reg  meta_411_lru; // @[ICache.scala 34:21]
  reg  meta_412_valid_0; // @[ICache.scala 34:21]
  reg  meta_412_valid_1; // @[ICache.scala 34:21]
  reg  meta_412_lru; // @[ICache.scala 34:21]
  reg  meta_413_valid_0; // @[ICache.scala 34:21]
  reg  meta_413_valid_1; // @[ICache.scala 34:21]
  reg  meta_413_lru; // @[ICache.scala 34:21]
  reg  meta_414_valid_0; // @[ICache.scala 34:21]
  reg  meta_414_valid_1; // @[ICache.scala 34:21]
  reg  meta_414_lru; // @[ICache.scala 34:21]
  reg  meta_415_valid_0; // @[ICache.scala 34:21]
  reg  meta_415_valid_1; // @[ICache.scala 34:21]
  reg  meta_415_lru; // @[ICache.scala 34:21]
  reg  meta_416_valid_0; // @[ICache.scala 34:21]
  reg  meta_416_valid_1; // @[ICache.scala 34:21]
  reg  meta_416_lru; // @[ICache.scala 34:21]
  reg  meta_417_valid_0; // @[ICache.scala 34:21]
  reg  meta_417_valid_1; // @[ICache.scala 34:21]
  reg  meta_417_lru; // @[ICache.scala 34:21]
  reg  meta_418_valid_0; // @[ICache.scala 34:21]
  reg  meta_418_valid_1; // @[ICache.scala 34:21]
  reg  meta_418_lru; // @[ICache.scala 34:21]
  reg  meta_419_valid_0; // @[ICache.scala 34:21]
  reg  meta_419_valid_1; // @[ICache.scala 34:21]
  reg  meta_419_lru; // @[ICache.scala 34:21]
  reg  meta_420_valid_0; // @[ICache.scala 34:21]
  reg  meta_420_valid_1; // @[ICache.scala 34:21]
  reg  meta_420_lru; // @[ICache.scala 34:21]
  reg  meta_421_valid_0; // @[ICache.scala 34:21]
  reg  meta_421_valid_1; // @[ICache.scala 34:21]
  reg  meta_421_lru; // @[ICache.scala 34:21]
  reg  meta_422_valid_0; // @[ICache.scala 34:21]
  reg  meta_422_valid_1; // @[ICache.scala 34:21]
  reg  meta_422_lru; // @[ICache.scala 34:21]
  reg  meta_423_valid_0; // @[ICache.scala 34:21]
  reg  meta_423_valid_1; // @[ICache.scala 34:21]
  reg  meta_423_lru; // @[ICache.scala 34:21]
  reg  meta_424_valid_0; // @[ICache.scala 34:21]
  reg  meta_424_valid_1; // @[ICache.scala 34:21]
  reg  meta_424_lru; // @[ICache.scala 34:21]
  reg  meta_425_valid_0; // @[ICache.scala 34:21]
  reg  meta_425_valid_1; // @[ICache.scala 34:21]
  reg  meta_425_lru; // @[ICache.scala 34:21]
  reg  meta_426_valid_0; // @[ICache.scala 34:21]
  reg  meta_426_valid_1; // @[ICache.scala 34:21]
  reg  meta_426_lru; // @[ICache.scala 34:21]
  reg  meta_427_valid_0; // @[ICache.scala 34:21]
  reg  meta_427_valid_1; // @[ICache.scala 34:21]
  reg  meta_427_lru; // @[ICache.scala 34:21]
  reg  meta_428_valid_0; // @[ICache.scala 34:21]
  reg  meta_428_valid_1; // @[ICache.scala 34:21]
  reg  meta_428_lru; // @[ICache.scala 34:21]
  reg  meta_429_valid_0; // @[ICache.scala 34:21]
  reg  meta_429_valid_1; // @[ICache.scala 34:21]
  reg  meta_429_lru; // @[ICache.scala 34:21]
  reg  meta_430_valid_0; // @[ICache.scala 34:21]
  reg  meta_430_valid_1; // @[ICache.scala 34:21]
  reg  meta_430_lru; // @[ICache.scala 34:21]
  reg  meta_431_valid_0; // @[ICache.scala 34:21]
  reg  meta_431_valid_1; // @[ICache.scala 34:21]
  reg  meta_431_lru; // @[ICache.scala 34:21]
  reg  meta_432_valid_0; // @[ICache.scala 34:21]
  reg  meta_432_valid_1; // @[ICache.scala 34:21]
  reg  meta_432_lru; // @[ICache.scala 34:21]
  reg  meta_433_valid_0; // @[ICache.scala 34:21]
  reg  meta_433_valid_1; // @[ICache.scala 34:21]
  reg  meta_433_lru; // @[ICache.scala 34:21]
  reg  meta_434_valid_0; // @[ICache.scala 34:21]
  reg  meta_434_valid_1; // @[ICache.scala 34:21]
  reg  meta_434_lru; // @[ICache.scala 34:21]
  reg  meta_435_valid_0; // @[ICache.scala 34:21]
  reg  meta_435_valid_1; // @[ICache.scala 34:21]
  reg  meta_435_lru; // @[ICache.scala 34:21]
  reg  meta_436_valid_0; // @[ICache.scala 34:21]
  reg  meta_436_valid_1; // @[ICache.scala 34:21]
  reg  meta_436_lru; // @[ICache.scala 34:21]
  reg  meta_437_valid_0; // @[ICache.scala 34:21]
  reg  meta_437_valid_1; // @[ICache.scala 34:21]
  reg  meta_437_lru; // @[ICache.scala 34:21]
  reg  meta_438_valid_0; // @[ICache.scala 34:21]
  reg  meta_438_valid_1; // @[ICache.scala 34:21]
  reg  meta_438_lru; // @[ICache.scala 34:21]
  reg  meta_439_valid_0; // @[ICache.scala 34:21]
  reg  meta_439_valid_1; // @[ICache.scala 34:21]
  reg  meta_439_lru; // @[ICache.scala 34:21]
  reg  meta_440_valid_0; // @[ICache.scala 34:21]
  reg  meta_440_valid_1; // @[ICache.scala 34:21]
  reg  meta_440_lru; // @[ICache.scala 34:21]
  reg  meta_441_valid_0; // @[ICache.scala 34:21]
  reg  meta_441_valid_1; // @[ICache.scala 34:21]
  reg  meta_441_lru; // @[ICache.scala 34:21]
  reg  meta_442_valid_0; // @[ICache.scala 34:21]
  reg  meta_442_valid_1; // @[ICache.scala 34:21]
  reg  meta_442_lru; // @[ICache.scala 34:21]
  reg  meta_443_valid_0; // @[ICache.scala 34:21]
  reg  meta_443_valid_1; // @[ICache.scala 34:21]
  reg  meta_443_lru; // @[ICache.scala 34:21]
  reg  meta_444_valid_0; // @[ICache.scala 34:21]
  reg  meta_444_valid_1; // @[ICache.scala 34:21]
  reg  meta_444_lru; // @[ICache.scala 34:21]
  reg  meta_445_valid_0; // @[ICache.scala 34:21]
  reg  meta_445_valid_1; // @[ICache.scala 34:21]
  reg  meta_445_lru; // @[ICache.scala 34:21]
  reg  meta_446_valid_0; // @[ICache.scala 34:21]
  reg  meta_446_valid_1; // @[ICache.scala 34:21]
  reg  meta_446_lru; // @[ICache.scala 34:21]
  reg  meta_447_valid_0; // @[ICache.scala 34:21]
  reg  meta_447_valid_1; // @[ICache.scala 34:21]
  reg  meta_447_lru; // @[ICache.scala 34:21]
  reg  meta_448_valid_0; // @[ICache.scala 34:21]
  reg  meta_448_valid_1; // @[ICache.scala 34:21]
  reg  meta_448_lru; // @[ICache.scala 34:21]
  reg  meta_449_valid_0; // @[ICache.scala 34:21]
  reg  meta_449_valid_1; // @[ICache.scala 34:21]
  reg  meta_449_lru; // @[ICache.scala 34:21]
  reg  meta_450_valid_0; // @[ICache.scala 34:21]
  reg  meta_450_valid_1; // @[ICache.scala 34:21]
  reg  meta_450_lru; // @[ICache.scala 34:21]
  reg  meta_451_valid_0; // @[ICache.scala 34:21]
  reg  meta_451_valid_1; // @[ICache.scala 34:21]
  reg  meta_451_lru; // @[ICache.scala 34:21]
  reg  meta_452_valid_0; // @[ICache.scala 34:21]
  reg  meta_452_valid_1; // @[ICache.scala 34:21]
  reg  meta_452_lru; // @[ICache.scala 34:21]
  reg  meta_453_valid_0; // @[ICache.scala 34:21]
  reg  meta_453_valid_1; // @[ICache.scala 34:21]
  reg  meta_453_lru; // @[ICache.scala 34:21]
  reg  meta_454_valid_0; // @[ICache.scala 34:21]
  reg  meta_454_valid_1; // @[ICache.scala 34:21]
  reg  meta_454_lru; // @[ICache.scala 34:21]
  reg  meta_455_valid_0; // @[ICache.scala 34:21]
  reg  meta_455_valid_1; // @[ICache.scala 34:21]
  reg  meta_455_lru; // @[ICache.scala 34:21]
  reg  meta_456_valid_0; // @[ICache.scala 34:21]
  reg  meta_456_valid_1; // @[ICache.scala 34:21]
  reg  meta_456_lru; // @[ICache.scala 34:21]
  reg  meta_457_valid_0; // @[ICache.scala 34:21]
  reg  meta_457_valid_1; // @[ICache.scala 34:21]
  reg  meta_457_lru; // @[ICache.scala 34:21]
  reg  meta_458_valid_0; // @[ICache.scala 34:21]
  reg  meta_458_valid_1; // @[ICache.scala 34:21]
  reg  meta_458_lru; // @[ICache.scala 34:21]
  reg  meta_459_valid_0; // @[ICache.scala 34:21]
  reg  meta_459_valid_1; // @[ICache.scala 34:21]
  reg  meta_459_lru; // @[ICache.scala 34:21]
  reg  meta_460_valid_0; // @[ICache.scala 34:21]
  reg  meta_460_valid_1; // @[ICache.scala 34:21]
  reg  meta_460_lru; // @[ICache.scala 34:21]
  reg  meta_461_valid_0; // @[ICache.scala 34:21]
  reg  meta_461_valid_1; // @[ICache.scala 34:21]
  reg  meta_461_lru; // @[ICache.scala 34:21]
  reg  meta_462_valid_0; // @[ICache.scala 34:21]
  reg  meta_462_valid_1; // @[ICache.scala 34:21]
  reg  meta_462_lru; // @[ICache.scala 34:21]
  reg  meta_463_valid_0; // @[ICache.scala 34:21]
  reg  meta_463_valid_1; // @[ICache.scala 34:21]
  reg  meta_463_lru; // @[ICache.scala 34:21]
  reg  meta_464_valid_0; // @[ICache.scala 34:21]
  reg  meta_464_valid_1; // @[ICache.scala 34:21]
  reg  meta_464_lru; // @[ICache.scala 34:21]
  reg  meta_465_valid_0; // @[ICache.scala 34:21]
  reg  meta_465_valid_1; // @[ICache.scala 34:21]
  reg  meta_465_lru; // @[ICache.scala 34:21]
  reg  meta_466_valid_0; // @[ICache.scala 34:21]
  reg  meta_466_valid_1; // @[ICache.scala 34:21]
  reg  meta_466_lru; // @[ICache.scala 34:21]
  reg  meta_467_valid_0; // @[ICache.scala 34:21]
  reg  meta_467_valid_1; // @[ICache.scala 34:21]
  reg  meta_467_lru; // @[ICache.scala 34:21]
  reg  meta_468_valid_0; // @[ICache.scala 34:21]
  reg  meta_468_valid_1; // @[ICache.scala 34:21]
  reg  meta_468_lru; // @[ICache.scala 34:21]
  reg  meta_469_valid_0; // @[ICache.scala 34:21]
  reg  meta_469_valid_1; // @[ICache.scala 34:21]
  reg  meta_469_lru; // @[ICache.scala 34:21]
  reg  meta_470_valid_0; // @[ICache.scala 34:21]
  reg  meta_470_valid_1; // @[ICache.scala 34:21]
  reg  meta_470_lru; // @[ICache.scala 34:21]
  reg  meta_471_valid_0; // @[ICache.scala 34:21]
  reg  meta_471_valid_1; // @[ICache.scala 34:21]
  reg  meta_471_lru; // @[ICache.scala 34:21]
  reg  meta_472_valid_0; // @[ICache.scala 34:21]
  reg  meta_472_valid_1; // @[ICache.scala 34:21]
  reg  meta_472_lru; // @[ICache.scala 34:21]
  reg  meta_473_valid_0; // @[ICache.scala 34:21]
  reg  meta_473_valid_1; // @[ICache.scala 34:21]
  reg  meta_473_lru; // @[ICache.scala 34:21]
  reg  meta_474_valid_0; // @[ICache.scala 34:21]
  reg  meta_474_valid_1; // @[ICache.scala 34:21]
  reg  meta_474_lru; // @[ICache.scala 34:21]
  reg  meta_475_valid_0; // @[ICache.scala 34:21]
  reg  meta_475_valid_1; // @[ICache.scala 34:21]
  reg  meta_475_lru; // @[ICache.scala 34:21]
  reg  meta_476_valid_0; // @[ICache.scala 34:21]
  reg  meta_476_valid_1; // @[ICache.scala 34:21]
  reg  meta_476_lru; // @[ICache.scala 34:21]
  reg  meta_477_valid_0; // @[ICache.scala 34:21]
  reg  meta_477_valid_1; // @[ICache.scala 34:21]
  reg  meta_477_lru; // @[ICache.scala 34:21]
  reg  meta_478_valid_0; // @[ICache.scala 34:21]
  reg  meta_478_valid_1; // @[ICache.scala 34:21]
  reg  meta_478_lru; // @[ICache.scala 34:21]
  reg  meta_479_valid_0; // @[ICache.scala 34:21]
  reg  meta_479_valid_1; // @[ICache.scala 34:21]
  reg  meta_479_lru; // @[ICache.scala 34:21]
  reg  meta_480_valid_0; // @[ICache.scala 34:21]
  reg  meta_480_valid_1; // @[ICache.scala 34:21]
  reg  meta_480_lru; // @[ICache.scala 34:21]
  reg  meta_481_valid_0; // @[ICache.scala 34:21]
  reg  meta_481_valid_1; // @[ICache.scala 34:21]
  reg  meta_481_lru; // @[ICache.scala 34:21]
  reg  meta_482_valid_0; // @[ICache.scala 34:21]
  reg  meta_482_valid_1; // @[ICache.scala 34:21]
  reg  meta_482_lru; // @[ICache.scala 34:21]
  reg  meta_483_valid_0; // @[ICache.scala 34:21]
  reg  meta_483_valid_1; // @[ICache.scala 34:21]
  reg  meta_483_lru; // @[ICache.scala 34:21]
  reg  meta_484_valid_0; // @[ICache.scala 34:21]
  reg  meta_484_valid_1; // @[ICache.scala 34:21]
  reg  meta_484_lru; // @[ICache.scala 34:21]
  reg  meta_485_valid_0; // @[ICache.scala 34:21]
  reg  meta_485_valid_1; // @[ICache.scala 34:21]
  reg  meta_485_lru; // @[ICache.scala 34:21]
  reg  meta_486_valid_0; // @[ICache.scala 34:21]
  reg  meta_486_valid_1; // @[ICache.scala 34:21]
  reg  meta_486_lru; // @[ICache.scala 34:21]
  reg  meta_487_valid_0; // @[ICache.scala 34:21]
  reg  meta_487_valid_1; // @[ICache.scala 34:21]
  reg  meta_487_lru; // @[ICache.scala 34:21]
  reg  meta_488_valid_0; // @[ICache.scala 34:21]
  reg  meta_488_valid_1; // @[ICache.scala 34:21]
  reg  meta_488_lru; // @[ICache.scala 34:21]
  reg  meta_489_valid_0; // @[ICache.scala 34:21]
  reg  meta_489_valid_1; // @[ICache.scala 34:21]
  reg  meta_489_lru; // @[ICache.scala 34:21]
  reg  meta_490_valid_0; // @[ICache.scala 34:21]
  reg  meta_490_valid_1; // @[ICache.scala 34:21]
  reg  meta_490_lru; // @[ICache.scala 34:21]
  reg  meta_491_valid_0; // @[ICache.scala 34:21]
  reg  meta_491_valid_1; // @[ICache.scala 34:21]
  reg  meta_491_lru; // @[ICache.scala 34:21]
  reg  meta_492_valid_0; // @[ICache.scala 34:21]
  reg  meta_492_valid_1; // @[ICache.scala 34:21]
  reg  meta_492_lru; // @[ICache.scala 34:21]
  reg  meta_493_valid_0; // @[ICache.scala 34:21]
  reg  meta_493_valid_1; // @[ICache.scala 34:21]
  reg  meta_493_lru; // @[ICache.scala 34:21]
  reg  meta_494_valid_0; // @[ICache.scala 34:21]
  reg  meta_494_valid_1; // @[ICache.scala 34:21]
  reg  meta_494_lru; // @[ICache.scala 34:21]
  reg  meta_495_valid_0; // @[ICache.scala 34:21]
  reg  meta_495_valid_1; // @[ICache.scala 34:21]
  reg  meta_495_lru; // @[ICache.scala 34:21]
  reg  meta_496_valid_0; // @[ICache.scala 34:21]
  reg  meta_496_valid_1; // @[ICache.scala 34:21]
  reg  meta_496_lru; // @[ICache.scala 34:21]
  reg  meta_497_valid_0; // @[ICache.scala 34:21]
  reg  meta_497_valid_1; // @[ICache.scala 34:21]
  reg  meta_497_lru; // @[ICache.scala 34:21]
  reg  meta_498_valid_0; // @[ICache.scala 34:21]
  reg  meta_498_valid_1; // @[ICache.scala 34:21]
  reg  meta_498_lru; // @[ICache.scala 34:21]
  reg  meta_499_valid_0; // @[ICache.scala 34:21]
  reg  meta_499_valid_1; // @[ICache.scala 34:21]
  reg  meta_499_lru; // @[ICache.scala 34:21]
  reg  meta_500_valid_0; // @[ICache.scala 34:21]
  reg  meta_500_valid_1; // @[ICache.scala 34:21]
  reg  meta_500_lru; // @[ICache.scala 34:21]
  reg  meta_501_valid_0; // @[ICache.scala 34:21]
  reg  meta_501_valid_1; // @[ICache.scala 34:21]
  reg  meta_501_lru; // @[ICache.scala 34:21]
  reg  meta_502_valid_0; // @[ICache.scala 34:21]
  reg  meta_502_valid_1; // @[ICache.scala 34:21]
  reg  meta_502_lru; // @[ICache.scala 34:21]
  reg  meta_503_valid_0; // @[ICache.scala 34:21]
  reg  meta_503_valid_1; // @[ICache.scala 34:21]
  reg  meta_503_lru; // @[ICache.scala 34:21]
  reg  meta_504_valid_0; // @[ICache.scala 34:21]
  reg  meta_504_valid_1; // @[ICache.scala 34:21]
  reg  meta_504_lru; // @[ICache.scala 34:21]
  reg  meta_505_valid_0; // @[ICache.scala 34:21]
  reg  meta_505_valid_1; // @[ICache.scala 34:21]
  reg  meta_505_lru; // @[ICache.scala 34:21]
  reg  meta_506_valid_0; // @[ICache.scala 34:21]
  reg  meta_506_valid_1; // @[ICache.scala 34:21]
  reg  meta_506_lru; // @[ICache.scala 34:21]
  reg  meta_507_valid_0; // @[ICache.scala 34:21]
  reg  meta_507_valid_1; // @[ICache.scala 34:21]
  reg  meta_507_lru; // @[ICache.scala 34:21]
  reg  meta_508_valid_0; // @[ICache.scala 34:21]
  reg  meta_508_valid_1; // @[ICache.scala 34:21]
  reg  meta_508_lru; // @[ICache.scala 34:21]
  reg  meta_509_valid_0; // @[ICache.scala 34:21]
  reg  meta_509_valid_1; // @[ICache.scala 34:21]
  reg  meta_509_lru; // @[ICache.scala 34:21]
  reg  meta_510_valid_0; // @[ICache.scala 34:21]
  reg  meta_510_valid_1; // @[ICache.scala 34:21]
  reg  meta_510_lru; // @[ICache.scala 34:21]
  reg  meta_511_valid_0; // @[ICache.scala 34:21]
  reg  meta_511_valid_1; // @[ICache.scala 34:21]
  reg  meta_511_lru; // @[ICache.scala 34:21]
  reg [16:0] tlb_vpn; // @[ICache.scala 40:20]
  reg [16:0] tlb_ppn; // @[ICache.scala 40:20]
  reg  tlb_uncached; // @[ICache.scala 40:20]
  reg  tlb_valid; // @[ICache.scala 40:20]
  reg [2:0] state; // @[ICache.scala 48:81]
  wire  direct_mapped = io_cpu_addr_0[31:30] == 2'h2; // @[ICache.scala 50:46]
  wire  uncached = direct_mapped ? io_cpu_addr_0[29] : tlb_uncached; // @[ICache.scala 51:26]
  wire [19:0] _inst_tag_T_1 = {3'h0,io_cpu_addr_0[28:12]}; // @[Cat.scala 33:92]
  wire [19:0] inst_tag = direct_mapped ? _inst_tag_T_1 : {{3'd0}, tlb_ppn}; // @[ICache.scala 52:26]
  wire [19:0] inst_vpn = io_cpu_addr_0[31:12]; // @[ICache.scala 53:37]
  wire [31:0] inst_pa = {inst_tag,io_cpu_addr_0[11:0]}; // @[Cat.scala 33:92]
  wire [19:0] _GEN_13515 = {{3'd0}, tlb_vpn}; // @[ICache.scala 56:50]
  wire  translation_ok = direct_mapped | _GEN_13515 == inst_vpn & tlb_valid; // @[ICache.scala 56:38]
  reg [5:0] replace_line_addr; // @[ICache.scala 58:38]
  wire  _bram_addr_choose_next_T_1 = state != 3'h4; // @[ICache.scala 59:62]
  wire  bram_addr_choose_next = ~(state != 3'h0 & state != 3'h4); // @[ICache.scala 59:31]
  wire [31:0] _GEN_1 = bram_addr_choose_next ? io_cpu_addr_1 : io_cpu_addr_0; // @[ICache.scala 61:{58,58}]
  wire [5:0] bram_line_addr = _GEN_1[11:6]; // @[ICache.scala 62:58]
  reg [7:0] data_wen_0; // @[ICache.scala 66:30]
  reg [7:0] data_wen_1; // @[ICache.scala 66:30]
  reg  tag_wen_0; // @[ICache.scala 67:30]
  reg  tag_wen_1; // @[ICache.scala 67:30]
  reg [16:0] tag_ram_wdata; // @[ICache.scala 68:30]
  wire [16:0] cache_tag_0 = tag_ram_io_way_0_r_data; // @[ICache.scala 64:28 131:30]
  wire [19:0] _GEN_13516 = {{3'd0}, cache_tag_0}; // @[ICache.scala 132:46]
  wire [5:0] va_line_addr = io_cpu_addr_0[11:6]; // @[ICache.scala 80:36]
  wire  _GEN_5 = 6'h1 == va_line_addr ? meta_1_valid_0 : meta_0_valid_0; // @[ICache.scala 132:{59,59}]
  wire  _GEN_6 = 6'h2 == va_line_addr ? meta_2_valid_0 : _GEN_5; // @[ICache.scala 132:{59,59}]
  wire  _GEN_7 = 6'h3 == va_line_addr ? meta_3_valid_0 : _GEN_6; // @[ICache.scala 132:{59,59}]
  wire  _GEN_8 = 6'h4 == va_line_addr ? meta_4_valid_0 : _GEN_7; // @[ICache.scala 132:{59,59}]
  wire  _GEN_9 = 6'h5 == va_line_addr ? meta_5_valid_0 : _GEN_8; // @[ICache.scala 132:{59,59}]
  wire  _GEN_10 = 6'h6 == va_line_addr ? meta_6_valid_0 : _GEN_9; // @[ICache.scala 132:{59,59}]
  wire  _GEN_11 = 6'h7 == va_line_addr ? meta_7_valid_0 : _GEN_10; // @[ICache.scala 132:{59,59}]
  wire  _GEN_12 = 6'h8 == va_line_addr ? meta_8_valid_0 : _GEN_11; // @[ICache.scala 132:{59,59}]
  wire  _GEN_13 = 6'h9 == va_line_addr ? meta_9_valid_0 : _GEN_12; // @[ICache.scala 132:{59,59}]
  wire  _GEN_14 = 6'ha == va_line_addr ? meta_10_valid_0 : _GEN_13; // @[ICache.scala 132:{59,59}]
  wire  _GEN_15 = 6'hb == va_line_addr ? meta_11_valid_0 : _GEN_14; // @[ICache.scala 132:{59,59}]
  wire  _GEN_16 = 6'hc == va_line_addr ? meta_12_valid_0 : _GEN_15; // @[ICache.scala 132:{59,59}]
  wire  _GEN_17 = 6'hd == va_line_addr ? meta_13_valid_0 : _GEN_16; // @[ICache.scala 132:{59,59}]
  wire  _GEN_18 = 6'he == va_line_addr ? meta_14_valid_0 : _GEN_17; // @[ICache.scala 132:{59,59}]
  wire  _GEN_19 = 6'hf == va_line_addr ? meta_15_valid_0 : _GEN_18; // @[ICache.scala 132:{59,59}]
  wire  _GEN_20 = 6'h10 == va_line_addr ? meta_16_valid_0 : _GEN_19; // @[ICache.scala 132:{59,59}]
  wire  _GEN_21 = 6'h11 == va_line_addr ? meta_17_valid_0 : _GEN_20; // @[ICache.scala 132:{59,59}]
  wire  _GEN_22 = 6'h12 == va_line_addr ? meta_18_valid_0 : _GEN_21; // @[ICache.scala 132:{59,59}]
  wire  _GEN_23 = 6'h13 == va_line_addr ? meta_19_valid_0 : _GEN_22; // @[ICache.scala 132:{59,59}]
  wire  _GEN_24 = 6'h14 == va_line_addr ? meta_20_valid_0 : _GEN_23; // @[ICache.scala 132:{59,59}]
  wire  _GEN_25 = 6'h15 == va_line_addr ? meta_21_valid_0 : _GEN_24; // @[ICache.scala 132:{59,59}]
  wire  _GEN_26 = 6'h16 == va_line_addr ? meta_22_valid_0 : _GEN_25; // @[ICache.scala 132:{59,59}]
  wire  _GEN_27 = 6'h17 == va_line_addr ? meta_23_valid_0 : _GEN_26; // @[ICache.scala 132:{59,59}]
  wire  _GEN_28 = 6'h18 == va_line_addr ? meta_24_valid_0 : _GEN_27; // @[ICache.scala 132:{59,59}]
  wire  _GEN_29 = 6'h19 == va_line_addr ? meta_25_valid_0 : _GEN_28; // @[ICache.scala 132:{59,59}]
  wire  _GEN_30 = 6'h1a == va_line_addr ? meta_26_valid_0 : _GEN_29; // @[ICache.scala 132:{59,59}]
  wire  _GEN_31 = 6'h1b == va_line_addr ? meta_27_valid_0 : _GEN_30; // @[ICache.scala 132:{59,59}]
  wire  _GEN_32 = 6'h1c == va_line_addr ? meta_28_valid_0 : _GEN_31; // @[ICache.scala 132:{59,59}]
  wire  _GEN_33 = 6'h1d == va_line_addr ? meta_29_valid_0 : _GEN_32; // @[ICache.scala 132:{59,59}]
  wire  _GEN_34 = 6'h1e == va_line_addr ? meta_30_valid_0 : _GEN_33; // @[ICache.scala 132:{59,59}]
  wire  _GEN_35 = 6'h1f == va_line_addr ? meta_31_valid_0 : _GEN_34; // @[ICache.scala 132:{59,59}]
  wire  _GEN_36 = 6'h20 == va_line_addr ? meta_32_valid_0 : _GEN_35; // @[ICache.scala 132:{59,59}]
  wire  _GEN_37 = 6'h21 == va_line_addr ? meta_33_valid_0 : _GEN_36; // @[ICache.scala 132:{59,59}]
  wire  _GEN_38 = 6'h22 == va_line_addr ? meta_34_valid_0 : _GEN_37; // @[ICache.scala 132:{59,59}]
  wire  _GEN_39 = 6'h23 == va_line_addr ? meta_35_valid_0 : _GEN_38; // @[ICache.scala 132:{59,59}]
  wire  _GEN_40 = 6'h24 == va_line_addr ? meta_36_valid_0 : _GEN_39; // @[ICache.scala 132:{59,59}]
  wire  _GEN_41 = 6'h25 == va_line_addr ? meta_37_valid_0 : _GEN_40; // @[ICache.scala 132:{59,59}]
  wire  _GEN_42 = 6'h26 == va_line_addr ? meta_38_valid_0 : _GEN_41; // @[ICache.scala 132:{59,59}]
  wire  _GEN_43 = 6'h27 == va_line_addr ? meta_39_valid_0 : _GEN_42; // @[ICache.scala 132:{59,59}]
  wire  _GEN_44 = 6'h28 == va_line_addr ? meta_40_valid_0 : _GEN_43; // @[ICache.scala 132:{59,59}]
  wire  _GEN_45 = 6'h29 == va_line_addr ? meta_41_valid_0 : _GEN_44; // @[ICache.scala 132:{59,59}]
  wire  _GEN_46 = 6'h2a == va_line_addr ? meta_42_valid_0 : _GEN_45; // @[ICache.scala 132:{59,59}]
  wire  _GEN_47 = 6'h2b == va_line_addr ? meta_43_valid_0 : _GEN_46; // @[ICache.scala 132:{59,59}]
  wire  _GEN_48 = 6'h2c == va_line_addr ? meta_44_valid_0 : _GEN_47; // @[ICache.scala 132:{59,59}]
  wire  _GEN_49 = 6'h2d == va_line_addr ? meta_45_valid_0 : _GEN_48; // @[ICache.scala 132:{59,59}]
  wire  _GEN_50 = 6'h2e == va_line_addr ? meta_46_valid_0 : _GEN_49; // @[ICache.scala 132:{59,59}]
  wire  _GEN_51 = 6'h2f == va_line_addr ? meta_47_valid_0 : _GEN_50; // @[ICache.scala 132:{59,59}]
  wire  _GEN_52 = 6'h30 == va_line_addr ? meta_48_valid_0 : _GEN_51; // @[ICache.scala 132:{59,59}]
  wire  _GEN_53 = 6'h31 == va_line_addr ? meta_49_valid_0 : _GEN_52; // @[ICache.scala 132:{59,59}]
  wire  _GEN_54 = 6'h32 == va_line_addr ? meta_50_valid_0 : _GEN_53; // @[ICache.scala 132:{59,59}]
  wire  _GEN_55 = 6'h33 == va_line_addr ? meta_51_valid_0 : _GEN_54; // @[ICache.scala 132:{59,59}]
  wire  _GEN_56 = 6'h34 == va_line_addr ? meta_52_valid_0 : _GEN_55; // @[ICache.scala 132:{59,59}]
  wire  _GEN_57 = 6'h35 == va_line_addr ? meta_53_valid_0 : _GEN_56; // @[ICache.scala 132:{59,59}]
  wire  _GEN_58 = 6'h36 == va_line_addr ? meta_54_valid_0 : _GEN_57; // @[ICache.scala 132:{59,59}]
  wire  _GEN_59 = 6'h37 == va_line_addr ? meta_55_valid_0 : _GEN_58; // @[ICache.scala 132:{59,59}]
  wire  _GEN_60 = 6'h38 == va_line_addr ? meta_56_valid_0 : _GEN_59; // @[ICache.scala 132:{59,59}]
  wire  _GEN_61 = 6'h39 == va_line_addr ? meta_57_valid_0 : _GEN_60; // @[ICache.scala 132:{59,59}]
  wire  _GEN_62 = 6'h3a == va_line_addr ? meta_58_valid_0 : _GEN_61; // @[ICache.scala 132:{59,59}]
  wire  _GEN_63 = 6'h3b == va_line_addr ? meta_59_valid_0 : _GEN_62; // @[ICache.scala 132:{59,59}]
  wire  _GEN_64 = 6'h3c == va_line_addr ? meta_60_valid_0 : _GEN_63; // @[ICache.scala 132:{59,59}]
  wire  _GEN_65 = 6'h3d == va_line_addr ? meta_61_valid_0 : _GEN_64; // @[ICache.scala 132:{59,59}]
  wire  _GEN_66 = 6'h3e == va_line_addr ? meta_62_valid_0 : _GEN_65; // @[ICache.scala 132:{59,59}]
  wire  _GEN_67 = 6'h3f == va_line_addr ? meta_63_valid_0 : _GEN_66; // @[ICache.scala 132:{59,59}]
  wire [6:0] _GEN_13517 = {{1'd0}, va_line_addr}; // @[ICache.scala 132:{59,59}]
  wire  _GEN_68 = 7'h40 == _GEN_13517 ? meta_64_valid_0 : _GEN_67; // @[ICache.scala 132:{59,59}]
  wire  _GEN_69 = 7'h41 == _GEN_13517 ? meta_65_valid_0 : _GEN_68; // @[ICache.scala 132:{59,59}]
  wire  _GEN_70 = 7'h42 == _GEN_13517 ? meta_66_valid_0 : _GEN_69; // @[ICache.scala 132:{59,59}]
  wire  _GEN_71 = 7'h43 == _GEN_13517 ? meta_67_valid_0 : _GEN_70; // @[ICache.scala 132:{59,59}]
  wire  _GEN_72 = 7'h44 == _GEN_13517 ? meta_68_valid_0 : _GEN_71; // @[ICache.scala 132:{59,59}]
  wire  _GEN_73 = 7'h45 == _GEN_13517 ? meta_69_valid_0 : _GEN_72; // @[ICache.scala 132:{59,59}]
  wire  _GEN_74 = 7'h46 == _GEN_13517 ? meta_70_valid_0 : _GEN_73; // @[ICache.scala 132:{59,59}]
  wire  _GEN_75 = 7'h47 == _GEN_13517 ? meta_71_valid_0 : _GEN_74; // @[ICache.scala 132:{59,59}]
  wire  _GEN_76 = 7'h48 == _GEN_13517 ? meta_72_valid_0 : _GEN_75; // @[ICache.scala 132:{59,59}]
  wire  _GEN_77 = 7'h49 == _GEN_13517 ? meta_73_valid_0 : _GEN_76; // @[ICache.scala 132:{59,59}]
  wire  _GEN_78 = 7'h4a == _GEN_13517 ? meta_74_valid_0 : _GEN_77; // @[ICache.scala 132:{59,59}]
  wire  _GEN_79 = 7'h4b == _GEN_13517 ? meta_75_valid_0 : _GEN_78; // @[ICache.scala 132:{59,59}]
  wire  _GEN_80 = 7'h4c == _GEN_13517 ? meta_76_valid_0 : _GEN_79; // @[ICache.scala 132:{59,59}]
  wire  _GEN_81 = 7'h4d == _GEN_13517 ? meta_77_valid_0 : _GEN_80; // @[ICache.scala 132:{59,59}]
  wire  _GEN_82 = 7'h4e == _GEN_13517 ? meta_78_valid_0 : _GEN_81; // @[ICache.scala 132:{59,59}]
  wire  _GEN_83 = 7'h4f == _GEN_13517 ? meta_79_valid_0 : _GEN_82; // @[ICache.scala 132:{59,59}]
  wire  _GEN_84 = 7'h50 == _GEN_13517 ? meta_80_valid_0 : _GEN_83; // @[ICache.scala 132:{59,59}]
  wire  _GEN_85 = 7'h51 == _GEN_13517 ? meta_81_valid_0 : _GEN_84; // @[ICache.scala 132:{59,59}]
  wire  _GEN_86 = 7'h52 == _GEN_13517 ? meta_82_valid_0 : _GEN_85; // @[ICache.scala 132:{59,59}]
  wire  _GEN_87 = 7'h53 == _GEN_13517 ? meta_83_valid_0 : _GEN_86; // @[ICache.scala 132:{59,59}]
  wire  _GEN_88 = 7'h54 == _GEN_13517 ? meta_84_valid_0 : _GEN_87; // @[ICache.scala 132:{59,59}]
  wire  _GEN_89 = 7'h55 == _GEN_13517 ? meta_85_valid_0 : _GEN_88; // @[ICache.scala 132:{59,59}]
  wire  _GEN_90 = 7'h56 == _GEN_13517 ? meta_86_valid_0 : _GEN_89; // @[ICache.scala 132:{59,59}]
  wire  _GEN_91 = 7'h57 == _GEN_13517 ? meta_87_valid_0 : _GEN_90; // @[ICache.scala 132:{59,59}]
  wire  _GEN_92 = 7'h58 == _GEN_13517 ? meta_88_valid_0 : _GEN_91; // @[ICache.scala 132:{59,59}]
  wire  _GEN_93 = 7'h59 == _GEN_13517 ? meta_89_valid_0 : _GEN_92; // @[ICache.scala 132:{59,59}]
  wire  _GEN_94 = 7'h5a == _GEN_13517 ? meta_90_valid_0 : _GEN_93; // @[ICache.scala 132:{59,59}]
  wire  _GEN_95 = 7'h5b == _GEN_13517 ? meta_91_valid_0 : _GEN_94; // @[ICache.scala 132:{59,59}]
  wire  _GEN_96 = 7'h5c == _GEN_13517 ? meta_92_valid_0 : _GEN_95; // @[ICache.scala 132:{59,59}]
  wire  _GEN_97 = 7'h5d == _GEN_13517 ? meta_93_valid_0 : _GEN_96; // @[ICache.scala 132:{59,59}]
  wire  _GEN_98 = 7'h5e == _GEN_13517 ? meta_94_valid_0 : _GEN_97; // @[ICache.scala 132:{59,59}]
  wire  _GEN_99 = 7'h5f == _GEN_13517 ? meta_95_valid_0 : _GEN_98; // @[ICache.scala 132:{59,59}]
  wire  _GEN_100 = 7'h60 == _GEN_13517 ? meta_96_valid_0 : _GEN_99; // @[ICache.scala 132:{59,59}]
  wire  _GEN_101 = 7'h61 == _GEN_13517 ? meta_97_valid_0 : _GEN_100; // @[ICache.scala 132:{59,59}]
  wire  _GEN_102 = 7'h62 == _GEN_13517 ? meta_98_valid_0 : _GEN_101; // @[ICache.scala 132:{59,59}]
  wire  _GEN_103 = 7'h63 == _GEN_13517 ? meta_99_valid_0 : _GEN_102; // @[ICache.scala 132:{59,59}]
  wire  _GEN_104 = 7'h64 == _GEN_13517 ? meta_100_valid_0 : _GEN_103; // @[ICache.scala 132:{59,59}]
  wire  _GEN_105 = 7'h65 == _GEN_13517 ? meta_101_valid_0 : _GEN_104; // @[ICache.scala 132:{59,59}]
  wire  _GEN_106 = 7'h66 == _GEN_13517 ? meta_102_valid_0 : _GEN_105; // @[ICache.scala 132:{59,59}]
  wire  _GEN_107 = 7'h67 == _GEN_13517 ? meta_103_valid_0 : _GEN_106; // @[ICache.scala 132:{59,59}]
  wire  _GEN_108 = 7'h68 == _GEN_13517 ? meta_104_valid_0 : _GEN_107; // @[ICache.scala 132:{59,59}]
  wire  _GEN_109 = 7'h69 == _GEN_13517 ? meta_105_valid_0 : _GEN_108; // @[ICache.scala 132:{59,59}]
  wire  _GEN_110 = 7'h6a == _GEN_13517 ? meta_106_valid_0 : _GEN_109; // @[ICache.scala 132:{59,59}]
  wire  _GEN_111 = 7'h6b == _GEN_13517 ? meta_107_valid_0 : _GEN_110; // @[ICache.scala 132:{59,59}]
  wire  _GEN_112 = 7'h6c == _GEN_13517 ? meta_108_valid_0 : _GEN_111; // @[ICache.scala 132:{59,59}]
  wire  _GEN_113 = 7'h6d == _GEN_13517 ? meta_109_valid_0 : _GEN_112; // @[ICache.scala 132:{59,59}]
  wire  _GEN_114 = 7'h6e == _GEN_13517 ? meta_110_valid_0 : _GEN_113; // @[ICache.scala 132:{59,59}]
  wire  _GEN_115 = 7'h6f == _GEN_13517 ? meta_111_valid_0 : _GEN_114; // @[ICache.scala 132:{59,59}]
  wire  _GEN_116 = 7'h70 == _GEN_13517 ? meta_112_valid_0 : _GEN_115; // @[ICache.scala 132:{59,59}]
  wire  _GEN_117 = 7'h71 == _GEN_13517 ? meta_113_valid_0 : _GEN_116; // @[ICache.scala 132:{59,59}]
  wire  _GEN_118 = 7'h72 == _GEN_13517 ? meta_114_valid_0 : _GEN_117; // @[ICache.scala 132:{59,59}]
  wire  _GEN_119 = 7'h73 == _GEN_13517 ? meta_115_valid_0 : _GEN_118; // @[ICache.scala 132:{59,59}]
  wire  _GEN_120 = 7'h74 == _GEN_13517 ? meta_116_valid_0 : _GEN_119; // @[ICache.scala 132:{59,59}]
  wire  _GEN_121 = 7'h75 == _GEN_13517 ? meta_117_valid_0 : _GEN_120; // @[ICache.scala 132:{59,59}]
  wire  _GEN_122 = 7'h76 == _GEN_13517 ? meta_118_valid_0 : _GEN_121; // @[ICache.scala 132:{59,59}]
  wire  _GEN_123 = 7'h77 == _GEN_13517 ? meta_119_valid_0 : _GEN_122; // @[ICache.scala 132:{59,59}]
  wire  _GEN_124 = 7'h78 == _GEN_13517 ? meta_120_valid_0 : _GEN_123; // @[ICache.scala 132:{59,59}]
  wire  _GEN_125 = 7'h79 == _GEN_13517 ? meta_121_valid_0 : _GEN_124; // @[ICache.scala 132:{59,59}]
  wire  _GEN_126 = 7'h7a == _GEN_13517 ? meta_122_valid_0 : _GEN_125; // @[ICache.scala 132:{59,59}]
  wire  _GEN_127 = 7'h7b == _GEN_13517 ? meta_123_valid_0 : _GEN_126; // @[ICache.scala 132:{59,59}]
  wire  _GEN_128 = 7'h7c == _GEN_13517 ? meta_124_valid_0 : _GEN_127; // @[ICache.scala 132:{59,59}]
  wire  _GEN_129 = 7'h7d == _GEN_13517 ? meta_125_valid_0 : _GEN_128; // @[ICache.scala 132:{59,59}]
  wire  _GEN_130 = 7'h7e == _GEN_13517 ? meta_126_valid_0 : _GEN_129; // @[ICache.scala 132:{59,59}]
  wire  _GEN_131 = 7'h7f == _GEN_13517 ? meta_127_valid_0 : _GEN_130; // @[ICache.scala 132:{59,59}]
  wire [7:0] _GEN_13581 = {{2'd0}, va_line_addr}; // @[ICache.scala 132:{59,59}]
  wire  _GEN_132 = 8'h80 == _GEN_13581 ? meta_128_valid_0 : _GEN_131; // @[ICache.scala 132:{59,59}]
  wire  _GEN_133 = 8'h81 == _GEN_13581 ? meta_129_valid_0 : _GEN_132; // @[ICache.scala 132:{59,59}]
  wire  _GEN_134 = 8'h82 == _GEN_13581 ? meta_130_valid_0 : _GEN_133; // @[ICache.scala 132:{59,59}]
  wire  _GEN_135 = 8'h83 == _GEN_13581 ? meta_131_valid_0 : _GEN_134; // @[ICache.scala 132:{59,59}]
  wire  _GEN_136 = 8'h84 == _GEN_13581 ? meta_132_valid_0 : _GEN_135; // @[ICache.scala 132:{59,59}]
  wire  _GEN_137 = 8'h85 == _GEN_13581 ? meta_133_valid_0 : _GEN_136; // @[ICache.scala 132:{59,59}]
  wire  _GEN_138 = 8'h86 == _GEN_13581 ? meta_134_valid_0 : _GEN_137; // @[ICache.scala 132:{59,59}]
  wire  _GEN_139 = 8'h87 == _GEN_13581 ? meta_135_valid_0 : _GEN_138; // @[ICache.scala 132:{59,59}]
  wire  _GEN_140 = 8'h88 == _GEN_13581 ? meta_136_valid_0 : _GEN_139; // @[ICache.scala 132:{59,59}]
  wire  _GEN_141 = 8'h89 == _GEN_13581 ? meta_137_valid_0 : _GEN_140; // @[ICache.scala 132:{59,59}]
  wire  _GEN_142 = 8'h8a == _GEN_13581 ? meta_138_valid_0 : _GEN_141; // @[ICache.scala 132:{59,59}]
  wire  _GEN_143 = 8'h8b == _GEN_13581 ? meta_139_valid_0 : _GEN_142; // @[ICache.scala 132:{59,59}]
  wire  _GEN_144 = 8'h8c == _GEN_13581 ? meta_140_valid_0 : _GEN_143; // @[ICache.scala 132:{59,59}]
  wire  _GEN_145 = 8'h8d == _GEN_13581 ? meta_141_valid_0 : _GEN_144; // @[ICache.scala 132:{59,59}]
  wire  _GEN_146 = 8'h8e == _GEN_13581 ? meta_142_valid_0 : _GEN_145; // @[ICache.scala 132:{59,59}]
  wire  _GEN_147 = 8'h8f == _GEN_13581 ? meta_143_valid_0 : _GEN_146; // @[ICache.scala 132:{59,59}]
  wire  _GEN_148 = 8'h90 == _GEN_13581 ? meta_144_valid_0 : _GEN_147; // @[ICache.scala 132:{59,59}]
  wire  _GEN_149 = 8'h91 == _GEN_13581 ? meta_145_valid_0 : _GEN_148; // @[ICache.scala 132:{59,59}]
  wire  _GEN_150 = 8'h92 == _GEN_13581 ? meta_146_valid_0 : _GEN_149; // @[ICache.scala 132:{59,59}]
  wire  _GEN_151 = 8'h93 == _GEN_13581 ? meta_147_valid_0 : _GEN_150; // @[ICache.scala 132:{59,59}]
  wire  _GEN_152 = 8'h94 == _GEN_13581 ? meta_148_valid_0 : _GEN_151; // @[ICache.scala 132:{59,59}]
  wire  _GEN_153 = 8'h95 == _GEN_13581 ? meta_149_valid_0 : _GEN_152; // @[ICache.scala 132:{59,59}]
  wire  _GEN_154 = 8'h96 == _GEN_13581 ? meta_150_valid_0 : _GEN_153; // @[ICache.scala 132:{59,59}]
  wire  _GEN_155 = 8'h97 == _GEN_13581 ? meta_151_valid_0 : _GEN_154; // @[ICache.scala 132:{59,59}]
  wire  _GEN_156 = 8'h98 == _GEN_13581 ? meta_152_valid_0 : _GEN_155; // @[ICache.scala 132:{59,59}]
  wire  _GEN_157 = 8'h99 == _GEN_13581 ? meta_153_valid_0 : _GEN_156; // @[ICache.scala 132:{59,59}]
  wire  _GEN_158 = 8'h9a == _GEN_13581 ? meta_154_valid_0 : _GEN_157; // @[ICache.scala 132:{59,59}]
  wire  _GEN_159 = 8'h9b == _GEN_13581 ? meta_155_valid_0 : _GEN_158; // @[ICache.scala 132:{59,59}]
  wire  _GEN_160 = 8'h9c == _GEN_13581 ? meta_156_valid_0 : _GEN_159; // @[ICache.scala 132:{59,59}]
  wire  _GEN_161 = 8'h9d == _GEN_13581 ? meta_157_valid_0 : _GEN_160; // @[ICache.scala 132:{59,59}]
  wire  _GEN_162 = 8'h9e == _GEN_13581 ? meta_158_valid_0 : _GEN_161; // @[ICache.scala 132:{59,59}]
  wire  _GEN_163 = 8'h9f == _GEN_13581 ? meta_159_valid_0 : _GEN_162; // @[ICache.scala 132:{59,59}]
  wire  _GEN_164 = 8'ha0 == _GEN_13581 ? meta_160_valid_0 : _GEN_163; // @[ICache.scala 132:{59,59}]
  wire  _GEN_165 = 8'ha1 == _GEN_13581 ? meta_161_valid_0 : _GEN_164; // @[ICache.scala 132:{59,59}]
  wire  _GEN_166 = 8'ha2 == _GEN_13581 ? meta_162_valid_0 : _GEN_165; // @[ICache.scala 132:{59,59}]
  wire  _GEN_167 = 8'ha3 == _GEN_13581 ? meta_163_valid_0 : _GEN_166; // @[ICache.scala 132:{59,59}]
  wire  _GEN_168 = 8'ha4 == _GEN_13581 ? meta_164_valid_0 : _GEN_167; // @[ICache.scala 132:{59,59}]
  wire  _GEN_169 = 8'ha5 == _GEN_13581 ? meta_165_valid_0 : _GEN_168; // @[ICache.scala 132:{59,59}]
  wire  _GEN_170 = 8'ha6 == _GEN_13581 ? meta_166_valid_0 : _GEN_169; // @[ICache.scala 132:{59,59}]
  wire  _GEN_171 = 8'ha7 == _GEN_13581 ? meta_167_valid_0 : _GEN_170; // @[ICache.scala 132:{59,59}]
  wire  _GEN_172 = 8'ha8 == _GEN_13581 ? meta_168_valid_0 : _GEN_171; // @[ICache.scala 132:{59,59}]
  wire  _GEN_173 = 8'ha9 == _GEN_13581 ? meta_169_valid_0 : _GEN_172; // @[ICache.scala 132:{59,59}]
  wire  _GEN_174 = 8'haa == _GEN_13581 ? meta_170_valid_0 : _GEN_173; // @[ICache.scala 132:{59,59}]
  wire  _GEN_175 = 8'hab == _GEN_13581 ? meta_171_valid_0 : _GEN_174; // @[ICache.scala 132:{59,59}]
  wire  _GEN_176 = 8'hac == _GEN_13581 ? meta_172_valid_0 : _GEN_175; // @[ICache.scala 132:{59,59}]
  wire  _GEN_177 = 8'had == _GEN_13581 ? meta_173_valid_0 : _GEN_176; // @[ICache.scala 132:{59,59}]
  wire  _GEN_178 = 8'hae == _GEN_13581 ? meta_174_valid_0 : _GEN_177; // @[ICache.scala 132:{59,59}]
  wire  _GEN_179 = 8'haf == _GEN_13581 ? meta_175_valid_0 : _GEN_178; // @[ICache.scala 132:{59,59}]
  wire  _GEN_180 = 8'hb0 == _GEN_13581 ? meta_176_valid_0 : _GEN_179; // @[ICache.scala 132:{59,59}]
  wire  _GEN_181 = 8'hb1 == _GEN_13581 ? meta_177_valid_0 : _GEN_180; // @[ICache.scala 132:{59,59}]
  wire  _GEN_182 = 8'hb2 == _GEN_13581 ? meta_178_valid_0 : _GEN_181; // @[ICache.scala 132:{59,59}]
  wire  _GEN_183 = 8'hb3 == _GEN_13581 ? meta_179_valid_0 : _GEN_182; // @[ICache.scala 132:{59,59}]
  wire  _GEN_184 = 8'hb4 == _GEN_13581 ? meta_180_valid_0 : _GEN_183; // @[ICache.scala 132:{59,59}]
  wire  _GEN_185 = 8'hb5 == _GEN_13581 ? meta_181_valid_0 : _GEN_184; // @[ICache.scala 132:{59,59}]
  wire  _GEN_186 = 8'hb6 == _GEN_13581 ? meta_182_valid_0 : _GEN_185; // @[ICache.scala 132:{59,59}]
  wire  _GEN_187 = 8'hb7 == _GEN_13581 ? meta_183_valid_0 : _GEN_186; // @[ICache.scala 132:{59,59}]
  wire  _GEN_188 = 8'hb8 == _GEN_13581 ? meta_184_valid_0 : _GEN_187; // @[ICache.scala 132:{59,59}]
  wire  _GEN_189 = 8'hb9 == _GEN_13581 ? meta_185_valid_0 : _GEN_188; // @[ICache.scala 132:{59,59}]
  wire  _GEN_190 = 8'hba == _GEN_13581 ? meta_186_valid_0 : _GEN_189; // @[ICache.scala 132:{59,59}]
  wire  _GEN_191 = 8'hbb == _GEN_13581 ? meta_187_valid_0 : _GEN_190; // @[ICache.scala 132:{59,59}]
  wire  _GEN_192 = 8'hbc == _GEN_13581 ? meta_188_valid_0 : _GEN_191; // @[ICache.scala 132:{59,59}]
  wire  _GEN_193 = 8'hbd == _GEN_13581 ? meta_189_valid_0 : _GEN_192; // @[ICache.scala 132:{59,59}]
  wire  _GEN_194 = 8'hbe == _GEN_13581 ? meta_190_valid_0 : _GEN_193; // @[ICache.scala 132:{59,59}]
  wire  _GEN_195 = 8'hbf == _GEN_13581 ? meta_191_valid_0 : _GEN_194; // @[ICache.scala 132:{59,59}]
  wire  _GEN_196 = 8'hc0 == _GEN_13581 ? meta_192_valid_0 : _GEN_195; // @[ICache.scala 132:{59,59}]
  wire  _GEN_197 = 8'hc1 == _GEN_13581 ? meta_193_valid_0 : _GEN_196; // @[ICache.scala 132:{59,59}]
  wire  _GEN_198 = 8'hc2 == _GEN_13581 ? meta_194_valid_0 : _GEN_197; // @[ICache.scala 132:{59,59}]
  wire  _GEN_199 = 8'hc3 == _GEN_13581 ? meta_195_valid_0 : _GEN_198; // @[ICache.scala 132:{59,59}]
  wire  _GEN_200 = 8'hc4 == _GEN_13581 ? meta_196_valid_0 : _GEN_199; // @[ICache.scala 132:{59,59}]
  wire  _GEN_201 = 8'hc5 == _GEN_13581 ? meta_197_valid_0 : _GEN_200; // @[ICache.scala 132:{59,59}]
  wire  _GEN_202 = 8'hc6 == _GEN_13581 ? meta_198_valid_0 : _GEN_201; // @[ICache.scala 132:{59,59}]
  wire  _GEN_203 = 8'hc7 == _GEN_13581 ? meta_199_valid_0 : _GEN_202; // @[ICache.scala 132:{59,59}]
  wire  _GEN_204 = 8'hc8 == _GEN_13581 ? meta_200_valid_0 : _GEN_203; // @[ICache.scala 132:{59,59}]
  wire  _GEN_205 = 8'hc9 == _GEN_13581 ? meta_201_valid_0 : _GEN_204; // @[ICache.scala 132:{59,59}]
  wire  _GEN_206 = 8'hca == _GEN_13581 ? meta_202_valid_0 : _GEN_205; // @[ICache.scala 132:{59,59}]
  wire  _GEN_207 = 8'hcb == _GEN_13581 ? meta_203_valid_0 : _GEN_206; // @[ICache.scala 132:{59,59}]
  wire  _GEN_208 = 8'hcc == _GEN_13581 ? meta_204_valid_0 : _GEN_207; // @[ICache.scala 132:{59,59}]
  wire  _GEN_209 = 8'hcd == _GEN_13581 ? meta_205_valid_0 : _GEN_208; // @[ICache.scala 132:{59,59}]
  wire  _GEN_210 = 8'hce == _GEN_13581 ? meta_206_valid_0 : _GEN_209; // @[ICache.scala 132:{59,59}]
  wire  _GEN_211 = 8'hcf == _GEN_13581 ? meta_207_valid_0 : _GEN_210; // @[ICache.scala 132:{59,59}]
  wire  _GEN_212 = 8'hd0 == _GEN_13581 ? meta_208_valid_0 : _GEN_211; // @[ICache.scala 132:{59,59}]
  wire  _GEN_213 = 8'hd1 == _GEN_13581 ? meta_209_valid_0 : _GEN_212; // @[ICache.scala 132:{59,59}]
  wire  _GEN_214 = 8'hd2 == _GEN_13581 ? meta_210_valid_0 : _GEN_213; // @[ICache.scala 132:{59,59}]
  wire  _GEN_215 = 8'hd3 == _GEN_13581 ? meta_211_valid_0 : _GEN_214; // @[ICache.scala 132:{59,59}]
  wire  _GEN_216 = 8'hd4 == _GEN_13581 ? meta_212_valid_0 : _GEN_215; // @[ICache.scala 132:{59,59}]
  wire  _GEN_217 = 8'hd5 == _GEN_13581 ? meta_213_valid_0 : _GEN_216; // @[ICache.scala 132:{59,59}]
  wire  _GEN_218 = 8'hd6 == _GEN_13581 ? meta_214_valid_0 : _GEN_217; // @[ICache.scala 132:{59,59}]
  wire  _GEN_219 = 8'hd7 == _GEN_13581 ? meta_215_valid_0 : _GEN_218; // @[ICache.scala 132:{59,59}]
  wire  _GEN_220 = 8'hd8 == _GEN_13581 ? meta_216_valid_0 : _GEN_219; // @[ICache.scala 132:{59,59}]
  wire  _GEN_221 = 8'hd9 == _GEN_13581 ? meta_217_valid_0 : _GEN_220; // @[ICache.scala 132:{59,59}]
  wire  _GEN_222 = 8'hda == _GEN_13581 ? meta_218_valid_0 : _GEN_221; // @[ICache.scala 132:{59,59}]
  wire  _GEN_223 = 8'hdb == _GEN_13581 ? meta_219_valid_0 : _GEN_222; // @[ICache.scala 132:{59,59}]
  wire  _GEN_224 = 8'hdc == _GEN_13581 ? meta_220_valid_0 : _GEN_223; // @[ICache.scala 132:{59,59}]
  wire  _GEN_225 = 8'hdd == _GEN_13581 ? meta_221_valid_0 : _GEN_224; // @[ICache.scala 132:{59,59}]
  wire  _GEN_226 = 8'hde == _GEN_13581 ? meta_222_valid_0 : _GEN_225; // @[ICache.scala 132:{59,59}]
  wire  _GEN_227 = 8'hdf == _GEN_13581 ? meta_223_valid_0 : _GEN_226; // @[ICache.scala 132:{59,59}]
  wire  _GEN_228 = 8'he0 == _GEN_13581 ? meta_224_valid_0 : _GEN_227; // @[ICache.scala 132:{59,59}]
  wire  _GEN_229 = 8'he1 == _GEN_13581 ? meta_225_valid_0 : _GEN_228; // @[ICache.scala 132:{59,59}]
  wire  _GEN_230 = 8'he2 == _GEN_13581 ? meta_226_valid_0 : _GEN_229; // @[ICache.scala 132:{59,59}]
  wire  _GEN_231 = 8'he3 == _GEN_13581 ? meta_227_valid_0 : _GEN_230; // @[ICache.scala 132:{59,59}]
  wire  _GEN_232 = 8'he4 == _GEN_13581 ? meta_228_valid_0 : _GEN_231; // @[ICache.scala 132:{59,59}]
  wire  _GEN_233 = 8'he5 == _GEN_13581 ? meta_229_valid_0 : _GEN_232; // @[ICache.scala 132:{59,59}]
  wire  _GEN_234 = 8'he6 == _GEN_13581 ? meta_230_valid_0 : _GEN_233; // @[ICache.scala 132:{59,59}]
  wire  _GEN_235 = 8'he7 == _GEN_13581 ? meta_231_valid_0 : _GEN_234; // @[ICache.scala 132:{59,59}]
  wire  _GEN_236 = 8'he8 == _GEN_13581 ? meta_232_valid_0 : _GEN_235; // @[ICache.scala 132:{59,59}]
  wire  _GEN_237 = 8'he9 == _GEN_13581 ? meta_233_valid_0 : _GEN_236; // @[ICache.scala 132:{59,59}]
  wire  _GEN_238 = 8'hea == _GEN_13581 ? meta_234_valid_0 : _GEN_237; // @[ICache.scala 132:{59,59}]
  wire  _GEN_239 = 8'heb == _GEN_13581 ? meta_235_valid_0 : _GEN_238; // @[ICache.scala 132:{59,59}]
  wire  _GEN_240 = 8'hec == _GEN_13581 ? meta_236_valid_0 : _GEN_239; // @[ICache.scala 132:{59,59}]
  wire  _GEN_241 = 8'hed == _GEN_13581 ? meta_237_valid_0 : _GEN_240; // @[ICache.scala 132:{59,59}]
  wire  _GEN_242 = 8'hee == _GEN_13581 ? meta_238_valid_0 : _GEN_241; // @[ICache.scala 132:{59,59}]
  wire  _GEN_243 = 8'hef == _GEN_13581 ? meta_239_valid_0 : _GEN_242; // @[ICache.scala 132:{59,59}]
  wire  _GEN_244 = 8'hf0 == _GEN_13581 ? meta_240_valid_0 : _GEN_243; // @[ICache.scala 132:{59,59}]
  wire  _GEN_245 = 8'hf1 == _GEN_13581 ? meta_241_valid_0 : _GEN_244; // @[ICache.scala 132:{59,59}]
  wire  _GEN_246 = 8'hf2 == _GEN_13581 ? meta_242_valid_0 : _GEN_245; // @[ICache.scala 132:{59,59}]
  wire  _GEN_247 = 8'hf3 == _GEN_13581 ? meta_243_valid_0 : _GEN_246; // @[ICache.scala 132:{59,59}]
  wire  _GEN_248 = 8'hf4 == _GEN_13581 ? meta_244_valid_0 : _GEN_247; // @[ICache.scala 132:{59,59}]
  wire  _GEN_249 = 8'hf5 == _GEN_13581 ? meta_245_valid_0 : _GEN_248; // @[ICache.scala 132:{59,59}]
  wire  _GEN_250 = 8'hf6 == _GEN_13581 ? meta_246_valid_0 : _GEN_249; // @[ICache.scala 132:{59,59}]
  wire  _GEN_251 = 8'hf7 == _GEN_13581 ? meta_247_valid_0 : _GEN_250; // @[ICache.scala 132:{59,59}]
  wire  _GEN_252 = 8'hf8 == _GEN_13581 ? meta_248_valid_0 : _GEN_251; // @[ICache.scala 132:{59,59}]
  wire  _GEN_253 = 8'hf9 == _GEN_13581 ? meta_249_valid_0 : _GEN_252; // @[ICache.scala 132:{59,59}]
  wire  _GEN_254 = 8'hfa == _GEN_13581 ? meta_250_valid_0 : _GEN_253; // @[ICache.scala 132:{59,59}]
  wire  _GEN_255 = 8'hfb == _GEN_13581 ? meta_251_valid_0 : _GEN_254; // @[ICache.scala 132:{59,59}]
  wire  _GEN_256 = 8'hfc == _GEN_13581 ? meta_252_valid_0 : _GEN_255; // @[ICache.scala 132:{59,59}]
  wire  _GEN_257 = 8'hfd == _GEN_13581 ? meta_253_valid_0 : _GEN_256; // @[ICache.scala 132:{59,59}]
  wire  _GEN_258 = 8'hfe == _GEN_13581 ? meta_254_valid_0 : _GEN_257; // @[ICache.scala 132:{59,59}]
  wire  _GEN_259 = 8'hff == _GEN_13581 ? meta_255_valid_0 : _GEN_258; // @[ICache.scala 132:{59,59}]
  wire [8:0] _GEN_13709 = {{3'd0}, va_line_addr}; // @[ICache.scala 132:{59,59}]
  wire  _GEN_260 = 9'h100 == _GEN_13709 ? meta_256_valid_0 : _GEN_259; // @[ICache.scala 132:{59,59}]
  wire  _GEN_261 = 9'h101 == _GEN_13709 ? meta_257_valid_0 : _GEN_260; // @[ICache.scala 132:{59,59}]
  wire  _GEN_262 = 9'h102 == _GEN_13709 ? meta_258_valid_0 : _GEN_261; // @[ICache.scala 132:{59,59}]
  wire  _GEN_263 = 9'h103 == _GEN_13709 ? meta_259_valid_0 : _GEN_262; // @[ICache.scala 132:{59,59}]
  wire  _GEN_264 = 9'h104 == _GEN_13709 ? meta_260_valid_0 : _GEN_263; // @[ICache.scala 132:{59,59}]
  wire  _GEN_265 = 9'h105 == _GEN_13709 ? meta_261_valid_0 : _GEN_264; // @[ICache.scala 132:{59,59}]
  wire  _GEN_266 = 9'h106 == _GEN_13709 ? meta_262_valid_0 : _GEN_265; // @[ICache.scala 132:{59,59}]
  wire  _GEN_267 = 9'h107 == _GEN_13709 ? meta_263_valid_0 : _GEN_266; // @[ICache.scala 132:{59,59}]
  wire  _GEN_268 = 9'h108 == _GEN_13709 ? meta_264_valid_0 : _GEN_267; // @[ICache.scala 132:{59,59}]
  wire  _GEN_269 = 9'h109 == _GEN_13709 ? meta_265_valid_0 : _GEN_268; // @[ICache.scala 132:{59,59}]
  wire  _GEN_270 = 9'h10a == _GEN_13709 ? meta_266_valid_0 : _GEN_269; // @[ICache.scala 132:{59,59}]
  wire  _GEN_271 = 9'h10b == _GEN_13709 ? meta_267_valid_0 : _GEN_270; // @[ICache.scala 132:{59,59}]
  wire  _GEN_272 = 9'h10c == _GEN_13709 ? meta_268_valid_0 : _GEN_271; // @[ICache.scala 132:{59,59}]
  wire  _GEN_273 = 9'h10d == _GEN_13709 ? meta_269_valid_0 : _GEN_272; // @[ICache.scala 132:{59,59}]
  wire  _GEN_274 = 9'h10e == _GEN_13709 ? meta_270_valid_0 : _GEN_273; // @[ICache.scala 132:{59,59}]
  wire  _GEN_275 = 9'h10f == _GEN_13709 ? meta_271_valid_0 : _GEN_274; // @[ICache.scala 132:{59,59}]
  wire  _GEN_276 = 9'h110 == _GEN_13709 ? meta_272_valid_0 : _GEN_275; // @[ICache.scala 132:{59,59}]
  wire  _GEN_277 = 9'h111 == _GEN_13709 ? meta_273_valid_0 : _GEN_276; // @[ICache.scala 132:{59,59}]
  wire  _GEN_278 = 9'h112 == _GEN_13709 ? meta_274_valid_0 : _GEN_277; // @[ICache.scala 132:{59,59}]
  wire  _GEN_279 = 9'h113 == _GEN_13709 ? meta_275_valid_0 : _GEN_278; // @[ICache.scala 132:{59,59}]
  wire  _GEN_280 = 9'h114 == _GEN_13709 ? meta_276_valid_0 : _GEN_279; // @[ICache.scala 132:{59,59}]
  wire  _GEN_281 = 9'h115 == _GEN_13709 ? meta_277_valid_0 : _GEN_280; // @[ICache.scala 132:{59,59}]
  wire  _GEN_282 = 9'h116 == _GEN_13709 ? meta_278_valid_0 : _GEN_281; // @[ICache.scala 132:{59,59}]
  wire  _GEN_283 = 9'h117 == _GEN_13709 ? meta_279_valid_0 : _GEN_282; // @[ICache.scala 132:{59,59}]
  wire  _GEN_284 = 9'h118 == _GEN_13709 ? meta_280_valid_0 : _GEN_283; // @[ICache.scala 132:{59,59}]
  wire  _GEN_285 = 9'h119 == _GEN_13709 ? meta_281_valid_0 : _GEN_284; // @[ICache.scala 132:{59,59}]
  wire  _GEN_286 = 9'h11a == _GEN_13709 ? meta_282_valid_0 : _GEN_285; // @[ICache.scala 132:{59,59}]
  wire  _GEN_287 = 9'h11b == _GEN_13709 ? meta_283_valid_0 : _GEN_286; // @[ICache.scala 132:{59,59}]
  wire  _GEN_288 = 9'h11c == _GEN_13709 ? meta_284_valid_0 : _GEN_287; // @[ICache.scala 132:{59,59}]
  wire  _GEN_289 = 9'h11d == _GEN_13709 ? meta_285_valid_0 : _GEN_288; // @[ICache.scala 132:{59,59}]
  wire  _GEN_290 = 9'h11e == _GEN_13709 ? meta_286_valid_0 : _GEN_289; // @[ICache.scala 132:{59,59}]
  wire  _GEN_291 = 9'h11f == _GEN_13709 ? meta_287_valid_0 : _GEN_290; // @[ICache.scala 132:{59,59}]
  wire  _GEN_292 = 9'h120 == _GEN_13709 ? meta_288_valid_0 : _GEN_291; // @[ICache.scala 132:{59,59}]
  wire  _GEN_293 = 9'h121 == _GEN_13709 ? meta_289_valid_0 : _GEN_292; // @[ICache.scala 132:{59,59}]
  wire  _GEN_294 = 9'h122 == _GEN_13709 ? meta_290_valid_0 : _GEN_293; // @[ICache.scala 132:{59,59}]
  wire  _GEN_295 = 9'h123 == _GEN_13709 ? meta_291_valid_0 : _GEN_294; // @[ICache.scala 132:{59,59}]
  wire  _GEN_296 = 9'h124 == _GEN_13709 ? meta_292_valid_0 : _GEN_295; // @[ICache.scala 132:{59,59}]
  wire  _GEN_297 = 9'h125 == _GEN_13709 ? meta_293_valid_0 : _GEN_296; // @[ICache.scala 132:{59,59}]
  wire  _GEN_298 = 9'h126 == _GEN_13709 ? meta_294_valid_0 : _GEN_297; // @[ICache.scala 132:{59,59}]
  wire  _GEN_299 = 9'h127 == _GEN_13709 ? meta_295_valid_0 : _GEN_298; // @[ICache.scala 132:{59,59}]
  wire  _GEN_300 = 9'h128 == _GEN_13709 ? meta_296_valid_0 : _GEN_299; // @[ICache.scala 132:{59,59}]
  wire  _GEN_301 = 9'h129 == _GEN_13709 ? meta_297_valid_0 : _GEN_300; // @[ICache.scala 132:{59,59}]
  wire  _GEN_302 = 9'h12a == _GEN_13709 ? meta_298_valid_0 : _GEN_301; // @[ICache.scala 132:{59,59}]
  wire  _GEN_303 = 9'h12b == _GEN_13709 ? meta_299_valid_0 : _GEN_302; // @[ICache.scala 132:{59,59}]
  wire  _GEN_304 = 9'h12c == _GEN_13709 ? meta_300_valid_0 : _GEN_303; // @[ICache.scala 132:{59,59}]
  wire  _GEN_305 = 9'h12d == _GEN_13709 ? meta_301_valid_0 : _GEN_304; // @[ICache.scala 132:{59,59}]
  wire  _GEN_306 = 9'h12e == _GEN_13709 ? meta_302_valid_0 : _GEN_305; // @[ICache.scala 132:{59,59}]
  wire  _GEN_307 = 9'h12f == _GEN_13709 ? meta_303_valid_0 : _GEN_306; // @[ICache.scala 132:{59,59}]
  wire  _GEN_308 = 9'h130 == _GEN_13709 ? meta_304_valid_0 : _GEN_307; // @[ICache.scala 132:{59,59}]
  wire  _GEN_309 = 9'h131 == _GEN_13709 ? meta_305_valid_0 : _GEN_308; // @[ICache.scala 132:{59,59}]
  wire  _GEN_310 = 9'h132 == _GEN_13709 ? meta_306_valid_0 : _GEN_309; // @[ICache.scala 132:{59,59}]
  wire  _GEN_311 = 9'h133 == _GEN_13709 ? meta_307_valid_0 : _GEN_310; // @[ICache.scala 132:{59,59}]
  wire  _GEN_312 = 9'h134 == _GEN_13709 ? meta_308_valid_0 : _GEN_311; // @[ICache.scala 132:{59,59}]
  wire  _GEN_313 = 9'h135 == _GEN_13709 ? meta_309_valid_0 : _GEN_312; // @[ICache.scala 132:{59,59}]
  wire  _GEN_314 = 9'h136 == _GEN_13709 ? meta_310_valid_0 : _GEN_313; // @[ICache.scala 132:{59,59}]
  wire  _GEN_315 = 9'h137 == _GEN_13709 ? meta_311_valid_0 : _GEN_314; // @[ICache.scala 132:{59,59}]
  wire  _GEN_316 = 9'h138 == _GEN_13709 ? meta_312_valid_0 : _GEN_315; // @[ICache.scala 132:{59,59}]
  wire  _GEN_317 = 9'h139 == _GEN_13709 ? meta_313_valid_0 : _GEN_316; // @[ICache.scala 132:{59,59}]
  wire  _GEN_318 = 9'h13a == _GEN_13709 ? meta_314_valid_0 : _GEN_317; // @[ICache.scala 132:{59,59}]
  wire  _GEN_319 = 9'h13b == _GEN_13709 ? meta_315_valid_0 : _GEN_318; // @[ICache.scala 132:{59,59}]
  wire  _GEN_320 = 9'h13c == _GEN_13709 ? meta_316_valid_0 : _GEN_319; // @[ICache.scala 132:{59,59}]
  wire  _GEN_321 = 9'h13d == _GEN_13709 ? meta_317_valid_0 : _GEN_320; // @[ICache.scala 132:{59,59}]
  wire  _GEN_322 = 9'h13e == _GEN_13709 ? meta_318_valid_0 : _GEN_321; // @[ICache.scala 132:{59,59}]
  wire  _GEN_323 = 9'h13f == _GEN_13709 ? meta_319_valid_0 : _GEN_322; // @[ICache.scala 132:{59,59}]
  wire  _GEN_324 = 9'h140 == _GEN_13709 ? meta_320_valid_0 : _GEN_323; // @[ICache.scala 132:{59,59}]
  wire  _GEN_325 = 9'h141 == _GEN_13709 ? meta_321_valid_0 : _GEN_324; // @[ICache.scala 132:{59,59}]
  wire  _GEN_326 = 9'h142 == _GEN_13709 ? meta_322_valid_0 : _GEN_325; // @[ICache.scala 132:{59,59}]
  wire  _GEN_327 = 9'h143 == _GEN_13709 ? meta_323_valid_0 : _GEN_326; // @[ICache.scala 132:{59,59}]
  wire  _GEN_328 = 9'h144 == _GEN_13709 ? meta_324_valid_0 : _GEN_327; // @[ICache.scala 132:{59,59}]
  wire  _GEN_329 = 9'h145 == _GEN_13709 ? meta_325_valid_0 : _GEN_328; // @[ICache.scala 132:{59,59}]
  wire  _GEN_330 = 9'h146 == _GEN_13709 ? meta_326_valid_0 : _GEN_329; // @[ICache.scala 132:{59,59}]
  wire  _GEN_331 = 9'h147 == _GEN_13709 ? meta_327_valid_0 : _GEN_330; // @[ICache.scala 132:{59,59}]
  wire  _GEN_332 = 9'h148 == _GEN_13709 ? meta_328_valid_0 : _GEN_331; // @[ICache.scala 132:{59,59}]
  wire  _GEN_333 = 9'h149 == _GEN_13709 ? meta_329_valid_0 : _GEN_332; // @[ICache.scala 132:{59,59}]
  wire  _GEN_334 = 9'h14a == _GEN_13709 ? meta_330_valid_0 : _GEN_333; // @[ICache.scala 132:{59,59}]
  wire  _GEN_335 = 9'h14b == _GEN_13709 ? meta_331_valid_0 : _GEN_334; // @[ICache.scala 132:{59,59}]
  wire  _GEN_336 = 9'h14c == _GEN_13709 ? meta_332_valid_0 : _GEN_335; // @[ICache.scala 132:{59,59}]
  wire  _GEN_337 = 9'h14d == _GEN_13709 ? meta_333_valid_0 : _GEN_336; // @[ICache.scala 132:{59,59}]
  wire  _GEN_338 = 9'h14e == _GEN_13709 ? meta_334_valid_0 : _GEN_337; // @[ICache.scala 132:{59,59}]
  wire  _GEN_339 = 9'h14f == _GEN_13709 ? meta_335_valid_0 : _GEN_338; // @[ICache.scala 132:{59,59}]
  wire  _GEN_340 = 9'h150 == _GEN_13709 ? meta_336_valid_0 : _GEN_339; // @[ICache.scala 132:{59,59}]
  wire  _GEN_341 = 9'h151 == _GEN_13709 ? meta_337_valid_0 : _GEN_340; // @[ICache.scala 132:{59,59}]
  wire  _GEN_342 = 9'h152 == _GEN_13709 ? meta_338_valid_0 : _GEN_341; // @[ICache.scala 132:{59,59}]
  wire  _GEN_343 = 9'h153 == _GEN_13709 ? meta_339_valid_0 : _GEN_342; // @[ICache.scala 132:{59,59}]
  wire  _GEN_344 = 9'h154 == _GEN_13709 ? meta_340_valid_0 : _GEN_343; // @[ICache.scala 132:{59,59}]
  wire  _GEN_345 = 9'h155 == _GEN_13709 ? meta_341_valid_0 : _GEN_344; // @[ICache.scala 132:{59,59}]
  wire  _GEN_346 = 9'h156 == _GEN_13709 ? meta_342_valid_0 : _GEN_345; // @[ICache.scala 132:{59,59}]
  wire  _GEN_347 = 9'h157 == _GEN_13709 ? meta_343_valid_0 : _GEN_346; // @[ICache.scala 132:{59,59}]
  wire  _GEN_348 = 9'h158 == _GEN_13709 ? meta_344_valid_0 : _GEN_347; // @[ICache.scala 132:{59,59}]
  wire  _GEN_349 = 9'h159 == _GEN_13709 ? meta_345_valid_0 : _GEN_348; // @[ICache.scala 132:{59,59}]
  wire  _GEN_350 = 9'h15a == _GEN_13709 ? meta_346_valid_0 : _GEN_349; // @[ICache.scala 132:{59,59}]
  wire  _GEN_351 = 9'h15b == _GEN_13709 ? meta_347_valid_0 : _GEN_350; // @[ICache.scala 132:{59,59}]
  wire  _GEN_352 = 9'h15c == _GEN_13709 ? meta_348_valid_0 : _GEN_351; // @[ICache.scala 132:{59,59}]
  wire  _GEN_353 = 9'h15d == _GEN_13709 ? meta_349_valid_0 : _GEN_352; // @[ICache.scala 132:{59,59}]
  wire  _GEN_354 = 9'h15e == _GEN_13709 ? meta_350_valid_0 : _GEN_353; // @[ICache.scala 132:{59,59}]
  wire  _GEN_355 = 9'h15f == _GEN_13709 ? meta_351_valid_0 : _GEN_354; // @[ICache.scala 132:{59,59}]
  wire  _GEN_356 = 9'h160 == _GEN_13709 ? meta_352_valid_0 : _GEN_355; // @[ICache.scala 132:{59,59}]
  wire  _GEN_357 = 9'h161 == _GEN_13709 ? meta_353_valid_0 : _GEN_356; // @[ICache.scala 132:{59,59}]
  wire  _GEN_358 = 9'h162 == _GEN_13709 ? meta_354_valid_0 : _GEN_357; // @[ICache.scala 132:{59,59}]
  wire  _GEN_359 = 9'h163 == _GEN_13709 ? meta_355_valid_0 : _GEN_358; // @[ICache.scala 132:{59,59}]
  wire  _GEN_360 = 9'h164 == _GEN_13709 ? meta_356_valid_0 : _GEN_359; // @[ICache.scala 132:{59,59}]
  wire  _GEN_361 = 9'h165 == _GEN_13709 ? meta_357_valid_0 : _GEN_360; // @[ICache.scala 132:{59,59}]
  wire  _GEN_362 = 9'h166 == _GEN_13709 ? meta_358_valid_0 : _GEN_361; // @[ICache.scala 132:{59,59}]
  wire  _GEN_363 = 9'h167 == _GEN_13709 ? meta_359_valid_0 : _GEN_362; // @[ICache.scala 132:{59,59}]
  wire  _GEN_364 = 9'h168 == _GEN_13709 ? meta_360_valid_0 : _GEN_363; // @[ICache.scala 132:{59,59}]
  wire  _GEN_365 = 9'h169 == _GEN_13709 ? meta_361_valid_0 : _GEN_364; // @[ICache.scala 132:{59,59}]
  wire  _GEN_366 = 9'h16a == _GEN_13709 ? meta_362_valid_0 : _GEN_365; // @[ICache.scala 132:{59,59}]
  wire  _GEN_367 = 9'h16b == _GEN_13709 ? meta_363_valid_0 : _GEN_366; // @[ICache.scala 132:{59,59}]
  wire  _GEN_368 = 9'h16c == _GEN_13709 ? meta_364_valid_0 : _GEN_367; // @[ICache.scala 132:{59,59}]
  wire  _GEN_369 = 9'h16d == _GEN_13709 ? meta_365_valid_0 : _GEN_368; // @[ICache.scala 132:{59,59}]
  wire  _GEN_370 = 9'h16e == _GEN_13709 ? meta_366_valid_0 : _GEN_369; // @[ICache.scala 132:{59,59}]
  wire  _GEN_371 = 9'h16f == _GEN_13709 ? meta_367_valid_0 : _GEN_370; // @[ICache.scala 132:{59,59}]
  wire  _GEN_372 = 9'h170 == _GEN_13709 ? meta_368_valid_0 : _GEN_371; // @[ICache.scala 132:{59,59}]
  wire  _GEN_373 = 9'h171 == _GEN_13709 ? meta_369_valid_0 : _GEN_372; // @[ICache.scala 132:{59,59}]
  wire  _GEN_374 = 9'h172 == _GEN_13709 ? meta_370_valid_0 : _GEN_373; // @[ICache.scala 132:{59,59}]
  wire  _GEN_375 = 9'h173 == _GEN_13709 ? meta_371_valid_0 : _GEN_374; // @[ICache.scala 132:{59,59}]
  wire  _GEN_376 = 9'h174 == _GEN_13709 ? meta_372_valid_0 : _GEN_375; // @[ICache.scala 132:{59,59}]
  wire  _GEN_377 = 9'h175 == _GEN_13709 ? meta_373_valid_0 : _GEN_376; // @[ICache.scala 132:{59,59}]
  wire  _GEN_378 = 9'h176 == _GEN_13709 ? meta_374_valid_0 : _GEN_377; // @[ICache.scala 132:{59,59}]
  wire  _GEN_379 = 9'h177 == _GEN_13709 ? meta_375_valid_0 : _GEN_378; // @[ICache.scala 132:{59,59}]
  wire  _GEN_380 = 9'h178 == _GEN_13709 ? meta_376_valid_0 : _GEN_379; // @[ICache.scala 132:{59,59}]
  wire  _GEN_381 = 9'h179 == _GEN_13709 ? meta_377_valid_0 : _GEN_380; // @[ICache.scala 132:{59,59}]
  wire  _GEN_382 = 9'h17a == _GEN_13709 ? meta_378_valid_0 : _GEN_381; // @[ICache.scala 132:{59,59}]
  wire  _GEN_383 = 9'h17b == _GEN_13709 ? meta_379_valid_0 : _GEN_382; // @[ICache.scala 132:{59,59}]
  wire  _GEN_384 = 9'h17c == _GEN_13709 ? meta_380_valid_0 : _GEN_383; // @[ICache.scala 132:{59,59}]
  wire  _GEN_385 = 9'h17d == _GEN_13709 ? meta_381_valid_0 : _GEN_384; // @[ICache.scala 132:{59,59}]
  wire  _GEN_386 = 9'h17e == _GEN_13709 ? meta_382_valid_0 : _GEN_385; // @[ICache.scala 132:{59,59}]
  wire  _GEN_387 = 9'h17f == _GEN_13709 ? meta_383_valid_0 : _GEN_386; // @[ICache.scala 132:{59,59}]
  wire  _GEN_388 = 9'h180 == _GEN_13709 ? meta_384_valid_0 : _GEN_387; // @[ICache.scala 132:{59,59}]
  wire  _GEN_389 = 9'h181 == _GEN_13709 ? meta_385_valid_0 : _GEN_388; // @[ICache.scala 132:{59,59}]
  wire  _GEN_390 = 9'h182 == _GEN_13709 ? meta_386_valid_0 : _GEN_389; // @[ICache.scala 132:{59,59}]
  wire  _GEN_391 = 9'h183 == _GEN_13709 ? meta_387_valid_0 : _GEN_390; // @[ICache.scala 132:{59,59}]
  wire  _GEN_392 = 9'h184 == _GEN_13709 ? meta_388_valid_0 : _GEN_391; // @[ICache.scala 132:{59,59}]
  wire  _GEN_393 = 9'h185 == _GEN_13709 ? meta_389_valid_0 : _GEN_392; // @[ICache.scala 132:{59,59}]
  wire  _GEN_394 = 9'h186 == _GEN_13709 ? meta_390_valid_0 : _GEN_393; // @[ICache.scala 132:{59,59}]
  wire  _GEN_395 = 9'h187 == _GEN_13709 ? meta_391_valid_0 : _GEN_394; // @[ICache.scala 132:{59,59}]
  wire  _GEN_396 = 9'h188 == _GEN_13709 ? meta_392_valid_0 : _GEN_395; // @[ICache.scala 132:{59,59}]
  wire  _GEN_397 = 9'h189 == _GEN_13709 ? meta_393_valid_0 : _GEN_396; // @[ICache.scala 132:{59,59}]
  wire  _GEN_398 = 9'h18a == _GEN_13709 ? meta_394_valid_0 : _GEN_397; // @[ICache.scala 132:{59,59}]
  wire  _GEN_399 = 9'h18b == _GEN_13709 ? meta_395_valid_0 : _GEN_398; // @[ICache.scala 132:{59,59}]
  wire  _GEN_400 = 9'h18c == _GEN_13709 ? meta_396_valid_0 : _GEN_399; // @[ICache.scala 132:{59,59}]
  wire  _GEN_401 = 9'h18d == _GEN_13709 ? meta_397_valid_0 : _GEN_400; // @[ICache.scala 132:{59,59}]
  wire  _GEN_402 = 9'h18e == _GEN_13709 ? meta_398_valid_0 : _GEN_401; // @[ICache.scala 132:{59,59}]
  wire  _GEN_403 = 9'h18f == _GEN_13709 ? meta_399_valid_0 : _GEN_402; // @[ICache.scala 132:{59,59}]
  wire  _GEN_404 = 9'h190 == _GEN_13709 ? meta_400_valid_0 : _GEN_403; // @[ICache.scala 132:{59,59}]
  wire  _GEN_405 = 9'h191 == _GEN_13709 ? meta_401_valid_0 : _GEN_404; // @[ICache.scala 132:{59,59}]
  wire  _GEN_406 = 9'h192 == _GEN_13709 ? meta_402_valid_0 : _GEN_405; // @[ICache.scala 132:{59,59}]
  wire  _GEN_407 = 9'h193 == _GEN_13709 ? meta_403_valid_0 : _GEN_406; // @[ICache.scala 132:{59,59}]
  wire  _GEN_408 = 9'h194 == _GEN_13709 ? meta_404_valid_0 : _GEN_407; // @[ICache.scala 132:{59,59}]
  wire  _GEN_409 = 9'h195 == _GEN_13709 ? meta_405_valid_0 : _GEN_408; // @[ICache.scala 132:{59,59}]
  wire  _GEN_410 = 9'h196 == _GEN_13709 ? meta_406_valid_0 : _GEN_409; // @[ICache.scala 132:{59,59}]
  wire  _GEN_411 = 9'h197 == _GEN_13709 ? meta_407_valid_0 : _GEN_410; // @[ICache.scala 132:{59,59}]
  wire  _GEN_412 = 9'h198 == _GEN_13709 ? meta_408_valid_0 : _GEN_411; // @[ICache.scala 132:{59,59}]
  wire  _GEN_413 = 9'h199 == _GEN_13709 ? meta_409_valid_0 : _GEN_412; // @[ICache.scala 132:{59,59}]
  wire  _GEN_414 = 9'h19a == _GEN_13709 ? meta_410_valid_0 : _GEN_413; // @[ICache.scala 132:{59,59}]
  wire  _GEN_415 = 9'h19b == _GEN_13709 ? meta_411_valid_0 : _GEN_414; // @[ICache.scala 132:{59,59}]
  wire  _GEN_416 = 9'h19c == _GEN_13709 ? meta_412_valid_0 : _GEN_415; // @[ICache.scala 132:{59,59}]
  wire  _GEN_417 = 9'h19d == _GEN_13709 ? meta_413_valid_0 : _GEN_416; // @[ICache.scala 132:{59,59}]
  wire  _GEN_418 = 9'h19e == _GEN_13709 ? meta_414_valid_0 : _GEN_417; // @[ICache.scala 132:{59,59}]
  wire  _GEN_419 = 9'h19f == _GEN_13709 ? meta_415_valid_0 : _GEN_418; // @[ICache.scala 132:{59,59}]
  wire  _GEN_420 = 9'h1a0 == _GEN_13709 ? meta_416_valid_0 : _GEN_419; // @[ICache.scala 132:{59,59}]
  wire  _GEN_421 = 9'h1a1 == _GEN_13709 ? meta_417_valid_0 : _GEN_420; // @[ICache.scala 132:{59,59}]
  wire  _GEN_422 = 9'h1a2 == _GEN_13709 ? meta_418_valid_0 : _GEN_421; // @[ICache.scala 132:{59,59}]
  wire  _GEN_423 = 9'h1a3 == _GEN_13709 ? meta_419_valid_0 : _GEN_422; // @[ICache.scala 132:{59,59}]
  wire  _GEN_424 = 9'h1a4 == _GEN_13709 ? meta_420_valid_0 : _GEN_423; // @[ICache.scala 132:{59,59}]
  wire  _GEN_425 = 9'h1a5 == _GEN_13709 ? meta_421_valid_0 : _GEN_424; // @[ICache.scala 132:{59,59}]
  wire  _GEN_426 = 9'h1a6 == _GEN_13709 ? meta_422_valid_0 : _GEN_425; // @[ICache.scala 132:{59,59}]
  wire  _GEN_427 = 9'h1a7 == _GEN_13709 ? meta_423_valid_0 : _GEN_426; // @[ICache.scala 132:{59,59}]
  wire  _GEN_428 = 9'h1a8 == _GEN_13709 ? meta_424_valid_0 : _GEN_427; // @[ICache.scala 132:{59,59}]
  wire  _GEN_429 = 9'h1a9 == _GEN_13709 ? meta_425_valid_0 : _GEN_428; // @[ICache.scala 132:{59,59}]
  wire  _GEN_430 = 9'h1aa == _GEN_13709 ? meta_426_valid_0 : _GEN_429; // @[ICache.scala 132:{59,59}]
  wire  _GEN_431 = 9'h1ab == _GEN_13709 ? meta_427_valid_0 : _GEN_430; // @[ICache.scala 132:{59,59}]
  wire  _GEN_432 = 9'h1ac == _GEN_13709 ? meta_428_valid_0 : _GEN_431; // @[ICache.scala 132:{59,59}]
  wire  _GEN_433 = 9'h1ad == _GEN_13709 ? meta_429_valid_0 : _GEN_432; // @[ICache.scala 132:{59,59}]
  wire  _GEN_434 = 9'h1ae == _GEN_13709 ? meta_430_valid_0 : _GEN_433; // @[ICache.scala 132:{59,59}]
  wire  _GEN_435 = 9'h1af == _GEN_13709 ? meta_431_valid_0 : _GEN_434; // @[ICache.scala 132:{59,59}]
  wire  _GEN_436 = 9'h1b0 == _GEN_13709 ? meta_432_valid_0 : _GEN_435; // @[ICache.scala 132:{59,59}]
  wire  _GEN_437 = 9'h1b1 == _GEN_13709 ? meta_433_valid_0 : _GEN_436; // @[ICache.scala 132:{59,59}]
  wire  _GEN_438 = 9'h1b2 == _GEN_13709 ? meta_434_valid_0 : _GEN_437; // @[ICache.scala 132:{59,59}]
  wire  _GEN_439 = 9'h1b3 == _GEN_13709 ? meta_435_valid_0 : _GEN_438; // @[ICache.scala 132:{59,59}]
  wire  _GEN_440 = 9'h1b4 == _GEN_13709 ? meta_436_valid_0 : _GEN_439; // @[ICache.scala 132:{59,59}]
  wire  _GEN_441 = 9'h1b5 == _GEN_13709 ? meta_437_valid_0 : _GEN_440; // @[ICache.scala 132:{59,59}]
  wire  _GEN_442 = 9'h1b6 == _GEN_13709 ? meta_438_valid_0 : _GEN_441; // @[ICache.scala 132:{59,59}]
  wire  _GEN_443 = 9'h1b7 == _GEN_13709 ? meta_439_valid_0 : _GEN_442; // @[ICache.scala 132:{59,59}]
  wire  _GEN_444 = 9'h1b8 == _GEN_13709 ? meta_440_valid_0 : _GEN_443; // @[ICache.scala 132:{59,59}]
  wire  _GEN_445 = 9'h1b9 == _GEN_13709 ? meta_441_valid_0 : _GEN_444; // @[ICache.scala 132:{59,59}]
  wire  _GEN_446 = 9'h1ba == _GEN_13709 ? meta_442_valid_0 : _GEN_445; // @[ICache.scala 132:{59,59}]
  wire  _GEN_447 = 9'h1bb == _GEN_13709 ? meta_443_valid_0 : _GEN_446; // @[ICache.scala 132:{59,59}]
  wire  _GEN_448 = 9'h1bc == _GEN_13709 ? meta_444_valid_0 : _GEN_447; // @[ICache.scala 132:{59,59}]
  wire  _GEN_449 = 9'h1bd == _GEN_13709 ? meta_445_valid_0 : _GEN_448; // @[ICache.scala 132:{59,59}]
  wire  _GEN_450 = 9'h1be == _GEN_13709 ? meta_446_valid_0 : _GEN_449; // @[ICache.scala 132:{59,59}]
  wire  _GEN_451 = 9'h1bf == _GEN_13709 ? meta_447_valid_0 : _GEN_450; // @[ICache.scala 132:{59,59}]
  wire  _GEN_452 = 9'h1c0 == _GEN_13709 ? meta_448_valid_0 : _GEN_451; // @[ICache.scala 132:{59,59}]
  wire  _GEN_453 = 9'h1c1 == _GEN_13709 ? meta_449_valid_0 : _GEN_452; // @[ICache.scala 132:{59,59}]
  wire  _GEN_454 = 9'h1c2 == _GEN_13709 ? meta_450_valid_0 : _GEN_453; // @[ICache.scala 132:{59,59}]
  wire  _GEN_455 = 9'h1c3 == _GEN_13709 ? meta_451_valid_0 : _GEN_454; // @[ICache.scala 132:{59,59}]
  wire  _GEN_456 = 9'h1c4 == _GEN_13709 ? meta_452_valid_0 : _GEN_455; // @[ICache.scala 132:{59,59}]
  wire  _GEN_457 = 9'h1c5 == _GEN_13709 ? meta_453_valid_0 : _GEN_456; // @[ICache.scala 132:{59,59}]
  wire  _GEN_458 = 9'h1c6 == _GEN_13709 ? meta_454_valid_0 : _GEN_457; // @[ICache.scala 132:{59,59}]
  wire  _GEN_459 = 9'h1c7 == _GEN_13709 ? meta_455_valid_0 : _GEN_458; // @[ICache.scala 132:{59,59}]
  wire  _GEN_460 = 9'h1c8 == _GEN_13709 ? meta_456_valid_0 : _GEN_459; // @[ICache.scala 132:{59,59}]
  wire  _GEN_461 = 9'h1c9 == _GEN_13709 ? meta_457_valid_0 : _GEN_460; // @[ICache.scala 132:{59,59}]
  wire  _GEN_462 = 9'h1ca == _GEN_13709 ? meta_458_valid_0 : _GEN_461; // @[ICache.scala 132:{59,59}]
  wire  _GEN_463 = 9'h1cb == _GEN_13709 ? meta_459_valid_0 : _GEN_462; // @[ICache.scala 132:{59,59}]
  wire  _GEN_464 = 9'h1cc == _GEN_13709 ? meta_460_valid_0 : _GEN_463; // @[ICache.scala 132:{59,59}]
  wire  _GEN_465 = 9'h1cd == _GEN_13709 ? meta_461_valid_0 : _GEN_464; // @[ICache.scala 132:{59,59}]
  wire  _GEN_466 = 9'h1ce == _GEN_13709 ? meta_462_valid_0 : _GEN_465; // @[ICache.scala 132:{59,59}]
  wire  _GEN_467 = 9'h1cf == _GEN_13709 ? meta_463_valid_0 : _GEN_466; // @[ICache.scala 132:{59,59}]
  wire  _GEN_468 = 9'h1d0 == _GEN_13709 ? meta_464_valid_0 : _GEN_467; // @[ICache.scala 132:{59,59}]
  wire  _GEN_469 = 9'h1d1 == _GEN_13709 ? meta_465_valid_0 : _GEN_468; // @[ICache.scala 132:{59,59}]
  wire  _GEN_470 = 9'h1d2 == _GEN_13709 ? meta_466_valid_0 : _GEN_469; // @[ICache.scala 132:{59,59}]
  wire  _GEN_471 = 9'h1d3 == _GEN_13709 ? meta_467_valid_0 : _GEN_470; // @[ICache.scala 132:{59,59}]
  wire  _GEN_472 = 9'h1d4 == _GEN_13709 ? meta_468_valid_0 : _GEN_471; // @[ICache.scala 132:{59,59}]
  wire  _GEN_473 = 9'h1d5 == _GEN_13709 ? meta_469_valid_0 : _GEN_472; // @[ICache.scala 132:{59,59}]
  wire  _GEN_474 = 9'h1d6 == _GEN_13709 ? meta_470_valid_0 : _GEN_473; // @[ICache.scala 132:{59,59}]
  wire  _GEN_475 = 9'h1d7 == _GEN_13709 ? meta_471_valid_0 : _GEN_474; // @[ICache.scala 132:{59,59}]
  wire  _GEN_476 = 9'h1d8 == _GEN_13709 ? meta_472_valid_0 : _GEN_475; // @[ICache.scala 132:{59,59}]
  wire  _GEN_477 = 9'h1d9 == _GEN_13709 ? meta_473_valid_0 : _GEN_476; // @[ICache.scala 132:{59,59}]
  wire  _GEN_478 = 9'h1da == _GEN_13709 ? meta_474_valid_0 : _GEN_477; // @[ICache.scala 132:{59,59}]
  wire  _GEN_479 = 9'h1db == _GEN_13709 ? meta_475_valid_0 : _GEN_478; // @[ICache.scala 132:{59,59}]
  wire  _GEN_480 = 9'h1dc == _GEN_13709 ? meta_476_valid_0 : _GEN_479; // @[ICache.scala 132:{59,59}]
  wire  _GEN_481 = 9'h1dd == _GEN_13709 ? meta_477_valid_0 : _GEN_480; // @[ICache.scala 132:{59,59}]
  wire  _GEN_482 = 9'h1de == _GEN_13709 ? meta_478_valid_0 : _GEN_481; // @[ICache.scala 132:{59,59}]
  wire  _GEN_483 = 9'h1df == _GEN_13709 ? meta_479_valid_0 : _GEN_482; // @[ICache.scala 132:{59,59}]
  wire  _GEN_484 = 9'h1e0 == _GEN_13709 ? meta_480_valid_0 : _GEN_483; // @[ICache.scala 132:{59,59}]
  wire  _GEN_485 = 9'h1e1 == _GEN_13709 ? meta_481_valid_0 : _GEN_484; // @[ICache.scala 132:{59,59}]
  wire  _GEN_486 = 9'h1e2 == _GEN_13709 ? meta_482_valid_0 : _GEN_485; // @[ICache.scala 132:{59,59}]
  wire  _GEN_487 = 9'h1e3 == _GEN_13709 ? meta_483_valid_0 : _GEN_486; // @[ICache.scala 132:{59,59}]
  wire  _GEN_488 = 9'h1e4 == _GEN_13709 ? meta_484_valid_0 : _GEN_487; // @[ICache.scala 132:{59,59}]
  wire  _GEN_489 = 9'h1e5 == _GEN_13709 ? meta_485_valid_0 : _GEN_488; // @[ICache.scala 132:{59,59}]
  wire  _GEN_490 = 9'h1e6 == _GEN_13709 ? meta_486_valid_0 : _GEN_489; // @[ICache.scala 132:{59,59}]
  wire  _GEN_491 = 9'h1e7 == _GEN_13709 ? meta_487_valid_0 : _GEN_490; // @[ICache.scala 132:{59,59}]
  wire  _GEN_492 = 9'h1e8 == _GEN_13709 ? meta_488_valid_0 : _GEN_491; // @[ICache.scala 132:{59,59}]
  wire  _GEN_493 = 9'h1e9 == _GEN_13709 ? meta_489_valid_0 : _GEN_492; // @[ICache.scala 132:{59,59}]
  wire  _GEN_494 = 9'h1ea == _GEN_13709 ? meta_490_valid_0 : _GEN_493; // @[ICache.scala 132:{59,59}]
  wire  _GEN_495 = 9'h1eb == _GEN_13709 ? meta_491_valid_0 : _GEN_494; // @[ICache.scala 132:{59,59}]
  wire  _GEN_496 = 9'h1ec == _GEN_13709 ? meta_492_valid_0 : _GEN_495; // @[ICache.scala 132:{59,59}]
  wire  _GEN_497 = 9'h1ed == _GEN_13709 ? meta_493_valid_0 : _GEN_496; // @[ICache.scala 132:{59,59}]
  wire  _GEN_498 = 9'h1ee == _GEN_13709 ? meta_494_valid_0 : _GEN_497; // @[ICache.scala 132:{59,59}]
  wire  _GEN_499 = 9'h1ef == _GEN_13709 ? meta_495_valid_0 : _GEN_498; // @[ICache.scala 132:{59,59}]
  wire  _GEN_500 = 9'h1f0 == _GEN_13709 ? meta_496_valid_0 : _GEN_499; // @[ICache.scala 132:{59,59}]
  wire  _GEN_501 = 9'h1f1 == _GEN_13709 ? meta_497_valid_0 : _GEN_500; // @[ICache.scala 132:{59,59}]
  wire  _GEN_502 = 9'h1f2 == _GEN_13709 ? meta_498_valid_0 : _GEN_501; // @[ICache.scala 132:{59,59}]
  wire  _GEN_503 = 9'h1f3 == _GEN_13709 ? meta_499_valid_0 : _GEN_502; // @[ICache.scala 132:{59,59}]
  wire  _GEN_504 = 9'h1f4 == _GEN_13709 ? meta_500_valid_0 : _GEN_503; // @[ICache.scala 132:{59,59}]
  wire  _GEN_505 = 9'h1f5 == _GEN_13709 ? meta_501_valid_0 : _GEN_504; // @[ICache.scala 132:{59,59}]
  wire  _GEN_506 = 9'h1f6 == _GEN_13709 ? meta_502_valid_0 : _GEN_505; // @[ICache.scala 132:{59,59}]
  wire  _GEN_507 = 9'h1f7 == _GEN_13709 ? meta_503_valid_0 : _GEN_506; // @[ICache.scala 132:{59,59}]
  wire  _GEN_508 = 9'h1f8 == _GEN_13709 ? meta_504_valid_0 : _GEN_507; // @[ICache.scala 132:{59,59}]
  wire  _GEN_509 = 9'h1f9 == _GEN_13709 ? meta_505_valid_0 : _GEN_508; // @[ICache.scala 132:{59,59}]
  wire  _GEN_510 = 9'h1fa == _GEN_13709 ? meta_506_valid_0 : _GEN_509; // @[ICache.scala 132:{59,59}]
  wire  _GEN_511 = 9'h1fb == _GEN_13709 ? meta_507_valid_0 : _GEN_510; // @[ICache.scala 132:{59,59}]
  wire  _GEN_512 = 9'h1fc == _GEN_13709 ? meta_508_valid_0 : _GEN_511; // @[ICache.scala 132:{59,59}]
  wire  _GEN_513 = 9'h1fd == _GEN_13709 ? meta_509_valid_0 : _GEN_512; // @[ICache.scala 132:{59,59}]
  wire  _GEN_514 = 9'h1fe == _GEN_13709 ? meta_510_valid_0 : _GEN_513; // @[ICache.scala 132:{59,59}]
  wire  _GEN_515 = 9'h1ff == _GEN_13709 ? meta_511_valid_0 : _GEN_514; // @[ICache.scala 132:{59,59}]
  wire  tag_compare_valid_0 = _GEN_13516 == inst_tag & _GEN_515; // @[ICache.scala 132:59]
  wire [16:0] cache_tag_1 = tag_ram_io_way_1_r_data; // @[ICache.scala 64:28 131:30]
  wire [19:0] _GEN_13965 = {{3'd0}, cache_tag_1}; // @[ICache.scala 132:46]
  wire  _GEN_517 = 6'h1 == va_line_addr ? meta_1_valid_1 : meta_0_valid_1; // @[ICache.scala 132:{59,59}]
  wire  _GEN_518 = 6'h2 == va_line_addr ? meta_2_valid_1 : _GEN_517; // @[ICache.scala 132:{59,59}]
  wire  _GEN_519 = 6'h3 == va_line_addr ? meta_3_valid_1 : _GEN_518; // @[ICache.scala 132:{59,59}]
  wire  _GEN_520 = 6'h4 == va_line_addr ? meta_4_valid_1 : _GEN_519; // @[ICache.scala 132:{59,59}]
  wire  _GEN_521 = 6'h5 == va_line_addr ? meta_5_valid_1 : _GEN_520; // @[ICache.scala 132:{59,59}]
  wire  _GEN_522 = 6'h6 == va_line_addr ? meta_6_valid_1 : _GEN_521; // @[ICache.scala 132:{59,59}]
  wire  _GEN_523 = 6'h7 == va_line_addr ? meta_7_valid_1 : _GEN_522; // @[ICache.scala 132:{59,59}]
  wire  _GEN_524 = 6'h8 == va_line_addr ? meta_8_valid_1 : _GEN_523; // @[ICache.scala 132:{59,59}]
  wire  _GEN_525 = 6'h9 == va_line_addr ? meta_9_valid_1 : _GEN_524; // @[ICache.scala 132:{59,59}]
  wire  _GEN_526 = 6'ha == va_line_addr ? meta_10_valid_1 : _GEN_525; // @[ICache.scala 132:{59,59}]
  wire  _GEN_527 = 6'hb == va_line_addr ? meta_11_valid_1 : _GEN_526; // @[ICache.scala 132:{59,59}]
  wire  _GEN_528 = 6'hc == va_line_addr ? meta_12_valid_1 : _GEN_527; // @[ICache.scala 132:{59,59}]
  wire  _GEN_529 = 6'hd == va_line_addr ? meta_13_valid_1 : _GEN_528; // @[ICache.scala 132:{59,59}]
  wire  _GEN_530 = 6'he == va_line_addr ? meta_14_valid_1 : _GEN_529; // @[ICache.scala 132:{59,59}]
  wire  _GEN_531 = 6'hf == va_line_addr ? meta_15_valid_1 : _GEN_530; // @[ICache.scala 132:{59,59}]
  wire  _GEN_532 = 6'h10 == va_line_addr ? meta_16_valid_1 : _GEN_531; // @[ICache.scala 132:{59,59}]
  wire  _GEN_533 = 6'h11 == va_line_addr ? meta_17_valid_1 : _GEN_532; // @[ICache.scala 132:{59,59}]
  wire  _GEN_534 = 6'h12 == va_line_addr ? meta_18_valid_1 : _GEN_533; // @[ICache.scala 132:{59,59}]
  wire  _GEN_535 = 6'h13 == va_line_addr ? meta_19_valid_1 : _GEN_534; // @[ICache.scala 132:{59,59}]
  wire  _GEN_536 = 6'h14 == va_line_addr ? meta_20_valid_1 : _GEN_535; // @[ICache.scala 132:{59,59}]
  wire  _GEN_537 = 6'h15 == va_line_addr ? meta_21_valid_1 : _GEN_536; // @[ICache.scala 132:{59,59}]
  wire  _GEN_538 = 6'h16 == va_line_addr ? meta_22_valid_1 : _GEN_537; // @[ICache.scala 132:{59,59}]
  wire  _GEN_539 = 6'h17 == va_line_addr ? meta_23_valid_1 : _GEN_538; // @[ICache.scala 132:{59,59}]
  wire  _GEN_540 = 6'h18 == va_line_addr ? meta_24_valid_1 : _GEN_539; // @[ICache.scala 132:{59,59}]
  wire  _GEN_541 = 6'h19 == va_line_addr ? meta_25_valid_1 : _GEN_540; // @[ICache.scala 132:{59,59}]
  wire  _GEN_542 = 6'h1a == va_line_addr ? meta_26_valid_1 : _GEN_541; // @[ICache.scala 132:{59,59}]
  wire  _GEN_543 = 6'h1b == va_line_addr ? meta_27_valid_1 : _GEN_542; // @[ICache.scala 132:{59,59}]
  wire  _GEN_544 = 6'h1c == va_line_addr ? meta_28_valid_1 : _GEN_543; // @[ICache.scala 132:{59,59}]
  wire  _GEN_545 = 6'h1d == va_line_addr ? meta_29_valid_1 : _GEN_544; // @[ICache.scala 132:{59,59}]
  wire  _GEN_546 = 6'h1e == va_line_addr ? meta_30_valid_1 : _GEN_545; // @[ICache.scala 132:{59,59}]
  wire  _GEN_547 = 6'h1f == va_line_addr ? meta_31_valid_1 : _GEN_546; // @[ICache.scala 132:{59,59}]
  wire  _GEN_548 = 6'h20 == va_line_addr ? meta_32_valid_1 : _GEN_547; // @[ICache.scala 132:{59,59}]
  wire  _GEN_549 = 6'h21 == va_line_addr ? meta_33_valid_1 : _GEN_548; // @[ICache.scala 132:{59,59}]
  wire  _GEN_550 = 6'h22 == va_line_addr ? meta_34_valid_1 : _GEN_549; // @[ICache.scala 132:{59,59}]
  wire  _GEN_551 = 6'h23 == va_line_addr ? meta_35_valid_1 : _GEN_550; // @[ICache.scala 132:{59,59}]
  wire  _GEN_552 = 6'h24 == va_line_addr ? meta_36_valid_1 : _GEN_551; // @[ICache.scala 132:{59,59}]
  wire  _GEN_553 = 6'h25 == va_line_addr ? meta_37_valid_1 : _GEN_552; // @[ICache.scala 132:{59,59}]
  wire  _GEN_554 = 6'h26 == va_line_addr ? meta_38_valid_1 : _GEN_553; // @[ICache.scala 132:{59,59}]
  wire  _GEN_555 = 6'h27 == va_line_addr ? meta_39_valid_1 : _GEN_554; // @[ICache.scala 132:{59,59}]
  wire  _GEN_556 = 6'h28 == va_line_addr ? meta_40_valid_1 : _GEN_555; // @[ICache.scala 132:{59,59}]
  wire  _GEN_557 = 6'h29 == va_line_addr ? meta_41_valid_1 : _GEN_556; // @[ICache.scala 132:{59,59}]
  wire  _GEN_558 = 6'h2a == va_line_addr ? meta_42_valid_1 : _GEN_557; // @[ICache.scala 132:{59,59}]
  wire  _GEN_559 = 6'h2b == va_line_addr ? meta_43_valid_1 : _GEN_558; // @[ICache.scala 132:{59,59}]
  wire  _GEN_560 = 6'h2c == va_line_addr ? meta_44_valid_1 : _GEN_559; // @[ICache.scala 132:{59,59}]
  wire  _GEN_561 = 6'h2d == va_line_addr ? meta_45_valid_1 : _GEN_560; // @[ICache.scala 132:{59,59}]
  wire  _GEN_562 = 6'h2e == va_line_addr ? meta_46_valid_1 : _GEN_561; // @[ICache.scala 132:{59,59}]
  wire  _GEN_563 = 6'h2f == va_line_addr ? meta_47_valid_1 : _GEN_562; // @[ICache.scala 132:{59,59}]
  wire  _GEN_564 = 6'h30 == va_line_addr ? meta_48_valid_1 : _GEN_563; // @[ICache.scala 132:{59,59}]
  wire  _GEN_565 = 6'h31 == va_line_addr ? meta_49_valid_1 : _GEN_564; // @[ICache.scala 132:{59,59}]
  wire  _GEN_566 = 6'h32 == va_line_addr ? meta_50_valid_1 : _GEN_565; // @[ICache.scala 132:{59,59}]
  wire  _GEN_567 = 6'h33 == va_line_addr ? meta_51_valid_1 : _GEN_566; // @[ICache.scala 132:{59,59}]
  wire  _GEN_568 = 6'h34 == va_line_addr ? meta_52_valid_1 : _GEN_567; // @[ICache.scala 132:{59,59}]
  wire  _GEN_569 = 6'h35 == va_line_addr ? meta_53_valid_1 : _GEN_568; // @[ICache.scala 132:{59,59}]
  wire  _GEN_570 = 6'h36 == va_line_addr ? meta_54_valid_1 : _GEN_569; // @[ICache.scala 132:{59,59}]
  wire  _GEN_571 = 6'h37 == va_line_addr ? meta_55_valid_1 : _GEN_570; // @[ICache.scala 132:{59,59}]
  wire  _GEN_572 = 6'h38 == va_line_addr ? meta_56_valid_1 : _GEN_571; // @[ICache.scala 132:{59,59}]
  wire  _GEN_573 = 6'h39 == va_line_addr ? meta_57_valid_1 : _GEN_572; // @[ICache.scala 132:{59,59}]
  wire  _GEN_574 = 6'h3a == va_line_addr ? meta_58_valid_1 : _GEN_573; // @[ICache.scala 132:{59,59}]
  wire  _GEN_575 = 6'h3b == va_line_addr ? meta_59_valid_1 : _GEN_574; // @[ICache.scala 132:{59,59}]
  wire  _GEN_576 = 6'h3c == va_line_addr ? meta_60_valid_1 : _GEN_575; // @[ICache.scala 132:{59,59}]
  wire  _GEN_577 = 6'h3d == va_line_addr ? meta_61_valid_1 : _GEN_576; // @[ICache.scala 132:{59,59}]
  wire  _GEN_578 = 6'h3e == va_line_addr ? meta_62_valid_1 : _GEN_577; // @[ICache.scala 132:{59,59}]
  wire  _GEN_579 = 6'h3f == va_line_addr ? meta_63_valid_1 : _GEN_578; // @[ICache.scala 132:{59,59}]
  wire  _GEN_580 = 7'h40 == _GEN_13517 ? meta_64_valid_1 : _GEN_579; // @[ICache.scala 132:{59,59}]
  wire  _GEN_581 = 7'h41 == _GEN_13517 ? meta_65_valid_1 : _GEN_580; // @[ICache.scala 132:{59,59}]
  wire  _GEN_582 = 7'h42 == _GEN_13517 ? meta_66_valid_1 : _GEN_581; // @[ICache.scala 132:{59,59}]
  wire  _GEN_583 = 7'h43 == _GEN_13517 ? meta_67_valid_1 : _GEN_582; // @[ICache.scala 132:{59,59}]
  wire  _GEN_584 = 7'h44 == _GEN_13517 ? meta_68_valid_1 : _GEN_583; // @[ICache.scala 132:{59,59}]
  wire  _GEN_585 = 7'h45 == _GEN_13517 ? meta_69_valid_1 : _GEN_584; // @[ICache.scala 132:{59,59}]
  wire  _GEN_586 = 7'h46 == _GEN_13517 ? meta_70_valid_1 : _GEN_585; // @[ICache.scala 132:{59,59}]
  wire  _GEN_587 = 7'h47 == _GEN_13517 ? meta_71_valid_1 : _GEN_586; // @[ICache.scala 132:{59,59}]
  wire  _GEN_588 = 7'h48 == _GEN_13517 ? meta_72_valid_1 : _GEN_587; // @[ICache.scala 132:{59,59}]
  wire  _GEN_589 = 7'h49 == _GEN_13517 ? meta_73_valid_1 : _GEN_588; // @[ICache.scala 132:{59,59}]
  wire  _GEN_590 = 7'h4a == _GEN_13517 ? meta_74_valid_1 : _GEN_589; // @[ICache.scala 132:{59,59}]
  wire  _GEN_591 = 7'h4b == _GEN_13517 ? meta_75_valid_1 : _GEN_590; // @[ICache.scala 132:{59,59}]
  wire  _GEN_592 = 7'h4c == _GEN_13517 ? meta_76_valid_1 : _GEN_591; // @[ICache.scala 132:{59,59}]
  wire  _GEN_593 = 7'h4d == _GEN_13517 ? meta_77_valid_1 : _GEN_592; // @[ICache.scala 132:{59,59}]
  wire  _GEN_594 = 7'h4e == _GEN_13517 ? meta_78_valid_1 : _GEN_593; // @[ICache.scala 132:{59,59}]
  wire  _GEN_595 = 7'h4f == _GEN_13517 ? meta_79_valid_1 : _GEN_594; // @[ICache.scala 132:{59,59}]
  wire  _GEN_596 = 7'h50 == _GEN_13517 ? meta_80_valid_1 : _GEN_595; // @[ICache.scala 132:{59,59}]
  wire  _GEN_597 = 7'h51 == _GEN_13517 ? meta_81_valid_1 : _GEN_596; // @[ICache.scala 132:{59,59}]
  wire  _GEN_598 = 7'h52 == _GEN_13517 ? meta_82_valid_1 : _GEN_597; // @[ICache.scala 132:{59,59}]
  wire  _GEN_599 = 7'h53 == _GEN_13517 ? meta_83_valid_1 : _GEN_598; // @[ICache.scala 132:{59,59}]
  wire  _GEN_600 = 7'h54 == _GEN_13517 ? meta_84_valid_1 : _GEN_599; // @[ICache.scala 132:{59,59}]
  wire  _GEN_601 = 7'h55 == _GEN_13517 ? meta_85_valid_1 : _GEN_600; // @[ICache.scala 132:{59,59}]
  wire  _GEN_602 = 7'h56 == _GEN_13517 ? meta_86_valid_1 : _GEN_601; // @[ICache.scala 132:{59,59}]
  wire  _GEN_603 = 7'h57 == _GEN_13517 ? meta_87_valid_1 : _GEN_602; // @[ICache.scala 132:{59,59}]
  wire  _GEN_604 = 7'h58 == _GEN_13517 ? meta_88_valid_1 : _GEN_603; // @[ICache.scala 132:{59,59}]
  wire  _GEN_605 = 7'h59 == _GEN_13517 ? meta_89_valid_1 : _GEN_604; // @[ICache.scala 132:{59,59}]
  wire  _GEN_606 = 7'h5a == _GEN_13517 ? meta_90_valid_1 : _GEN_605; // @[ICache.scala 132:{59,59}]
  wire  _GEN_607 = 7'h5b == _GEN_13517 ? meta_91_valid_1 : _GEN_606; // @[ICache.scala 132:{59,59}]
  wire  _GEN_608 = 7'h5c == _GEN_13517 ? meta_92_valid_1 : _GEN_607; // @[ICache.scala 132:{59,59}]
  wire  _GEN_609 = 7'h5d == _GEN_13517 ? meta_93_valid_1 : _GEN_608; // @[ICache.scala 132:{59,59}]
  wire  _GEN_610 = 7'h5e == _GEN_13517 ? meta_94_valid_1 : _GEN_609; // @[ICache.scala 132:{59,59}]
  wire  _GEN_611 = 7'h5f == _GEN_13517 ? meta_95_valid_1 : _GEN_610; // @[ICache.scala 132:{59,59}]
  wire  _GEN_612 = 7'h60 == _GEN_13517 ? meta_96_valid_1 : _GEN_611; // @[ICache.scala 132:{59,59}]
  wire  _GEN_613 = 7'h61 == _GEN_13517 ? meta_97_valid_1 : _GEN_612; // @[ICache.scala 132:{59,59}]
  wire  _GEN_614 = 7'h62 == _GEN_13517 ? meta_98_valid_1 : _GEN_613; // @[ICache.scala 132:{59,59}]
  wire  _GEN_615 = 7'h63 == _GEN_13517 ? meta_99_valid_1 : _GEN_614; // @[ICache.scala 132:{59,59}]
  wire  _GEN_616 = 7'h64 == _GEN_13517 ? meta_100_valid_1 : _GEN_615; // @[ICache.scala 132:{59,59}]
  wire  _GEN_617 = 7'h65 == _GEN_13517 ? meta_101_valid_1 : _GEN_616; // @[ICache.scala 132:{59,59}]
  wire  _GEN_618 = 7'h66 == _GEN_13517 ? meta_102_valid_1 : _GEN_617; // @[ICache.scala 132:{59,59}]
  wire  _GEN_619 = 7'h67 == _GEN_13517 ? meta_103_valid_1 : _GEN_618; // @[ICache.scala 132:{59,59}]
  wire  _GEN_620 = 7'h68 == _GEN_13517 ? meta_104_valid_1 : _GEN_619; // @[ICache.scala 132:{59,59}]
  wire  _GEN_621 = 7'h69 == _GEN_13517 ? meta_105_valid_1 : _GEN_620; // @[ICache.scala 132:{59,59}]
  wire  _GEN_622 = 7'h6a == _GEN_13517 ? meta_106_valid_1 : _GEN_621; // @[ICache.scala 132:{59,59}]
  wire  _GEN_623 = 7'h6b == _GEN_13517 ? meta_107_valid_1 : _GEN_622; // @[ICache.scala 132:{59,59}]
  wire  _GEN_624 = 7'h6c == _GEN_13517 ? meta_108_valid_1 : _GEN_623; // @[ICache.scala 132:{59,59}]
  wire  _GEN_625 = 7'h6d == _GEN_13517 ? meta_109_valid_1 : _GEN_624; // @[ICache.scala 132:{59,59}]
  wire  _GEN_626 = 7'h6e == _GEN_13517 ? meta_110_valid_1 : _GEN_625; // @[ICache.scala 132:{59,59}]
  wire  _GEN_627 = 7'h6f == _GEN_13517 ? meta_111_valid_1 : _GEN_626; // @[ICache.scala 132:{59,59}]
  wire  _GEN_628 = 7'h70 == _GEN_13517 ? meta_112_valid_1 : _GEN_627; // @[ICache.scala 132:{59,59}]
  wire  _GEN_629 = 7'h71 == _GEN_13517 ? meta_113_valid_1 : _GEN_628; // @[ICache.scala 132:{59,59}]
  wire  _GEN_630 = 7'h72 == _GEN_13517 ? meta_114_valid_1 : _GEN_629; // @[ICache.scala 132:{59,59}]
  wire  _GEN_631 = 7'h73 == _GEN_13517 ? meta_115_valid_1 : _GEN_630; // @[ICache.scala 132:{59,59}]
  wire  _GEN_632 = 7'h74 == _GEN_13517 ? meta_116_valid_1 : _GEN_631; // @[ICache.scala 132:{59,59}]
  wire  _GEN_633 = 7'h75 == _GEN_13517 ? meta_117_valid_1 : _GEN_632; // @[ICache.scala 132:{59,59}]
  wire  _GEN_634 = 7'h76 == _GEN_13517 ? meta_118_valid_1 : _GEN_633; // @[ICache.scala 132:{59,59}]
  wire  _GEN_635 = 7'h77 == _GEN_13517 ? meta_119_valid_1 : _GEN_634; // @[ICache.scala 132:{59,59}]
  wire  _GEN_636 = 7'h78 == _GEN_13517 ? meta_120_valid_1 : _GEN_635; // @[ICache.scala 132:{59,59}]
  wire  _GEN_637 = 7'h79 == _GEN_13517 ? meta_121_valid_1 : _GEN_636; // @[ICache.scala 132:{59,59}]
  wire  _GEN_638 = 7'h7a == _GEN_13517 ? meta_122_valid_1 : _GEN_637; // @[ICache.scala 132:{59,59}]
  wire  _GEN_639 = 7'h7b == _GEN_13517 ? meta_123_valid_1 : _GEN_638; // @[ICache.scala 132:{59,59}]
  wire  _GEN_640 = 7'h7c == _GEN_13517 ? meta_124_valid_1 : _GEN_639; // @[ICache.scala 132:{59,59}]
  wire  _GEN_641 = 7'h7d == _GEN_13517 ? meta_125_valid_1 : _GEN_640; // @[ICache.scala 132:{59,59}]
  wire  _GEN_642 = 7'h7e == _GEN_13517 ? meta_126_valid_1 : _GEN_641; // @[ICache.scala 132:{59,59}]
  wire  _GEN_643 = 7'h7f == _GEN_13517 ? meta_127_valid_1 : _GEN_642; // @[ICache.scala 132:{59,59}]
  wire  _GEN_644 = 8'h80 == _GEN_13581 ? meta_128_valid_1 : _GEN_643; // @[ICache.scala 132:{59,59}]
  wire  _GEN_645 = 8'h81 == _GEN_13581 ? meta_129_valid_1 : _GEN_644; // @[ICache.scala 132:{59,59}]
  wire  _GEN_646 = 8'h82 == _GEN_13581 ? meta_130_valid_1 : _GEN_645; // @[ICache.scala 132:{59,59}]
  wire  _GEN_647 = 8'h83 == _GEN_13581 ? meta_131_valid_1 : _GEN_646; // @[ICache.scala 132:{59,59}]
  wire  _GEN_648 = 8'h84 == _GEN_13581 ? meta_132_valid_1 : _GEN_647; // @[ICache.scala 132:{59,59}]
  wire  _GEN_649 = 8'h85 == _GEN_13581 ? meta_133_valid_1 : _GEN_648; // @[ICache.scala 132:{59,59}]
  wire  _GEN_650 = 8'h86 == _GEN_13581 ? meta_134_valid_1 : _GEN_649; // @[ICache.scala 132:{59,59}]
  wire  _GEN_651 = 8'h87 == _GEN_13581 ? meta_135_valid_1 : _GEN_650; // @[ICache.scala 132:{59,59}]
  wire  _GEN_652 = 8'h88 == _GEN_13581 ? meta_136_valid_1 : _GEN_651; // @[ICache.scala 132:{59,59}]
  wire  _GEN_653 = 8'h89 == _GEN_13581 ? meta_137_valid_1 : _GEN_652; // @[ICache.scala 132:{59,59}]
  wire  _GEN_654 = 8'h8a == _GEN_13581 ? meta_138_valid_1 : _GEN_653; // @[ICache.scala 132:{59,59}]
  wire  _GEN_655 = 8'h8b == _GEN_13581 ? meta_139_valid_1 : _GEN_654; // @[ICache.scala 132:{59,59}]
  wire  _GEN_656 = 8'h8c == _GEN_13581 ? meta_140_valid_1 : _GEN_655; // @[ICache.scala 132:{59,59}]
  wire  _GEN_657 = 8'h8d == _GEN_13581 ? meta_141_valid_1 : _GEN_656; // @[ICache.scala 132:{59,59}]
  wire  _GEN_658 = 8'h8e == _GEN_13581 ? meta_142_valid_1 : _GEN_657; // @[ICache.scala 132:{59,59}]
  wire  _GEN_659 = 8'h8f == _GEN_13581 ? meta_143_valid_1 : _GEN_658; // @[ICache.scala 132:{59,59}]
  wire  _GEN_660 = 8'h90 == _GEN_13581 ? meta_144_valid_1 : _GEN_659; // @[ICache.scala 132:{59,59}]
  wire  _GEN_661 = 8'h91 == _GEN_13581 ? meta_145_valid_1 : _GEN_660; // @[ICache.scala 132:{59,59}]
  wire  _GEN_662 = 8'h92 == _GEN_13581 ? meta_146_valid_1 : _GEN_661; // @[ICache.scala 132:{59,59}]
  wire  _GEN_663 = 8'h93 == _GEN_13581 ? meta_147_valid_1 : _GEN_662; // @[ICache.scala 132:{59,59}]
  wire  _GEN_664 = 8'h94 == _GEN_13581 ? meta_148_valid_1 : _GEN_663; // @[ICache.scala 132:{59,59}]
  wire  _GEN_665 = 8'h95 == _GEN_13581 ? meta_149_valid_1 : _GEN_664; // @[ICache.scala 132:{59,59}]
  wire  _GEN_666 = 8'h96 == _GEN_13581 ? meta_150_valid_1 : _GEN_665; // @[ICache.scala 132:{59,59}]
  wire  _GEN_667 = 8'h97 == _GEN_13581 ? meta_151_valid_1 : _GEN_666; // @[ICache.scala 132:{59,59}]
  wire  _GEN_668 = 8'h98 == _GEN_13581 ? meta_152_valid_1 : _GEN_667; // @[ICache.scala 132:{59,59}]
  wire  _GEN_669 = 8'h99 == _GEN_13581 ? meta_153_valid_1 : _GEN_668; // @[ICache.scala 132:{59,59}]
  wire  _GEN_670 = 8'h9a == _GEN_13581 ? meta_154_valid_1 : _GEN_669; // @[ICache.scala 132:{59,59}]
  wire  _GEN_671 = 8'h9b == _GEN_13581 ? meta_155_valid_1 : _GEN_670; // @[ICache.scala 132:{59,59}]
  wire  _GEN_672 = 8'h9c == _GEN_13581 ? meta_156_valid_1 : _GEN_671; // @[ICache.scala 132:{59,59}]
  wire  _GEN_673 = 8'h9d == _GEN_13581 ? meta_157_valid_1 : _GEN_672; // @[ICache.scala 132:{59,59}]
  wire  _GEN_674 = 8'h9e == _GEN_13581 ? meta_158_valid_1 : _GEN_673; // @[ICache.scala 132:{59,59}]
  wire  _GEN_675 = 8'h9f == _GEN_13581 ? meta_159_valid_1 : _GEN_674; // @[ICache.scala 132:{59,59}]
  wire  _GEN_676 = 8'ha0 == _GEN_13581 ? meta_160_valid_1 : _GEN_675; // @[ICache.scala 132:{59,59}]
  wire  _GEN_677 = 8'ha1 == _GEN_13581 ? meta_161_valid_1 : _GEN_676; // @[ICache.scala 132:{59,59}]
  wire  _GEN_678 = 8'ha2 == _GEN_13581 ? meta_162_valid_1 : _GEN_677; // @[ICache.scala 132:{59,59}]
  wire  _GEN_679 = 8'ha3 == _GEN_13581 ? meta_163_valid_1 : _GEN_678; // @[ICache.scala 132:{59,59}]
  wire  _GEN_680 = 8'ha4 == _GEN_13581 ? meta_164_valid_1 : _GEN_679; // @[ICache.scala 132:{59,59}]
  wire  _GEN_681 = 8'ha5 == _GEN_13581 ? meta_165_valid_1 : _GEN_680; // @[ICache.scala 132:{59,59}]
  wire  _GEN_682 = 8'ha6 == _GEN_13581 ? meta_166_valid_1 : _GEN_681; // @[ICache.scala 132:{59,59}]
  wire  _GEN_683 = 8'ha7 == _GEN_13581 ? meta_167_valid_1 : _GEN_682; // @[ICache.scala 132:{59,59}]
  wire  _GEN_684 = 8'ha8 == _GEN_13581 ? meta_168_valid_1 : _GEN_683; // @[ICache.scala 132:{59,59}]
  wire  _GEN_685 = 8'ha9 == _GEN_13581 ? meta_169_valid_1 : _GEN_684; // @[ICache.scala 132:{59,59}]
  wire  _GEN_686 = 8'haa == _GEN_13581 ? meta_170_valid_1 : _GEN_685; // @[ICache.scala 132:{59,59}]
  wire  _GEN_687 = 8'hab == _GEN_13581 ? meta_171_valid_1 : _GEN_686; // @[ICache.scala 132:{59,59}]
  wire  _GEN_688 = 8'hac == _GEN_13581 ? meta_172_valid_1 : _GEN_687; // @[ICache.scala 132:{59,59}]
  wire  _GEN_689 = 8'had == _GEN_13581 ? meta_173_valid_1 : _GEN_688; // @[ICache.scala 132:{59,59}]
  wire  _GEN_690 = 8'hae == _GEN_13581 ? meta_174_valid_1 : _GEN_689; // @[ICache.scala 132:{59,59}]
  wire  _GEN_691 = 8'haf == _GEN_13581 ? meta_175_valid_1 : _GEN_690; // @[ICache.scala 132:{59,59}]
  wire  _GEN_692 = 8'hb0 == _GEN_13581 ? meta_176_valid_1 : _GEN_691; // @[ICache.scala 132:{59,59}]
  wire  _GEN_693 = 8'hb1 == _GEN_13581 ? meta_177_valid_1 : _GEN_692; // @[ICache.scala 132:{59,59}]
  wire  _GEN_694 = 8'hb2 == _GEN_13581 ? meta_178_valid_1 : _GEN_693; // @[ICache.scala 132:{59,59}]
  wire  _GEN_695 = 8'hb3 == _GEN_13581 ? meta_179_valid_1 : _GEN_694; // @[ICache.scala 132:{59,59}]
  wire  _GEN_696 = 8'hb4 == _GEN_13581 ? meta_180_valid_1 : _GEN_695; // @[ICache.scala 132:{59,59}]
  wire  _GEN_697 = 8'hb5 == _GEN_13581 ? meta_181_valid_1 : _GEN_696; // @[ICache.scala 132:{59,59}]
  wire  _GEN_698 = 8'hb6 == _GEN_13581 ? meta_182_valid_1 : _GEN_697; // @[ICache.scala 132:{59,59}]
  wire  _GEN_699 = 8'hb7 == _GEN_13581 ? meta_183_valid_1 : _GEN_698; // @[ICache.scala 132:{59,59}]
  wire  _GEN_700 = 8'hb8 == _GEN_13581 ? meta_184_valid_1 : _GEN_699; // @[ICache.scala 132:{59,59}]
  wire  _GEN_701 = 8'hb9 == _GEN_13581 ? meta_185_valid_1 : _GEN_700; // @[ICache.scala 132:{59,59}]
  wire  _GEN_702 = 8'hba == _GEN_13581 ? meta_186_valid_1 : _GEN_701; // @[ICache.scala 132:{59,59}]
  wire  _GEN_703 = 8'hbb == _GEN_13581 ? meta_187_valid_1 : _GEN_702; // @[ICache.scala 132:{59,59}]
  wire  _GEN_704 = 8'hbc == _GEN_13581 ? meta_188_valid_1 : _GEN_703; // @[ICache.scala 132:{59,59}]
  wire  _GEN_705 = 8'hbd == _GEN_13581 ? meta_189_valid_1 : _GEN_704; // @[ICache.scala 132:{59,59}]
  wire  _GEN_706 = 8'hbe == _GEN_13581 ? meta_190_valid_1 : _GEN_705; // @[ICache.scala 132:{59,59}]
  wire  _GEN_707 = 8'hbf == _GEN_13581 ? meta_191_valid_1 : _GEN_706; // @[ICache.scala 132:{59,59}]
  wire  _GEN_708 = 8'hc0 == _GEN_13581 ? meta_192_valid_1 : _GEN_707; // @[ICache.scala 132:{59,59}]
  wire  _GEN_709 = 8'hc1 == _GEN_13581 ? meta_193_valid_1 : _GEN_708; // @[ICache.scala 132:{59,59}]
  wire  _GEN_710 = 8'hc2 == _GEN_13581 ? meta_194_valid_1 : _GEN_709; // @[ICache.scala 132:{59,59}]
  wire  _GEN_711 = 8'hc3 == _GEN_13581 ? meta_195_valid_1 : _GEN_710; // @[ICache.scala 132:{59,59}]
  wire  _GEN_712 = 8'hc4 == _GEN_13581 ? meta_196_valid_1 : _GEN_711; // @[ICache.scala 132:{59,59}]
  wire  _GEN_713 = 8'hc5 == _GEN_13581 ? meta_197_valid_1 : _GEN_712; // @[ICache.scala 132:{59,59}]
  wire  _GEN_714 = 8'hc6 == _GEN_13581 ? meta_198_valid_1 : _GEN_713; // @[ICache.scala 132:{59,59}]
  wire  _GEN_715 = 8'hc7 == _GEN_13581 ? meta_199_valid_1 : _GEN_714; // @[ICache.scala 132:{59,59}]
  wire  _GEN_716 = 8'hc8 == _GEN_13581 ? meta_200_valid_1 : _GEN_715; // @[ICache.scala 132:{59,59}]
  wire  _GEN_717 = 8'hc9 == _GEN_13581 ? meta_201_valid_1 : _GEN_716; // @[ICache.scala 132:{59,59}]
  wire  _GEN_718 = 8'hca == _GEN_13581 ? meta_202_valid_1 : _GEN_717; // @[ICache.scala 132:{59,59}]
  wire  _GEN_719 = 8'hcb == _GEN_13581 ? meta_203_valid_1 : _GEN_718; // @[ICache.scala 132:{59,59}]
  wire  _GEN_720 = 8'hcc == _GEN_13581 ? meta_204_valid_1 : _GEN_719; // @[ICache.scala 132:{59,59}]
  wire  _GEN_721 = 8'hcd == _GEN_13581 ? meta_205_valid_1 : _GEN_720; // @[ICache.scala 132:{59,59}]
  wire  _GEN_722 = 8'hce == _GEN_13581 ? meta_206_valid_1 : _GEN_721; // @[ICache.scala 132:{59,59}]
  wire  _GEN_723 = 8'hcf == _GEN_13581 ? meta_207_valid_1 : _GEN_722; // @[ICache.scala 132:{59,59}]
  wire  _GEN_724 = 8'hd0 == _GEN_13581 ? meta_208_valid_1 : _GEN_723; // @[ICache.scala 132:{59,59}]
  wire  _GEN_725 = 8'hd1 == _GEN_13581 ? meta_209_valid_1 : _GEN_724; // @[ICache.scala 132:{59,59}]
  wire  _GEN_726 = 8'hd2 == _GEN_13581 ? meta_210_valid_1 : _GEN_725; // @[ICache.scala 132:{59,59}]
  wire  _GEN_727 = 8'hd3 == _GEN_13581 ? meta_211_valid_1 : _GEN_726; // @[ICache.scala 132:{59,59}]
  wire  _GEN_728 = 8'hd4 == _GEN_13581 ? meta_212_valid_1 : _GEN_727; // @[ICache.scala 132:{59,59}]
  wire  _GEN_729 = 8'hd5 == _GEN_13581 ? meta_213_valid_1 : _GEN_728; // @[ICache.scala 132:{59,59}]
  wire  _GEN_730 = 8'hd6 == _GEN_13581 ? meta_214_valid_1 : _GEN_729; // @[ICache.scala 132:{59,59}]
  wire  _GEN_731 = 8'hd7 == _GEN_13581 ? meta_215_valid_1 : _GEN_730; // @[ICache.scala 132:{59,59}]
  wire  _GEN_732 = 8'hd8 == _GEN_13581 ? meta_216_valid_1 : _GEN_731; // @[ICache.scala 132:{59,59}]
  wire  _GEN_733 = 8'hd9 == _GEN_13581 ? meta_217_valid_1 : _GEN_732; // @[ICache.scala 132:{59,59}]
  wire  _GEN_734 = 8'hda == _GEN_13581 ? meta_218_valid_1 : _GEN_733; // @[ICache.scala 132:{59,59}]
  wire  _GEN_735 = 8'hdb == _GEN_13581 ? meta_219_valid_1 : _GEN_734; // @[ICache.scala 132:{59,59}]
  wire  _GEN_736 = 8'hdc == _GEN_13581 ? meta_220_valid_1 : _GEN_735; // @[ICache.scala 132:{59,59}]
  wire  _GEN_737 = 8'hdd == _GEN_13581 ? meta_221_valid_1 : _GEN_736; // @[ICache.scala 132:{59,59}]
  wire  _GEN_738 = 8'hde == _GEN_13581 ? meta_222_valid_1 : _GEN_737; // @[ICache.scala 132:{59,59}]
  wire  _GEN_739 = 8'hdf == _GEN_13581 ? meta_223_valid_1 : _GEN_738; // @[ICache.scala 132:{59,59}]
  wire  _GEN_740 = 8'he0 == _GEN_13581 ? meta_224_valid_1 : _GEN_739; // @[ICache.scala 132:{59,59}]
  wire  _GEN_741 = 8'he1 == _GEN_13581 ? meta_225_valid_1 : _GEN_740; // @[ICache.scala 132:{59,59}]
  wire  _GEN_742 = 8'he2 == _GEN_13581 ? meta_226_valid_1 : _GEN_741; // @[ICache.scala 132:{59,59}]
  wire  _GEN_743 = 8'he3 == _GEN_13581 ? meta_227_valid_1 : _GEN_742; // @[ICache.scala 132:{59,59}]
  wire  _GEN_744 = 8'he4 == _GEN_13581 ? meta_228_valid_1 : _GEN_743; // @[ICache.scala 132:{59,59}]
  wire  _GEN_745 = 8'he5 == _GEN_13581 ? meta_229_valid_1 : _GEN_744; // @[ICache.scala 132:{59,59}]
  wire  _GEN_746 = 8'he6 == _GEN_13581 ? meta_230_valid_1 : _GEN_745; // @[ICache.scala 132:{59,59}]
  wire  _GEN_747 = 8'he7 == _GEN_13581 ? meta_231_valid_1 : _GEN_746; // @[ICache.scala 132:{59,59}]
  wire  _GEN_748 = 8'he8 == _GEN_13581 ? meta_232_valid_1 : _GEN_747; // @[ICache.scala 132:{59,59}]
  wire  _GEN_749 = 8'he9 == _GEN_13581 ? meta_233_valid_1 : _GEN_748; // @[ICache.scala 132:{59,59}]
  wire  _GEN_750 = 8'hea == _GEN_13581 ? meta_234_valid_1 : _GEN_749; // @[ICache.scala 132:{59,59}]
  wire  _GEN_751 = 8'heb == _GEN_13581 ? meta_235_valid_1 : _GEN_750; // @[ICache.scala 132:{59,59}]
  wire  _GEN_752 = 8'hec == _GEN_13581 ? meta_236_valid_1 : _GEN_751; // @[ICache.scala 132:{59,59}]
  wire  _GEN_753 = 8'hed == _GEN_13581 ? meta_237_valid_1 : _GEN_752; // @[ICache.scala 132:{59,59}]
  wire  _GEN_754 = 8'hee == _GEN_13581 ? meta_238_valid_1 : _GEN_753; // @[ICache.scala 132:{59,59}]
  wire  _GEN_755 = 8'hef == _GEN_13581 ? meta_239_valid_1 : _GEN_754; // @[ICache.scala 132:{59,59}]
  wire  _GEN_756 = 8'hf0 == _GEN_13581 ? meta_240_valid_1 : _GEN_755; // @[ICache.scala 132:{59,59}]
  wire  _GEN_757 = 8'hf1 == _GEN_13581 ? meta_241_valid_1 : _GEN_756; // @[ICache.scala 132:{59,59}]
  wire  _GEN_758 = 8'hf2 == _GEN_13581 ? meta_242_valid_1 : _GEN_757; // @[ICache.scala 132:{59,59}]
  wire  _GEN_759 = 8'hf3 == _GEN_13581 ? meta_243_valid_1 : _GEN_758; // @[ICache.scala 132:{59,59}]
  wire  _GEN_760 = 8'hf4 == _GEN_13581 ? meta_244_valid_1 : _GEN_759; // @[ICache.scala 132:{59,59}]
  wire  _GEN_761 = 8'hf5 == _GEN_13581 ? meta_245_valid_1 : _GEN_760; // @[ICache.scala 132:{59,59}]
  wire  _GEN_762 = 8'hf6 == _GEN_13581 ? meta_246_valid_1 : _GEN_761; // @[ICache.scala 132:{59,59}]
  wire  _GEN_763 = 8'hf7 == _GEN_13581 ? meta_247_valid_1 : _GEN_762; // @[ICache.scala 132:{59,59}]
  wire  _GEN_764 = 8'hf8 == _GEN_13581 ? meta_248_valid_1 : _GEN_763; // @[ICache.scala 132:{59,59}]
  wire  _GEN_765 = 8'hf9 == _GEN_13581 ? meta_249_valid_1 : _GEN_764; // @[ICache.scala 132:{59,59}]
  wire  _GEN_766 = 8'hfa == _GEN_13581 ? meta_250_valid_1 : _GEN_765; // @[ICache.scala 132:{59,59}]
  wire  _GEN_767 = 8'hfb == _GEN_13581 ? meta_251_valid_1 : _GEN_766; // @[ICache.scala 132:{59,59}]
  wire  _GEN_768 = 8'hfc == _GEN_13581 ? meta_252_valid_1 : _GEN_767; // @[ICache.scala 132:{59,59}]
  wire  _GEN_769 = 8'hfd == _GEN_13581 ? meta_253_valid_1 : _GEN_768; // @[ICache.scala 132:{59,59}]
  wire  _GEN_770 = 8'hfe == _GEN_13581 ? meta_254_valid_1 : _GEN_769; // @[ICache.scala 132:{59,59}]
  wire  _GEN_771 = 8'hff == _GEN_13581 ? meta_255_valid_1 : _GEN_770; // @[ICache.scala 132:{59,59}]
  wire  _GEN_772 = 9'h100 == _GEN_13709 ? meta_256_valid_1 : _GEN_771; // @[ICache.scala 132:{59,59}]
  wire  _GEN_773 = 9'h101 == _GEN_13709 ? meta_257_valid_1 : _GEN_772; // @[ICache.scala 132:{59,59}]
  wire  _GEN_774 = 9'h102 == _GEN_13709 ? meta_258_valid_1 : _GEN_773; // @[ICache.scala 132:{59,59}]
  wire  _GEN_775 = 9'h103 == _GEN_13709 ? meta_259_valid_1 : _GEN_774; // @[ICache.scala 132:{59,59}]
  wire  _GEN_776 = 9'h104 == _GEN_13709 ? meta_260_valid_1 : _GEN_775; // @[ICache.scala 132:{59,59}]
  wire  _GEN_777 = 9'h105 == _GEN_13709 ? meta_261_valid_1 : _GEN_776; // @[ICache.scala 132:{59,59}]
  wire  _GEN_778 = 9'h106 == _GEN_13709 ? meta_262_valid_1 : _GEN_777; // @[ICache.scala 132:{59,59}]
  wire  _GEN_779 = 9'h107 == _GEN_13709 ? meta_263_valid_1 : _GEN_778; // @[ICache.scala 132:{59,59}]
  wire  _GEN_780 = 9'h108 == _GEN_13709 ? meta_264_valid_1 : _GEN_779; // @[ICache.scala 132:{59,59}]
  wire  _GEN_781 = 9'h109 == _GEN_13709 ? meta_265_valid_1 : _GEN_780; // @[ICache.scala 132:{59,59}]
  wire  _GEN_782 = 9'h10a == _GEN_13709 ? meta_266_valid_1 : _GEN_781; // @[ICache.scala 132:{59,59}]
  wire  _GEN_783 = 9'h10b == _GEN_13709 ? meta_267_valid_1 : _GEN_782; // @[ICache.scala 132:{59,59}]
  wire  _GEN_784 = 9'h10c == _GEN_13709 ? meta_268_valid_1 : _GEN_783; // @[ICache.scala 132:{59,59}]
  wire  _GEN_785 = 9'h10d == _GEN_13709 ? meta_269_valid_1 : _GEN_784; // @[ICache.scala 132:{59,59}]
  wire  _GEN_786 = 9'h10e == _GEN_13709 ? meta_270_valid_1 : _GEN_785; // @[ICache.scala 132:{59,59}]
  wire  _GEN_787 = 9'h10f == _GEN_13709 ? meta_271_valid_1 : _GEN_786; // @[ICache.scala 132:{59,59}]
  wire  _GEN_788 = 9'h110 == _GEN_13709 ? meta_272_valid_1 : _GEN_787; // @[ICache.scala 132:{59,59}]
  wire  _GEN_789 = 9'h111 == _GEN_13709 ? meta_273_valid_1 : _GEN_788; // @[ICache.scala 132:{59,59}]
  wire  _GEN_790 = 9'h112 == _GEN_13709 ? meta_274_valid_1 : _GEN_789; // @[ICache.scala 132:{59,59}]
  wire  _GEN_791 = 9'h113 == _GEN_13709 ? meta_275_valid_1 : _GEN_790; // @[ICache.scala 132:{59,59}]
  wire  _GEN_792 = 9'h114 == _GEN_13709 ? meta_276_valid_1 : _GEN_791; // @[ICache.scala 132:{59,59}]
  wire  _GEN_793 = 9'h115 == _GEN_13709 ? meta_277_valid_1 : _GEN_792; // @[ICache.scala 132:{59,59}]
  wire  _GEN_794 = 9'h116 == _GEN_13709 ? meta_278_valid_1 : _GEN_793; // @[ICache.scala 132:{59,59}]
  wire  _GEN_795 = 9'h117 == _GEN_13709 ? meta_279_valid_1 : _GEN_794; // @[ICache.scala 132:{59,59}]
  wire  _GEN_796 = 9'h118 == _GEN_13709 ? meta_280_valid_1 : _GEN_795; // @[ICache.scala 132:{59,59}]
  wire  _GEN_797 = 9'h119 == _GEN_13709 ? meta_281_valid_1 : _GEN_796; // @[ICache.scala 132:{59,59}]
  wire  _GEN_798 = 9'h11a == _GEN_13709 ? meta_282_valid_1 : _GEN_797; // @[ICache.scala 132:{59,59}]
  wire  _GEN_799 = 9'h11b == _GEN_13709 ? meta_283_valid_1 : _GEN_798; // @[ICache.scala 132:{59,59}]
  wire  _GEN_800 = 9'h11c == _GEN_13709 ? meta_284_valid_1 : _GEN_799; // @[ICache.scala 132:{59,59}]
  wire  _GEN_801 = 9'h11d == _GEN_13709 ? meta_285_valid_1 : _GEN_800; // @[ICache.scala 132:{59,59}]
  wire  _GEN_802 = 9'h11e == _GEN_13709 ? meta_286_valid_1 : _GEN_801; // @[ICache.scala 132:{59,59}]
  wire  _GEN_803 = 9'h11f == _GEN_13709 ? meta_287_valid_1 : _GEN_802; // @[ICache.scala 132:{59,59}]
  wire  _GEN_804 = 9'h120 == _GEN_13709 ? meta_288_valid_1 : _GEN_803; // @[ICache.scala 132:{59,59}]
  wire  _GEN_805 = 9'h121 == _GEN_13709 ? meta_289_valid_1 : _GEN_804; // @[ICache.scala 132:{59,59}]
  wire  _GEN_806 = 9'h122 == _GEN_13709 ? meta_290_valid_1 : _GEN_805; // @[ICache.scala 132:{59,59}]
  wire  _GEN_807 = 9'h123 == _GEN_13709 ? meta_291_valid_1 : _GEN_806; // @[ICache.scala 132:{59,59}]
  wire  _GEN_808 = 9'h124 == _GEN_13709 ? meta_292_valid_1 : _GEN_807; // @[ICache.scala 132:{59,59}]
  wire  _GEN_809 = 9'h125 == _GEN_13709 ? meta_293_valid_1 : _GEN_808; // @[ICache.scala 132:{59,59}]
  wire  _GEN_810 = 9'h126 == _GEN_13709 ? meta_294_valid_1 : _GEN_809; // @[ICache.scala 132:{59,59}]
  wire  _GEN_811 = 9'h127 == _GEN_13709 ? meta_295_valid_1 : _GEN_810; // @[ICache.scala 132:{59,59}]
  wire  _GEN_812 = 9'h128 == _GEN_13709 ? meta_296_valid_1 : _GEN_811; // @[ICache.scala 132:{59,59}]
  wire  _GEN_813 = 9'h129 == _GEN_13709 ? meta_297_valid_1 : _GEN_812; // @[ICache.scala 132:{59,59}]
  wire  _GEN_814 = 9'h12a == _GEN_13709 ? meta_298_valid_1 : _GEN_813; // @[ICache.scala 132:{59,59}]
  wire  _GEN_815 = 9'h12b == _GEN_13709 ? meta_299_valid_1 : _GEN_814; // @[ICache.scala 132:{59,59}]
  wire  _GEN_816 = 9'h12c == _GEN_13709 ? meta_300_valid_1 : _GEN_815; // @[ICache.scala 132:{59,59}]
  wire  _GEN_817 = 9'h12d == _GEN_13709 ? meta_301_valid_1 : _GEN_816; // @[ICache.scala 132:{59,59}]
  wire  _GEN_818 = 9'h12e == _GEN_13709 ? meta_302_valid_1 : _GEN_817; // @[ICache.scala 132:{59,59}]
  wire  _GEN_819 = 9'h12f == _GEN_13709 ? meta_303_valid_1 : _GEN_818; // @[ICache.scala 132:{59,59}]
  wire  _GEN_820 = 9'h130 == _GEN_13709 ? meta_304_valid_1 : _GEN_819; // @[ICache.scala 132:{59,59}]
  wire  _GEN_821 = 9'h131 == _GEN_13709 ? meta_305_valid_1 : _GEN_820; // @[ICache.scala 132:{59,59}]
  wire  _GEN_822 = 9'h132 == _GEN_13709 ? meta_306_valid_1 : _GEN_821; // @[ICache.scala 132:{59,59}]
  wire  _GEN_823 = 9'h133 == _GEN_13709 ? meta_307_valid_1 : _GEN_822; // @[ICache.scala 132:{59,59}]
  wire  _GEN_824 = 9'h134 == _GEN_13709 ? meta_308_valid_1 : _GEN_823; // @[ICache.scala 132:{59,59}]
  wire  _GEN_825 = 9'h135 == _GEN_13709 ? meta_309_valid_1 : _GEN_824; // @[ICache.scala 132:{59,59}]
  wire  _GEN_826 = 9'h136 == _GEN_13709 ? meta_310_valid_1 : _GEN_825; // @[ICache.scala 132:{59,59}]
  wire  _GEN_827 = 9'h137 == _GEN_13709 ? meta_311_valid_1 : _GEN_826; // @[ICache.scala 132:{59,59}]
  wire  _GEN_828 = 9'h138 == _GEN_13709 ? meta_312_valid_1 : _GEN_827; // @[ICache.scala 132:{59,59}]
  wire  _GEN_829 = 9'h139 == _GEN_13709 ? meta_313_valid_1 : _GEN_828; // @[ICache.scala 132:{59,59}]
  wire  _GEN_830 = 9'h13a == _GEN_13709 ? meta_314_valid_1 : _GEN_829; // @[ICache.scala 132:{59,59}]
  wire  _GEN_831 = 9'h13b == _GEN_13709 ? meta_315_valid_1 : _GEN_830; // @[ICache.scala 132:{59,59}]
  wire  _GEN_832 = 9'h13c == _GEN_13709 ? meta_316_valid_1 : _GEN_831; // @[ICache.scala 132:{59,59}]
  wire  _GEN_833 = 9'h13d == _GEN_13709 ? meta_317_valid_1 : _GEN_832; // @[ICache.scala 132:{59,59}]
  wire  _GEN_834 = 9'h13e == _GEN_13709 ? meta_318_valid_1 : _GEN_833; // @[ICache.scala 132:{59,59}]
  wire  _GEN_835 = 9'h13f == _GEN_13709 ? meta_319_valid_1 : _GEN_834; // @[ICache.scala 132:{59,59}]
  wire  _GEN_836 = 9'h140 == _GEN_13709 ? meta_320_valid_1 : _GEN_835; // @[ICache.scala 132:{59,59}]
  wire  _GEN_837 = 9'h141 == _GEN_13709 ? meta_321_valid_1 : _GEN_836; // @[ICache.scala 132:{59,59}]
  wire  _GEN_838 = 9'h142 == _GEN_13709 ? meta_322_valid_1 : _GEN_837; // @[ICache.scala 132:{59,59}]
  wire  _GEN_839 = 9'h143 == _GEN_13709 ? meta_323_valid_1 : _GEN_838; // @[ICache.scala 132:{59,59}]
  wire  _GEN_840 = 9'h144 == _GEN_13709 ? meta_324_valid_1 : _GEN_839; // @[ICache.scala 132:{59,59}]
  wire  _GEN_841 = 9'h145 == _GEN_13709 ? meta_325_valid_1 : _GEN_840; // @[ICache.scala 132:{59,59}]
  wire  _GEN_842 = 9'h146 == _GEN_13709 ? meta_326_valid_1 : _GEN_841; // @[ICache.scala 132:{59,59}]
  wire  _GEN_843 = 9'h147 == _GEN_13709 ? meta_327_valid_1 : _GEN_842; // @[ICache.scala 132:{59,59}]
  wire  _GEN_844 = 9'h148 == _GEN_13709 ? meta_328_valid_1 : _GEN_843; // @[ICache.scala 132:{59,59}]
  wire  _GEN_845 = 9'h149 == _GEN_13709 ? meta_329_valid_1 : _GEN_844; // @[ICache.scala 132:{59,59}]
  wire  _GEN_846 = 9'h14a == _GEN_13709 ? meta_330_valid_1 : _GEN_845; // @[ICache.scala 132:{59,59}]
  wire  _GEN_847 = 9'h14b == _GEN_13709 ? meta_331_valid_1 : _GEN_846; // @[ICache.scala 132:{59,59}]
  wire  _GEN_848 = 9'h14c == _GEN_13709 ? meta_332_valid_1 : _GEN_847; // @[ICache.scala 132:{59,59}]
  wire  _GEN_849 = 9'h14d == _GEN_13709 ? meta_333_valid_1 : _GEN_848; // @[ICache.scala 132:{59,59}]
  wire  _GEN_850 = 9'h14e == _GEN_13709 ? meta_334_valid_1 : _GEN_849; // @[ICache.scala 132:{59,59}]
  wire  _GEN_851 = 9'h14f == _GEN_13709 ? meta_335_valid_1 : _GEN_850; // @[ICache.scala 132:{59,59}]
  wire  _GEN_852 = 9'h150 == _GEN_13709 ? meta_336_valid_1 : _GEN_851; // @[ICache.scala 132:{59,59}]
  wire  _GEN_853 = 9'h151 == _GEN_13709 ? meta_337_valid_1 : _GEN_852; // @[ICache.scala 132:{59,59}]
  wire  _GEN_854 = 9'h152 == _GEN_13709 ? meta_338_valid_1 : _GEN_853; // @[ICache.scala 132:{59,59}]
  wire  _GEN_855 = 9'h153 == _GEN_13709 ? meta_339_valid_1 : _GEN_854; // @[ICache.scala 132:{59,59}]
  wire  _GEN_856 = 9'h154 == _GEN_13709 ? meta_340_valid_1 : _GEN_855; // @[ICache.scala 132:{59,59}]
  wire  _GEN_857 = 9'h155 == _GEN_13709 ? meta_341_valid_1 : _GEN_856; // @[ICache.scala 132:{59,59}]
  wire  _GEN_858 = 9'h156 == _GEN_13709 ? meta_342_valid_1 : _GEN_857; // @[ICache.scala 132:{59,59}]
  wire  _GEN_859 = 9'h157 == _GEN_13709 ? meta_343_valid_1 : _GEN_858; // @[ICache.scala 132:{59,59}]
  wire  _GEN_860 = 9'h158 == _GEN_13709 ? meta_344_valid_1 : _GEN_859; // @[ICache.scala 132:{59,59}]
  wire  _GEN_861 = 9'h159 == _GEN_13709 ? meta_345_valid_1 : _GEN_860; // @[ICache.scala 132:{59,59}]
  wire  _GEN_862 = 9'h15a == _GEN_13709 ? meta_346_valid_1 : _GEN_861; // @[ICache.scala 132:{59,59}]
  wire  _GEN_863 = 9'h15b == _GEN_13709 ? meta_347_valid_1 : _GEN_862; // @[ICache.scala 132:{59,59}]
  wire  _GEN_864 = 9'h15c == _GEN_13709 ? meta_348_valid_1 : _GEN_863; // @[ICache.scala 132:{59,59}]
  wire  _GEN_865 = 9'h15d == _GEN_13709 ? meta_349_valid_1 : _GEN_864; // @[ICache.scala 132:{59,59}]
  wire  _GEN_866 = 9'h15e == _GEN_13709 ? meta_350_valid_1 : _GEN_865; // @[ICache.scala 132:{59,59}]
  wire  _GEN_867 = 9'h15f == _GEN_13709 ? meta_351_valid_1 : _GEN_866; // @[ICache.scala 132:{59,59}]
  wire  _GEN_868 = 9'h160 == _GEN_13709 ? meta_352_valid_1 : _GEN_867; // @[ICache.scala 132:{59,59}]
  wire  _GEN_869 = 9'h161 == _GEN_13709 ? meta_353_valid_1 : _GEN_868; // @[ICache.scala 132:{59,59}]
  wire  _GEN_870 = 9'h162 == _GEN_13709 ? meta_354_valid_1 : _GEN_869; // @[ICache.scala 132:{59,59}]
  wire  _GEN_871 = 9'h163 == _GEN_13709 ? meta_355_valid_1 : _GEN_870; // @[ICache.scala 132:{59,59}]
  wire  _GEN_872 = 9'h164 == _GEN_13709 ? meta_356_valid_1 : _GEN_871; // @[ICache.scala 132:{59,59}]
  wire  _GEN_873 = 9'h165 == _GEN_13709 ? meta_357_valid_1 : _GEN_872; // @[ICache.scala 132:{59,59}]
  wire  _GEN_874 = 9'h166 == _GEN_13709 ? meta_358_valid_1 : _GEN_873; // @[ICache.scala 132:{59,59}]
  wire  _GEN_875 = 9'h167 == _GEN_13709 ? meta_359_valid_1 : _GEN_874; // @[ICache.scala 132:{59,59}]
  wire  _GEN_876 = 9'h168 == _GEN_13709 ? meta_360_valid_1 : _GEN_875; // @[ICache.scala 132:{59,59}]
  wire  _GEN_877 = 9'h169 == _GEN_13709 ? meta_361_valid_1 : _GEN_876; // @[ICache.scala 132:{59,59}]
  wire  _GEN_878 = 9'h16a == _GEN_13709 ? meta_362_valid_1 : _GEN_877; // @[ICache.scala 132:{59,59}]
  wire  _GEN_879 = 9'h16b == _GEN_13709 ? meta_363_valid_1 : _GEN_878; // @[ICache.scala 132:{59,59}]
  wire  _GEN_880 = 9'h16c == _GEN_13709 ? meta_364_valid_1 : _GEN_879; // @[ICache.scala 132:{59,59}]
  wire  _GEN_881 = 9'h16d == _GEN_13709 ? meta_365_valid_1 : _GEN_880; // @[ICache.scala 132:{59,59}]
  wire  _GEN_882 = 9'h16e == _GEN_13709 ? meta_366_valid_1 : _GEN_881; // @[ICache.scala 132:{59,59}]
  wire  _GEN_883 = 9'h16f == _GEN_13709 ? meta_367_valid_1 : _GEN_882; // @[ICache.scala 132:{59,59}]
  wire  _GEN_884 = 9'h170 == _GEN_13709 ? meta_368_valid_1 : _GEN_883; // @[ICache.scala 132:{59,59}]
  wire  _GEN_885 = 9'h171 == _GEN_13709 ? meta_369_valid_1 : _GEN_884; // @[ICache.scala 132:{59,59}]
  wire  _GEN_886 = 9'h172 == _GEN_13709 ? meta_370_valid_1 : _GEN_885; // @[ICache.scala 132:{59,59}]
  wire  _GEN_887 = 9'h173 == _GEN_13709 ? meta_371_valid_1 : _GEN_886; // @[ICache.scala 132:{59,59}]
  wire  _GEN_888 = 9'h174 == _GEN_13709 ? meta_372_valid_1 : _GEN_887; // @[ICache.scala 132:{59,59}]
  wire  _GEN_889 = 9'h175 == _GEN_13709 ? meta_373_valid_1 : _GEN_888; // @[ICache.scala 132:{59,59}]
  wire  _GEN_890 = 9'h176 == _GEN_13709 ? meta_374_valid_1 : _GEN_889; // @[ICache.scala 132:{59,59}]
  wire  _GEN_891 = 9'h177 == _GEN_13709 ? meta_375_valid_1 : _GEN_890; // @[ICache.scala 132:{59,59}]
  wire  _GEN_892 = 9'h178 == _GEN_13709 ? meta_376_valid_1 : _GEN_891; // @[ICache.scala 132:{59,59}]
  wire  _GEN_893 = 9'h179 == _GEN_13709 ? meta_377_valid_1 : _GEN_892; // @[ICache.scala 132:{59,59}]
  wire  _GEN_894 = 9'h17a == _GEN_13709 ? meta_378_valid_1 : _GEN_893; // @[ICache.scala 132:{59,59}]
  wire  _GEN_895 = 9'h17b == _GEN_13709 ? meta_379_valid_1 : _GEN_894; // @[ICache.scala 132:{59,59}]
  wire  _GEN_896 = 9'h17c == _GEN_13709 ? meta_380_valid_1 : _GEN_895; // @[ICache.scala 132:{59,59}]
  wire  _GEN_897 = 9'h17d == _GEN_13709 ? meta_381_valid_1 : _GEN_896; // @[ICache.scala 132:{59,59}]
  wire  _GEN_898 = 9'h17e == _GEN_13709 ? meta_382_valid_1 : _GEN_897; // @[ICache.scala 132:{59,59}]
  wire  _GEN_899 = 9'h17f == _GEN_13709 ? meta_383_valid_1 : _GEN_898; // @[ICache.scala 132:{59,59}]
  wire  _GEN_900 = 9'h180 == _GEN_13709 ? meta_384_valid_1 : _GEN_899; // @[ICache.scala 132:{59,59}]
  wire  _GEN_901 = 9'h181 == _GEN_13709 ? meta_385_valid_1 : _GEN_900; // @[ICache.scala 132:{59,59}]
  wire  _GEN_902 = 9'h182 == _GEN_13709 ? meta_386_valid_1 : _GEN_901; // @[ICache.scala 132:{59,59}]
  wire  _GEN_903 = 9'h183 == _GEN_13709 ? meta_387_valid_1 : _GEN_902; // @[ICache.scala 132:{59,59}]
  wire  _GEN_904 = 9'h184 == _GEN_13709 ? meta_388_valid_1 : _GEN_903; // @[ICache.scala 132:{59,59}]
  wire  _GEN_905 = 9'h185 == _GEN_13709 ? meta_389_valid_1 : _GEN_904; // @[ICache.scala 132:{59,59}]
  wire  _GEN_906 = 9'h186 == _GEN_13709 ? meta_390_valid_1 : _GEN_905; // @[ICache.scala 132:{59,59}]
  wire  _GEN_907 = 9'h187 == _GEN_13709 ? meta_391_valid_1 : _GEN_906; // @[ICache.scala 132:{59,59}]
  wire  _GEN_908 = 9'h188 == _GEN_13709 ? meta_392_valid_1 : _GEN_907; // @[ICache.scala 132:{59,59}]
  wire  _GEN_909 = 9'h189 == _GEN_13709 ? meta_393_valid_1 : _GEN_908; // @[ICache.scala 132:{59,59}]
  wire  _GEN_910 = 9'h18a == _GEN_13709 ? meta_394_valid_1 : _GEN_909; // @[ICache.scala 132:{59,59}]
  wire  _GEN_911 = 9'h18b == _GEN_13709 ? meta_395_valid_1 : _GEN_910; // @[ICache.scala 132:{59,59}]
  wire  _GEN_912 = 9'h18c == _GEN_13709 ? meta_396_valid_1 : _GEN_911; // @[ICache.scala 132:{59,59}]
  wire  _GEN_913 = 9'h18d == _GEN_13709 ? meta_397_valid_1 : _GEN_912; // @[ICache.scala 132:{59,59}]
  wire  _GEN_914 = 9'h18e == _GEN_13709 ? meta_398_valid_1 : _GEN_913; // @[ICache.scala 132:{59,59}]
  wire  _GEN_915 = 9'h18f == _GEN_13709 ? meta_399_valid_1 : _GEN_914; // @[ICache.scala 132:{59,59}]
  wire  _GEN_916 = 9'h190 == _GEN_13709 ? meta_400_valid_1 : _GEN_915; // @[ICache.scala 132:{59,59}]
  wire  _GEN_917 = 9'h191 == _GEN_13709 ? meta_401_valid_1 : _GEN_916; // @[ICache.scala 132:{59,59}]
  wire  _GEN_918 = 9'h192 == _GEN_13709 ? meta_402_valid_1 : _GEN_917; // @[ICache.scala 132:{59,59}]
  wire  _GEN_919 = 9'h193 == _GEN_13709 ? meta_403_valid_1 : _GEN_918; // @[ICache.scala 132:{59,59}]
  wire  _GEN_920 = 9'h194 == _GEN_13709 ? meta_404_valid_1 : _GEN_919; // @[ICache.scala 132:{59,59}]
  wire  _GEN_921 = 9'h195 == _GEN_13709 ? meta_405_valid_1 : _GEN_920; // @[ICache.scala 132:{59,59}]
  wire  _GEN_922 = 9'h196 == _GEN_13709 ? meta_406_valid_1 : _GEN_921; // @[ICache.scala 132:{59,59}]
  wire  _GEN_923 = 9'h197 == _GEN_13709 ? meta_407_valid_1 : _GEN_922; // @[ICache.scala 132:{59,59}]
  wire  _GEN_924 = 9'h198 == _GEN_13709 ? meta_408_valid_1 : _GEN_923; // @[ICache.scala 132:{59,59}]
  wire  _GEN_925 = 9'h199 == _GEN_13709 ? meta_409_valid_1 : _GEN_924; // @[ICache.scala 132:{59,59}]
  wire  _GEN_926 = 9'h19a == _GEN_13709 ? meta_410_valid_1 : _GEN_925; // @[ICache.scala 132:{59,59}]
  wire  _GEN_927 = 9'h19b == _GEN_13709 ? meta_411_valid_1 : _GEN_926; // @[ICache.scala 132:{59,59}]
  wire  _GEN_928 = 9'h19c == _GEN_13709 ? meta_412_valid_1 : _GEN_927; // @[ICache.scala 132:{59,59}]
  wire  _GEN_929 = 9'h19d == _GEN_13709 ? meta_413_valid_1 : _GEN_928; // @[ICache.scala 132:{59,59}]
  wire  _GEN_930 = 9'h19e == _GEN_13709 ? meta_414_valid_1 : _GEN_929; // @[ICache.scala 132:{59,59}]
  wire  _GEN_931 = 9'h19f == _GEN_13709 ? meta_415_valid_1 : _GEN_930; // @[ICache.scala 132:{59,59}]
  wire  _GEN_932 = 9'h1a0 == _GEN_13709 ? meta_416_valid_1 : _GEN_931; // @[ICache.scala 132:{59,59}]
  wire  _GEN_933 = 9'h1a1 == _GEN_13709 ? meta_417_valid_1 : _GEN_932; // @[ICache.scala 132:{59,59}]
  wire  _GEN_934 = 9'h1a2 == _GEN_13709 ? meta_418_valid_1 : _GEN_933; // @[ICache.scala 132:{59,59}]
  wire  _GEN_935 = 9'h1a3 == _GEN_13709 ? meta_419_valid_1 : _GEN_934; // @[ICache.scala 132:{59,59}]
  wire  _GEN_936 = 9'h1a4 == _GEN_13709 ? meta_420_valid_1 : _GEN_935; // @[ICache.scala 132:{59,59}]
  wire  _GEN_937 = 9'h1a5 == _GEN_13709 ? meta_421_valid_1 : _GEN_936; // @[ICache.scala 132:{59,59}]
  wire  _GEN_938 = 9'h1a6 == _GEN_13709 ? meta_422_valid_1 : _GEN_937; // @[ICache.scala 132:{59,59}]
  wire  _GEN_939 = 9'h1a7 == _GEN_13709 ? meta_423_valid_1 : _GEN_938; // @[ICache.scala 132:{59,59}]
  wire  _GEN_940 = 9'h1a8 == _GEN_13709 ? meta_424_valid_1 : _GEN_939; // @[ICache.scala 132:{59,59}]
  wire  _GEN_941 = 9'h1a9 == _GEN_13709 ? meta_425_valid_1 : _GEN_940; // @[ICache.scala 132:{59,59}]
  wire  _GEN_942 = 9'h1aa == _GEN_13709 ? meta_426_valid_1 : _GEN_941; // @[ICache.scala 132:{59,59}]
  wire  _GEN_943 = 9'h1ab == _GEN_13709 ? meta_427_valid_1 : _GEN_942; // @[ICache.scala 132:{59,59}]
  wire  _GEN_944 = 9'h1ac == _GEN_13709 ? meta_428_valid_1 : _GEN_943; // @[ICache.scala 132:{59,59}]
  wire  _GEN_945 = 9'h1ad == _GEN_13709 ? meta_429_valid_1 : _GEN_944; // @[ICache.scala 132:{59,59}]
  wire  _GEN_946 = 9'h1ae == _GEN_13709 ? meta_430_valid_1 : _GEN_945; // @[ICache.scala 132:{59,59}]
  wire  _GEN_947 = 9'h1af == _GEN_13709 ? meta_431_valid_1 : _GEN_946; // @[ICache.scala 132:{59,59}]
  wire  _GEN_948 = 9'h1b0 == _GEN_13709 ? meta_432_valid_1 : _GEN_947; // @[ICache.scala 132:{59,59}]
  wire  _GEN_949 = 9'h1b1 == _GEN_13709 ? meta_433_valid_1 : _GEN_948; // @[ICache.scala 132:{59,59}]
  wire  _GEN_950 = 9'h1b2 == _GEN_13709 ? meta_434_valid_1 : _GEN_949; // @[ICache.scala 132:{59,59}]
  wire  _GEN_951 = 9'h1b3 == _GEN_13709 ? meta_435_valid_1 : _GEN_950; // @[ICache.scala 132:{59,59}]
  wire  _GEN_952 = 9'h1b4 == _GEN_13709 ? meta_436_valid_1 : _GEN_951; // @[ICache.scala 132:{59,59}]
  wire  _GEN_953 = 9'h1b5 == _GEN_13709 ? meta_437_valid_1 : _GEN_952; // @[ICache.scala 132:{59,59}]
  wire  _GEN_954 = 9'h1b6 == _GEN_13709 ? meta_438_valid_1 : _GEN_953; // @[ICache.scala 132:{59,59}]
  wire  _GEN_955 = 9'h1b7 == _GEN_13709 ? meta_439_valid_1 : _GEN_954; // @[ICache.scala 132:{59,59}]
  wire  _GEN_956 = 9'h1b8 == _GEN_13709 ? meta_440_valid_1 : _GEN_955; // @[ICache.scala 132:{59,59}]
  wire  _GEN_957 = 9'h1b9 == _GEN_13709 ? meta_441_valid_1 : _GEN_956; // @[ICache.scala 132:{59,59}]
  wire  _GEN_958 = 9'h1ba == _GEN_13709 ? meta_442_valid_1 : _GEN_957; // @[ICache.scala 132:{59,59}]
  wire  _GEN_959 = 9'h1bb == _GEN_13709 ? meta_443_valid_1 : _GEN_958; // @[ICache.scala 132:{59,59}]
  wire  _GEN_960 = 9'h1bc == _GEN_13709 ? meta_444_valid_1 : _GEN_959; // @[ICache.scala 132:{59,59}]
  wire  _GEN_961 = 9'h1bd == _GEN_13709 ? meta_445_valid_1 : _GEN_960; // @[ICache.scala 132:{59,59}]
  wire  _GEN_962 = 9'h1be == _GEN_13709 ? meta_446_valid_1 : _GEN_961; // @[ICache.scala 132:{59,59}]
  wire  _GEN_963 = 9'h1bf == _GEN_13709 ? meta_447_valid_1 : _GEN_962; // @[ICache.scala 132:{59,59}]
  wire  _GEN_964 = 9'h1c0 == _GEN_13709 ? meta_448_valid_1 : _GEN_963; // @[ICache.scala 132:{59,59}]
  wire  _GEN_965 = 9'h1c1 == _GEN_13709 ? meta_449_valid_1 : _GEN_964; // @[ICache.scala 132:{59,59}]
  wire  _GEN_966 = 9'h1c2 == _GEN_13709 ? meta_450_valid_1 : _GEN_965; // @[ICache.scala 132:{59,59}]
  wire  _GEN_967 = 9'h1c3 == _GEN_13709 ? meta_451_valid_1 : _GEN_966; // @[ICache.scala 132:{59,59}]
  wire  _GEN_968 = 9'h1c4 == _GEN_13709 ? meta_452_valid_1 : _GEN_967; // @[ICache.scala 132:{59,59}]
  wire  _GEN_969 = 9'h1c5 == _GEN_13709 ? meta_453_valid_1 : _GEN_968; // @[ICache.scala 132:{59,59}]
  wire  _GEN_970 = 9'h1c6 == _GEN_13709 ? meta_454_valid_1 : _GEN_969; // @[ICache.scala 132:{59,59}]
  wire  _GEN_971 = 9'h1c7 == _GEN_13709 ? meta_455_valid_1 : _GEN_970; // @[ICache.scala 132:{59,59}]
  wire  _GEN_972 = 9'h1c8 == _GEN_13709 ? meta_456_valid_1 : _GEN_971; // @[ICache.scala 132:{59,59}]
  wire  _GEN_973 = 9'h1c9 == _GEN_13709 ? meta_457_valid_1 : _GEN_972; // @[ICache.scala 132:{59,59}]
  wire  _GEN_974 = 9'h1ca == _GEN_13709 ? meta_458_valid_1 : _GEN_973; // @[ICache.scala 132:{59,59}]
  wire  _GEN_975 = 9'h1cb == _GEN_13709 ? meta_459_valid_1 : _GEN_974; // @[ICache.scala 132:{59,59}]
  wire  _GEN_976 = 9'h1cc == _GEN_13709 ? meta_460_valid_1 : _GEN_975; // @[ICache.scala 132:{59,59}]
  wire  _GEN_977 = 9'h1cd == _GEN_13709 ? meta_461_valid_1 : _GEN_976; // @[ICache.scala 132:{59,59}]
  wire  _GEN_978 = 9'h1ce == _GEN_13709 ? meta_462_valid_1 : _GEN_977; // @[ICache.scala 132:{59,59}]
  wire  _GEN_979 = 9'h1cf == _GEN_13709 ? meta_463_valid_1 : _GEN_978; // @[ICache.scala 132:{59,59}]
  wire  _GEN_980 = 9'h1d0 == _GEN_13709 ? meta_464_valid_1 : _GEN_979; // @[ICache.scala 132:{59,59}]
  wire  _GEN_981 = 9'h1d1 == _GEN_13709 ? meta_465_valid_1 : _GEN_980; // @[ICache.scala 132:{59,59}]
  wire  _GEN_982 = 9'h1d2 == _GEN_13709 ? meta_466_valid_1 : _GEN_981; // @[ICache.scala 132:{59,59}]
  wire  _GEN_983 = 9'h1d3 == _GEN_13709 ? meta_467_valid_1 : _GEN_982; // @[ICache.scala 132:{59,59}]
  wire  _GEN_984 = 9'h1d4 == _GEN_13709 ? meta_468_valid_1 : _GEN_983; // @[ICache.scala 132:{59,59}]
  wire  _GEN_985 = 9'h1d5 == _GEN_13709 ? meta_469_valid_1 : _GEN_984; // @[ICache.scala 132:{59,59}]
  wire  _GEN_986 = 9'h1d6 == _GEN_13709 ? meta_470_valid_1 : _GEN_985; // @[ICache.scala 132:{59,59}]
  wire  _GEN_987 = 9'h1d7 == _GEN_13709 ? meta_471_valid_1 : _GEN_986; // @[ICache.scala 132:{59,59}]
  wire  _GEN_988 = 9'h1d8 == _GEN_13709 ? meta_472_valid_1 : _GEN_987; // @[ICache.scala 132:{59,59}]
  wire  _GEN_989 = 9'h1d9 == _GEN_13709 ? meta_473_valid_1 : _GEN_988; // @[ICache.scala 132:{59,59}]
  wire  _GEN_990 = 9'h1da == _GEN_13709 ? meta_474_valid_1 : _GEN_989; // @[ICache.scala 132:{59,59}]
  wire  _GEN_991 = 9'h1db == _GEN_13709 ? meta_475_valid_1 : _GEN_990; // @[ICache.scala 132:{59,59}]
  wire  _GEN_992 = 9'h1dc == _GEN_13709 ? meta_476_valid_1 : _GEN_991; // @[ICache.scala 132:{59,59}]
  wire  _GEN_993 = 9'h1dd == _GEN_13709 ? meta_477_valid_1 : _GEN_992; // @[ICache.scala 132:{59,59}]
  wire  _GEN_994 = 9'h1de == _GEN_13709 ? meta_478_valid_1 : _GEN_993; // @[ICache.scala 132:{59,59}]
  wire  _GEN_995 = 9'h1df == _GEN_13709 ? meta_479_valid_1 : _GEN_994; // @[ICache.scala 132:{59,59}]
  wire  _GEN_996 = 9'h1e0 == _GEN_13709 ? meta_480_valid_1 : _GEN_995; // @[ICache.scala 132:{59,59}]
  wire  _GEN_997 = 9'h1e1 == _GEN_13709 ? meta_481_valid_1 : _GEN_996; // @[ICache.scala 132:{59,59}]
  wire  _GEN_998 = 9'h1e2 == _GEN_13709 ? meta_482_valid_1 : _GEN_997; // @[ICache.scala 132:{59,59}]
  wire  _GEN_999 = 9'h1e3 == _GEN_13709 ? meta_483_valid_1 : _GEN_998; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1000 = 9'h1e4 == _GEN_13709 ? meta_484_valid_1 : _GEN_999; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1001 = 9'h1e5 == _GEN_13709 ? meta_485_valid_1 : _GEN_1000; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1002 = 9'h1e6 == _GEN_13709 ? meta_486_valid_1 : _GEN_1001; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1003 = 9'h1e7 == _GEN_13709 ? meta_487_valid_1 : _GEN_1002; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1004 = 9'h1e8 == _GEN_13709 ? meta_488_valid_1 : _GEN_1003; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1005 = 9'h1e9 == _GEN_13709 ? meta_489_valid_1 : _GEN_1004; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1006 = 9'h1ea == _GEN_13709 ? meta_490_valid_1 : _GEN_1005; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1007 = 9'h1eb == _GEN_13709 ? meta_491_valid_1 : _GEN_1006; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1008 = 9'h1ec == _GEN_13709 ? meta_492_valid_1 : _GEN_1007; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1009 = 9'h1ed == _GEN_13709 ? meta_493_valid_1 : _GEN_1008; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1010 = 9'h1ee == _GEN_13709 ? meta_494_valid_1 : _GEN_1009; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1011 = 9'h1ef == _GEN_13709 ? meta_495_valid_1 : _GEN_1010; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1012 = 9'h1f0 == _GEN_13709 ? meta_496_valid_1 : _GEN_1011; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1013 = 9'h1f1 == _GEN_13709 ? meta_497_valid_1 : _GEN_1012; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1014 = 9'h1f2 == _GEN_13709 ? meta_498_valid_1 : _GEN_1013; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1015 = 9'h1f3 == _GEN_13709 ? meta_499_valid_1 : _GEN_1014; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1016 = 9'h1f4 == _GEN_13709 ? meta_500_valid_1 : _GEN_1015; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1017 = 9'h1f5 == _GEN_13709 ? meta_501_valid_1 : _GEN_1016; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1018 = 9'h1f6 == _GEN_13709 ? meta_502_valid_1 : _GEN_1017; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1019 = 9'h1f7 == _GEN_13709 ? meta_503_valid_1 : _GEN_1018; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1020 = 9'h1f8 == _GEN_13709 ? meta_504_valid_1 : _GEN_1019; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1021 = 9'h1f9 == _GEN_13709 ? meta_505_valid_1 : _GEN_1020; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1022 = 9'h1fa == _GEN_13709 ? meta_506_valid_1 : _GEN_1021; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1023 = 9'h1fb == _GEN_13709 ? meta_507_valid_1 : _GEN_1022; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1024 = 9'h1fc == _GEN_13709 ? meta_508_valid_1 : _GEN_1023; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1025 = 9'h1fd == _GEN_13709 ? meta_509_valid_1 : _GEN_1024; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1026 = 9'h1fe == _GEN_13709 ? meta_510_valid_1 : _GEN_1025; // @[ICache.scala 132:{59,59}]
  wire  _GEN_1027 = 9'h1ff == _GEN_13709 ? meta_511_valid_1 : _GEN_1026; // @[ICache.scala 132:{59,59}]
  wire  tag_compare_valid_1 = _GEN_13965 == inst_tag & _GEN_1027; // @[ICache.scala 132:59]
  wire  cache_hit = tag_compare_valid_0 | tag_compare_valid_1; // @[ICache.scala 71:55]
  wire  cache_hit_available = cache_hit & translation_ok & ~uncached; // @[ICache.scala 72:57]
  wire  cache_inst_ok_1 = cache_hit_available & ~io_cpu_addr_0[2]; // @[ICache.scala 76:43]
  wire [5:0] fence_index = io_cpu_fence_addr[11:6]; // @[ICache.scala 81:39]
  wire [63:0] cache_data_0 = bank_ram_io_way_0_r_data; // @[ICache.scala 122:19 63:28]
  wire [63:0] cache_data_1 = bank_ram_io_way_1_r_data; // @[ICache.scala 122:19 63:28]
  wire [63:0] _GEN_3 = tag_compare_valid_1 ? cache_data_1 : cache_data_0; // @[ICache.scala 86:{28,28}]
  wire [31:0] cache_inst_0 = io_cpu_addr_0[2] ? _GEN_3[63:32] : _GEN_3[31:0]; // @[ICache.scala 84:23]
  reg [31:0] saved_0_inst; // @[ICache.scala 91:22]
  reg  saved_0_valid; // @[ICache.scala 91:22]
  reg [31:0] saved_1_inst; // @[ICache.scala 91:22]
  reg  saved_1_valid; // @[ICache.scala 91:22]
  wire  _io_cpu_icache_stall_T = state == 3'h0; // @[ICache.scala 99:11]
  wire  _io_cpu_icache_stall_T_2 = ~cache_hit_available & io_cpu_req; // @[ICache.scala 100:27]
  wire  _io_cpu_inst_valid_0_T_1 = _io_cpu_icache_stall_T ? cache_hit_available : saved_0_valid; // @[ICache.scala 104:30]
  wire  _io_cpu_inst_valid_1_T_1 = _io_cpu_icache_stall_T ? cache_inst_ok_1 : saved_1_valid; // @[ICache.scala 105:30]
  reg [4:0] axi_cnt; // @[ICache.scala 109:24]
  wire [63:0] _bank_ram_io_way_0_w_data_T_1 = {io_axi_r_bits_data,32'h0}; // @[Cat.scala 33:92]
  wire [63:0] _bank_ram_io_way_0_w_data_T_2 = {32'h0,io_axi_r_bits_data}; // @[Cat.scala 33:92]
  wire  _T = ~io_cpu_icache_stall; // @[ICache.scala 135:28]
  wire  _T_2 = ~io_cpu_cpu_stall; // @[ICache.scala 135:52]
  wire  _GEN_1028 = io_cpu_fence_tlb & ~io_cpu_icache_stall & ~io_cpu_cpu_stall ? 1'h0 : tlb_valid; // @[ICache.scala 135:{71,83} 40:20]
  wire  _GEN_1029 = 6'h0 == fence_index ? 1'h0 : meta_0_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1030 = 6'h1 == fence_index ? 1'h0 : meta_1_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1031 = 6'h2 == fence_index ? 1'h0 : meta_2_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1032 = 6'h3 == fence_index ? 1'h0 : meta_3_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1033 = 6'h4 == fence_index ? 1'h0 : meta_4_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1034 = 6'h5 == fence_index ? 1'h0 : meta_5_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1035 = 6'h6 == fence_index ? 1'h0 : meta_6_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1036 = 6'h7 == fence_index ? 1'h0 : meta_7_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1037 = 6'h8 == fence_index ? 1'h0 : meta_8_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1038 = 6'h9 == fence_index ? 1'h0 : meta_9_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1039 = 6'ha == fence_index ? 1'h0 : meta_10_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1040 = 6'hb == fence_index ? 1'h0 : meta_11_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1041 = 6'hc == fence_index ? 1'h0 : meta_12_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1042 = 6'hd == fence_index ? 1'h0 : meta_13_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1043 = 6'he == fence_index ? 1'h0 : meta_14_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1044 = 6'hf == fence_index ? 1'h0 : meta_15_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1045 = 6'h10 == fence_index ? 1'h0 : meta_16_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1046 = 6'h11 == fence_index ? 1'h0 : meta_17_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1047 = 6'h12 == fence_index ? 1'h0 : meta_18_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1048 = 6'h13 == fence_index ? 1'h0 : meta_19_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1049 = 6'h14 == fence_index ? 1'h0 : meta_20_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1050 = 6'h15 == fence_index ? 1'h0 : meta_21_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1051 = 6'h16 == fence_index ? 1'h0 : meta_22_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1052 = 6'h17 == fence_index ? 1'h0 : meta_23_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1053 = 6'h18 == fence_index ? 1'h0 : meta_24_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1054 = 6'h19 == fence_index ? 1'h0 : meta_25_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1055 = 6'h1a == fence_index ? 1'h0 : meta_26_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1056 = 6'h1b == fence_index ? 1'h0 : meta_27_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1057 = 6'h1c == fence_index ? 1'h0 : meta_28_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1058 = 6'h1d == fence_index ? 1'h0 : meta_29_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1059 = 6'h1e == fence_index ? 1'h0 : meta_30_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1060 = 6'h1f == fence_index ? 1'h0 : meta_31_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1061 = 6'h20 == fence_index ? 1'h0 : meta_32_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1062 = 6'h21 == fence_index ? 1'h0 : meta_33_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1063 = 6'h22 == fence_index ? 1'h0 : meta_34_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1064 = 6'h23 == fence_index ? 1'h0 : meta_35_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1065 = 6'h24 == fence_index ? 1'h0 : meta_36_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1066 = 6'h25 == fence_index ? 1'h0 : meta_37_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1067 = 6'h26 == fence_index ? 1'h0 : meta_38_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1068 = 6'h27 == fence_index ? 1'h0 : meta_39_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1069 = 6'h28 == fence_index ? 1'h0 : meta_40_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1070 = 6'h29 == fence_index ? 1'h0 : meta_41_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1071 = 6'h2a == fence_index ? 1'h0 : meta_42_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1072 = 6'h2b == fence_index ? 1'h0 : meta_43_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1073 = 6'h2c == fence_index ? 1'h0 : meta_44_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1074 = 6'h2d == fence_index ? 1'h0 : meta_45_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1075 = 6'h2e == fence_index ? 1'h0 : meta_46_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1076 = 6'h2f == fence_index ? 1'h0 : meta_47_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1077 = 6'h30 == fence_index ? 1'h0 : meta_48_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1078 = 6'h31 == fence_index ? 1'h0 : meta_49_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1079 = 6'h32 == fence_index ? 1'h0 : meta_50_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1080 = 6'h33 == fence_index ? 1'h0 : meta_51_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1081 = 6'h34 == fence_index ? 1'h0 : meta_52_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1082 = 6'h35 == fence_index ? 1'h0 : meta_53_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1083 = 6'h36 == fence_index ? 1'h0 : meta_54_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1084 = 6'h37 == fence_index ? 1'h0 : meta_55_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1085 = 6'h38 == fence_index ? 1'h0 : meta_56_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1086 = 6'h39 == fence_index ? 1'h0 : meta_57_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1087 = 6'h3a == fence_index ? 1'h0 : meta_58_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1088 = 6'h3b == fence_index ? 1'h0 : meta_59_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1089 = 6'h3c == fence_index ? 1'h0 : meta_60_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1090 = 6'h3d == fence_index ? 1'h0 : meta_61_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1091 = 6'h3e == fence_index ? 1'h0 : meta_62_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1092 = 6'h3f == fence_index ? 1'h0 : meta_63_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire [6:0] _GEN_14414 = {{1'd0}, fence_index}; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1093 = 7'h40 == _GEN_14414 ? 1'h0 : meta_64_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1094 = 7'h41 == _GEN_14414 ? 1'h0 : meta_65_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1095 = 7'h42 == _GEN_14414 ? 1'h0 : meta_66_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1096 = 7'h43 == _GEN_14414 ? 1'h0 : meta_67_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1097 = 7'h44 == _GEN_14414 ? 1'h0 : meta_68_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1098 = 7'h45 == _GEN_14414 ? 1'h0 : meta_69_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1099 = 7'h46 == _GEN_14414 ? 1'h0 : meta_70_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1100 = 7'h47 == _GEN_14414 ? 1'h0 : meta_71_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1101 = 7'h48 == _GEN_14414 ? 1'h0 : meta_72_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1102 = 7'h49 == _GEN_14414 ? 1'h0 : meta_73_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1103 = 7'h4a == _GEN_14414 ? 1'h0 : meta_74_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1104 = 7'h4b == _GEN_14414 ? 1'h0 : meta_75_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1105 = 7'h4c == _GEN_14414 ? 1'h0 : meta_76_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1106 = 7'h4d == _GEN_14414 ? 1'h0 : meta_77_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1107 = 7'h4e == _GEN_14414 ? 1'h0 : meta_78_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1108 = 7'h4f == _GEN_14414 ? 1'h0 : meta_79_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1109 = 7'h50 == _GEN_14414 ? 1'h0 : meta_80_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1110 = 7'h51 == _GEN_14414 ? 1'h0 : meta_81_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1111 = 7'h52 == _GEN_14414 ? 1'h0 : meta_82_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1112 = 7'h53 == _GEN_14414 ? 1'h0 : meta_83_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1113 = 7'h54 == _GEN_14414 ? 1'h0 : meta_84_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1114 = 7'h55 == _GEN_14414 ? 1'h0 : meta_85_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1115 = 7'h56 == _GEN_14414 ? 1'h0 : meta_86_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1116 = 7'h57 == _GEN_14414 ? 1'h0 : meta_87_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1117 = 7'h58 == _GEN_14414 ? 1'h0 : meta_88_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1118 = 7'h59 == _GEN_14414 ? 1'h0 : meta_89_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1119 = 7'h5a == _GEN_14414 ? 1'h0 : meta_90_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1120 = 7'h5b == _GEN_14414 ? 1'h0 : meta_91_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1121 = 7'h5c == _GEN_14414 ? 1'h0 : meta_92_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1122 = 7'h5d == _GEN_14414 ? 1'h0 : meta_93_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1123 = 7'h5e == _GEN_14414 ? 1'h0 : meta_94_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1124 = 7'h5f == _GEN_14414 ? 1'h0 : meta_95_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1125 = 7'h60 == _GEN_14414 ? 1'h0 : meta_96_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1126 = 7'h61 == _GEN_14414 ? 1'h0 : meta_97_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1127 = 7'h62 == _GEN_14414 ? 1'h0 : meta_98_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1128 = 7'h63 == _GEN_14414 ? 1'h0 : meta_99_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1129 = 7'h64 == _GEN_14414 ? 1'h0 : meta_100_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1130 = 7'h65 == _GEN_14414 ? 1'h0 : meta_101_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1131 = 7'h66 == _GEN_14414 ? 1'h0 : meta_102_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1132 = 7'h67 == _GEN_14414 ? 1'h0 : meta_103_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1133 = 7'h68 == _GEN_14414 ? 1'h0 : meta_104_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1134 = 7'h69 == _GEN_14414 ? 1'h0 : meta_105_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1135 = 7'h6a == _GEN_14414 ? 1'h0 : meta_106_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1136 = 7'h6b == _GEN_14414 ? 1'h0 : meta_107_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1137 = 7'h6c == _GEN_14414 ? 1'h0 : meta_108_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1138 = 7'h6d == _GEN_14414 ? 1'h0 : meta_109_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1139 = 7'h6e == _GEN_14414 ? 1'h0 : meta_110_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1140 = 7'h6f == _GEN_14414 ? 1'h0 : meta_111_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1141 = 7'h70 == _GEN_14414 ? 1'h0 : meta_112_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1142 = 7'h71 == _GEN_14414 ? 1'h0 : meta_113_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1143 = 7'h72 == _GEN_14414 ? 1'h0 : meta_114_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1144 = 7'h73 == _GEN_14414 ? 1'h0 : meta_115_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1145 = 7'h74 == _GEN_14414 ? 1'h0 : meta_116_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1146 = 7'h75 == _GEN_14414 ? 1'h0 : meta_117_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1147 = 7'h76 == _GEN_14414 ? 1'h0 : meta_118_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1148 = 7'h77 == _GEN_14414 ? 1'h0 : meta_119_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1149 = 7'h78 == _GEN_14414 ? 1'h0 : meta_120_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1150 = 7'h79 == _GEN_14414 ? 1'h0 : meta_121_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1151 = 7'h7a == _GEN_14414 ? 1'h0 : meta_122_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1152 = 7'h7b == _GEN_14414 ? 1'h0 : meta_123_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1153 = 7'h7c == _GEN_14414 ? 1'h0 : meta_124_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1154 = 7'h7d == _GEN_14414 ? 1'h0 : meta_125_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1155 = 7'h7e == _GEN_14414 ? 1'h0 : meta_126_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1156 = 7'h7f == _GEN_14414 ? 1'h0 : meta_127_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire [7:0] _GEN_14478 = {{2'd0}, fence_index}; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1157 = 8'h80 == _GEN_14478 ? 1'h0 : meta_128_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1158 = 8'h81 == _GEN_14478 ? 1'h0 : meta_129_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1159 = 8'h82 == _GEN_14478 ? 1'h0 : meta_130_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1160 = 8'h83 == _GEN_14478 ? 1'h0 : meta_131_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1161 = 8'h84 == _GEN_14478 ? 1'h0 : meta_132_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1162 = 8'h85 == _GEN_14478 ? 1'h0 : meta_133_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1163 = 8'h86 == _GEN_14478 ? 1'h0 : meta_134_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1164 = 8'h87 == _GEN_14478 ? 1'h0 : meta_135_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1165 = 8'h88 == _GEN_14478 ? 1'h0 : meta_136_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1166 = 8'h89 == _GEN_14478 ? 1'h0 : meta_137_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1167 = 8'h8a == _GEN_14478 ? 1'h0 : meta_138_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1168 = 8'h8b == _GEN_14478 ? 1'h0 : meta_139_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1169 = 8'h8c == _GEN_14478 ? 1'h0 : meta_140_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1170 = 8'h8d == _GEN_14478 ? 1'h0 : meta_141_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1171 = 8'h8e == _GEN_14478 ? 1'h0 : meta_142_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1172 = 8'h8f == _GEN_14478 ? 1'h0 : meta_143_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1173 = 8'h90 == _GEN_14478 ? 1'h0 : meta_144_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1174 = 8'h91 == _GEN_14478 ? 1'h0 : meta_145_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1175 = 8'h92 == _GEN_14478 ? 1'h0 : meta_146_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1176 = 8'h93 == _GEN_14478 ? 1'h0 : meta_147_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1177 = 8'h94 == _GEN_14478 ? 1'h0 : meta_148_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1178 = 8'h95 == _GEN_14478 ? 1'h0 : meta_149_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1179 = 8'h96 == _GEN_14478 ? 1'h0 : meta_150_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1180 = 8'h97 == _GEN_14478 ? 1'h0 : meta_151_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1181 = 8'h98 == _GEN_14478 ? 1'h0 : meta_152_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1182 = 8'h99 == _GEN_14478 ? 1'h0 : meta_153_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1183 = 8'h9a == _GEN_14478 ? 1'h0 : meta_154_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1184 = 8'h9b == _GEN_14478 ? 1'h0 : meta_155_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1185 = 8'h9c == _GEN_14478 ? 1'h0 : meta_156_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1186 = 8'h9d == _GEN_14478 ? 1'h0 : meta_157_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1187 = 8'h9e == _GEN_14478 ? 1'h0 : meta_158_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1188 = 8'h9f == _GEN_14478 ? 1'h0 : meta_159_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1189 = 8'ha0 == _GEN_14478 ? 1'h0 : meta_160_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1190 = 8'ha1 == _GEN_14478 ? 1'h0 : meta_161_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1191 = 8'ha2 == _GEN_14478 ? 1'h0 : meta_162_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1192 = 8'ha3 == _GEN_14478 ? 1'h0 : meta_163_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1193 = 8'ha4 == _GEN_14478 ? 1'h0 : meta_164_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1194 = 8'ha5 == _GEN_14478 ? 1'h0 : meta_165_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1195 = 8'ha6 == _GEN_14478 ? 1'h0 : meta_166_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1196 = 8'ha7 == _GEN_14478 ? 1'h0 : meta_167_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1197 = 8'ha8 == _GEN_14478 ? 1'h0 : meta_168_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1198 = 8'ha9 == _GEN_14478 ? 1'h0 : meta_169_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1199 = 8'haa == _GEN_14478 ? 1'h0 : meta_170_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1200 = 8'hab == _GEN_14478 ? 1'h0 : meta_171_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1201 = 8'hac == _GEN_14478 ? 1'h0 : meta_172_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1202 = 8'had == _GEN_14478 ? 1'h0 : meta_173_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1203 = 8'hae == _GEN_14478 ? 1'h0 : meta_174_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1204 = 8'haf == _GEN_14478 ? 1'h0 : meta_175_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1205 = 8'hb0 == _GEN_14478 ? 1'h0 : meta_176_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1206 = 8'hb1 == _GEN_14478 ? 1'h0 : meta_177_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1207 = 8'hb2 == _GEN_14478 ? 1'h0 : meta_178_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1208 = 8'hb3 == _GEN_14478 ? 1'h0 : meta_179_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1209 = 8'hb4 == _GEN_14478 ? 1'h0 : meta_180_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1210 = 8'hb5 == _GEN_14478 ? 1'h0 : meta_181_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1211 = 8'hb6 == _GEN_14478 ? 1'h0 : meta_182_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1212 = 8'hb7 == _GEN_14478 ? 1'h0 : meta_183_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1213 = 8'hb8 == _GEN_14478 ? 1'h0 : meta_184_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1214 = 8'hb9 == _GEN_14478 ? 1'h0 : meta_185_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1215 = 8'hba == _GEN_14478 ? 1'h0 : meta_186_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1216 = 8'hbb == _GEN_14478 ? 1'h0 : meta_187_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1217 = 8'hbc == _GEN_14478 ? 1'h0 : meta_188_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1218 = 8'hbd == _GEN_14478 ? 1'h0 : meta_189_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1219 = 8'hbe == _GEN_14478 ? 1'h0 : meta_190_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1220 = 8'hbf == _GEN_14478 ? 1'h0 : meta_191_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1221 = 8'hc0 == _GEN_14478 ? 1'h0 : meta_192_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1222 = 8'hc1 == _GEN_14478 ? 1'h0 : meta_193_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1223 = 8'hc2 == _GEN_14478 ? 1'h0 : meta_194_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1224 = 8'hc3 == _GEN_14478 ? 1'h0 : meta_195_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1225 = 8'hc4 == _GEN_14478 ? 1'h0 : meta_196_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1226 = 8'hc5 == _GEN_14478 ? 1'h0 : meta_197_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1227 = 8'hc6 == _GEN_14478 ? 1'h0 : meta_198_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1228 = 8'hc7 == _GEN_14478 ? 1'h0 : meta_199_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1229 = 8'hc8 == _GEN_14478 ? 1'h0 : meta_200_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1230 = 8'hc9 == _GEN_14478 ? 1'h0 : meta_201_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1231 = 8'hca == _GEN_14478 ? 1'h0 : meta_202_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1232 = 8'hcb == _GEN_14478 ? 1'h0 : meta_203_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1233 = 8'hcc == _GEN_14478 ? 1'h0 : meta_204_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1234 = 8'hcd == _GEN_14478 ? 1'h0 : meta_205_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1235 = 8'hce == _GEN_14478 ? 1'h0 : meta_206_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1236 = 8'hcf == _GEN_14478 ? 1'h0 : meta_207_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1237 = 8'hd0 == _GEN_14478 ? 1'h0 : meta_208_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1238 = 8'hd1 == _GEN_14478 ? 1'h0 : meta_209_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1239 = 8'hd2 == _GEN_14478 ? 1'h0 : meta_210_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1240 = 8'hd3 == _GEN_14478 ? 1'h0 : meta_211_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1241 = 8'hd4 == _GEN_14478 ? 1'h0 : meta_212_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1242 = 8'hd5 == _GEN_14478 ? 1'h0 : meta_213_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1243 = 8'hd6 == _GEN_14478 ? 1'h0 : meta_214_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1244 = 8'hd7 == _GEN_14478 ? 1'h0 : meta_215_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1245 = 8'hd8 == _GEN_14478 ? 1'h0 : meta_216_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1246 = 8'hd9 == _GEN_14478 ? 1'h0 : meta_217_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1247 = 8'hda == _GEN_14478 ? 1'h0 : meta_218_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1248 = 8'hdb == _GEN_14478 ? 1'h0 : meta_219_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1249 = 8'hdc == _GEN_14478 ? 1'h0 : meta_220_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1250 = 8'hdd == _GEN_14478 ? 1'h0 : meta_221_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1251 = 8'hde == _GEN_14478 ? 1'h0 : meta_222_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1252 = 8'hdf == _GEN_14478 ? 1'h0 : meta_223_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1253 = 8'he0 == _GEN_14478 ? 1'h0 : meta_224_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1254 = 8'he1 == _GEN_14478 ? 1'h0 : meta_225_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1255 = 8'he2 == _GEN_14478 ? 1'h0 : meta_226_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1256 = 8'he3 == _GEN_14478 ? 1'h0 : meta_227_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1257 = 8'he4 == _GEN_14478 ? 1'h0 : meta_228_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1258 = 8'he5 == _GEN_14478 ? 1'h0 : meta_229_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1259 = 8'he6 == _GEN_14478 ? 1'h0 : meta_230_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1260 = 8'he7 == _GEN_14478 ? 1'h0 : meta_231_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1261 = 8'he8 == _GEN_14478 ? 1'h0 : meta_232_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1262 = 8'he9 == _GEN_14478 ? 1'h0 : meta_233_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1263 = 8'hea == _GEN_14478 ? 1'h0 : meta_234_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1264 = 8'heb == _GEN_14478 ? 1'h0 : meta_235_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1265 = 8'hec == _GEN_14478 ? 1'h0 : meta_236_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1266 = 8'hed == _GEN_14478 ? 1'h0 : meta_237_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1267 = 8'hee == _GEN_14478 ? 1'h0 : meta_238_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1268 = 8'hef == _GEN_14478 ? 1'h0 : meta_239_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1269 = 8'hf0 == _GEN_14478 ? 1'h0 : meta_240_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1270 = 8'hf1 == _GEN_14478 ? 1'h0 : meta_241_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1271 = 8'hf2 == _GEN_14478 ? 1'h0 : meta_242_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1272 = 8'hf3 == _GEN_14478 ? 1'h0 : meta_243_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1273 = 8'hf4 == _GEN_14478 ? 1'h0 : meta_244_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1274 = 8'hf5 == _GEN_14478 ? 1'h0 : meta_245_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1275 = 8'hf6 == _GEN_14478 ? 1'h0 : meta_246_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1276 = 8'hf7 == _GEN_14478 ? 1'h0 : meta_247_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1277 = 8'hf8 == _GEN_14478 ? 1'h0 : meta_248_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1278 = 8'hf9 == _GEN_14478 ? 1'h0 : meta_249_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1279 = 8'hfa == _GEN_14478 ? 1'h0 : meta_250_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1280 = 8'hfb == _GEN_14478 ? 1'h0 : meta_251_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1281 = 8'hfc == _GEN_14478 ? 1'h0 : meta_252_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1282 = 8'hfd == _GEN_14478 ? 1'h0 : meta_253_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1283 = 8'hfe == _GEN_14478 ? 1'h0 : meta_254_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1284 = 8'hff == _GEN_14478 ? 1'h0 : meta_255_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire [8:0] _GEN_14606 = {{3'd0}, fence_index}; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1285 = 9'h100 == _GEN_14606 ? 1'h0 : meta_256_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1286 = 9'h101 == _GEN_14606 ? 1'h0 : meta_257_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1287 = 9'h102 == _GEN_14606 ? 1'h0 : meta_258_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1288 = 9'h103 == _GEN_14606 ? 1'h0 : meta_259_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1289 = 9'h104 == _GEN_14606 ? 1'h0 : meta_260_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1290 = 9'h105 == _GEN_14606 ? 1'h0 : meta_261_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1291 = 9'h106 == _GEN_14606 ? 1'h0 : meta_262_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1292 = 9'h107 == _GEN_14606 ? 1'h0 : meta_263_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1293 = 9'h108 == _GEN_14606 ? 1'h0 : meta_264_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1294 = 9'h109 == _GEN_14606 ? 1'h0 : meta_265_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1295 = 9'h10a == _GEN_14606 ? 1'h0 : meta_266_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1296 = 9'h10b == _GEN_14606 ? 1'h0 : meta_267_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1297 = 9'h10c == _GEN_14606 ? 1'h0 : meta_268_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1298 = 9'h10d == _GEN_14606 ? 1'h0 : meta_269_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1299 = 9'h10e == _GEN_14606 ? 1'h0 : meta_270_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1300 = 9'h10f == _GEN_14606 ? 1'h0 : meta_271_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1301 = 9'h110 == _GEN_14606 ? 1'h0 : meta_272_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1302 = 9'h111 == _GEN_14606 ? 1'h0 : meta_273_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1303 = 9'h112 == _GEN_14606 ? 1'h0 : meta_274_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1304 = 9'h113 == _GEN_14606 ? 1'h0 : meta_275_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1305 = 9'h114 == _GEN_14606 ? 1'h0 : meta_276_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1306 = 9'h115 == _GEN_14606 ? 1'h0 : meta_277_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1307 = 9'h116 == _GEN_14606 ? 1'h0 : meta_278_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1308 = 9'h117 == _GEN_14606 ? 1'h0 : meta_279_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1309 = 9'h118 == _GEN_14606 ? 1'h0 : meta_280_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1310 = 9'h119 == _GEN_14606 ? 1'h0 : meta_281_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1311 = 9'h11a == _GEN_14606 ? 1'h0 : meta_282_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1312 = 9'h11b == _GEN_14606 ? 1'h0 : meta_283_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1313 = 9'h11c == _GEN_14606 ? 1'h0 : meta_284_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1314 = 9'h11d == _GEN_14606 ? 1'h0 : meta_285_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1315 = 9'h11e == _GEN_14606 ? 1'h0 : meta_286_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1316 = 9'h11f == _GEN_14606 ? 1'h0 : meta_287_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1317 = 9'h120 == _GEN_14606 ? 1'h0 : meta_288_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1318 = 9'h121 == _GEN_14606 ? 1'h0 : meta_289_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1319 = 9'h122 == _GEN_14606 ? 1'h0 : meta_290_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1320 = 9'h123 == _GEN_14606 ? 1'h0 : meta_291_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1321 = 9'h124 == _GEN_14606 ? 1'h0 : meta_292_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1322 = 9'h125 == _GEN_14606 ? 1'h0 : meta_293_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1323 = 9'h126 == _GEN_14606 ? 1'h0 : meta_294_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1324 = 9'h127 == _GEN_14606 ? 1'h0 : meta_295_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1325 = 9'h128 == _GEN_14606 ? 1'h0 : meta_296_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1326 = 9'h129 == _GEN_14606 ? 1'h0 : meta_297_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1327 = 9'h12a == _GEN_14606 ? 1'h0 : meta_298_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1328 = 9'h12b == _GEN_14606 ? 1'h0 : meta_299_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1329 = 9'h12c == _GEN_14606 ? 1'h0 : meta_300_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1330 = 9'h12d == _GEN_14606 ? 1'h0 : meta_301_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1331 = 9'h12e == _GEN_14606 ? 1'h0 : meta_302_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1332 = 9'h12f == _GEN_14606 ? 1'h0 : meta_303_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1333 = 9'h130 == _GEN_14606 ? 1'h0 : meta_304_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1334 = 9'h131 == _GEN_14606 ? 1'h0 : meta_305_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1335 = 9'h132 == _GEN_14606 ? 1'h0 : meta_306_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1336 = 9'h133 == _GEN_14606 ? 1'h0 : meta_307_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1337 = 9'h134 == _GEN_14606 ? 1'h0 : meta_308_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1338 = 9'h135 == _GEN_14606 ? 1'h0 : meta_309_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1339 = 9'h136 == _GEN_14606 ? 1'h0 : meta_310_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1340 = 9'h137 == _GEN_14606 ? 1'h0 : meta_311_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1341 = 9'h138 == _GEN_14606 ? 1'h0 : meta_312_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1342 = 9'h139 == _GEN_14606 ? 1'h0 : meta_313_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1343 = 9'h13a == _GEN_14606 ? 1'h0 : meta_314_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1344 = 9'h13b == _GEN_14606 ? 1'h0 : meta_315_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1345 = 9'h13c == _GEN_14606 ? 1'h0 : meta_316_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1346 = 9'h13d == _GEN_14606 ? 1'h0 : meta_317_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1347 = 9'h13e == _GEN_14606 ? 1'h0 : meta_318_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1348 = 9'h13f == _GEN_14606 ? 1'h0 : meta_319_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1349 = 9'h140 == _GEN_14606 ? 1'h0 : meta_320_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1350 = 9'h141 == _GEN_14606 ? 1'h0 : meta_321_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1351 = 9'h142 == _GEN_14606 ? 1'h0 : meta_322_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1352 = 9'h143 == _GEN_14606 ? 1'h0 : meta_323_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1353 = 9'h144 == _GEN_14606 ? 1'h0 : meta_324_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1354 = 9'h145 == _GEN_14606 ? 1'h0 : meta_325_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1355 = 9'h146 == _GEN_14606 ? 1'h0 : meta_326_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1356 = 9'h147 == _GEN_14606 ? 1'h0 : meta_327_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1357 = 9'h148 == _GEN_14606 ? 1'h0 : meta_328_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1358 = 9'h149 == _GEN_14606 ? 1'h0 : meta_329_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1359 = 9'h14a == _GEN_14606 ? 1'h0 : meta_330_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1360 = 9'h14b == _GEN_14606 ? 1'h0 : meta_331_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1361 = 9'h14c == _GEN_14606 ? 1'h0 : meta_332_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1362 = 9'h14d == _GEN_14606 ? 1'h0 : meta_333_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1363 = 9'h14e == _GEN_14606 ? 1'h0 : meta_334_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1364 = 9'h14f == _GEN_14606 ? 1'h0 : meta_335_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1365 = 9'h150 == _GEN_14606 ? 1'h0 : meta_336_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1366 = 9'h151 == _GEN_14606 ? 1'h0 : meta_337_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1367 = 9'h152 == _GEN_14606 ? 1'h0 : meta_338_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1368 = 9'h153 == _GEN_14606 ? 1'h0 : meta_339_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1369 = 9'h154 == _GEN_14606 ? 1'h0 : meta_340_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1370 = 9'h155 == _GEN_14606 ? 1'h0 : meta_341_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1371 = 9'h156 == _GEN_14606 ? 1'h0 : meta_342_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1372 = 9'h157 == _GEN_14606 ? 1'h0 : meta_343_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1373 = 9'h158 == _GEN_14606 ? 1'h0 : meta_344_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1374 = 9'h159 == _GEN_14606 ? 1'h0 : meta_345_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1375 = 9'h15a == _GEN_14606 ? 1'h0 : meta_346_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1376 = 9'h15b == _GEN_14606 ? 1'h0 : meta_347_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1377 = 9'h15c == _GEN_14606 ? 1'h0 : meta_348_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1378 = 9'h15d == _GEN_14606 ? 1'h0 : meta_349_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1379 = 9'h15e == _GEN_14606 ? 1'h0 : meta_350_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1380 = 9'h15f == _GEN_14606 ? 1'h0 : meta_351_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1381 = 9'h160 == _GEN_14606 ? 1'h0 : meta_352_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1382 = 9'h161 == _GEN_14606 ? 1'h0 : meta_353_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1383 = 9'h162 == _GEN_14606 ? 1'h0 : meta_354_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1384 = 9'h163 == _GEN_14606 ? 1'h0 : meta_355_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1385 = 9'h164 == _GEN_14606 ? 1'h0 : meta_356_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1386 = 9'h165 == _GEN_14606 ? 1'h0 : meta_357_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1387 = 9'h166 == _GEN_14606 ? 1'h0 : meta_358_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1388 = 9'h167 == _GEN_14606 ? 1'h0 : meta_359_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1389 = 9'h168 == _GEN_14606 ? 1'h0 : meta_360_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1390 = 9'h169 == _GEN_14606 ? 1'h0 : meta_361_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1391 = 9'h16a == _GEN_14606 ? 1'h0 : meta_362_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1392 = 9'h16b == _GEN_14606 ? 1'h0 : meta_363_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1393 = 9'h16c == _GEN_14606 ? 1'h0 : meta_364_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1394 = 9'h16d == _GEN_14606 ? 1'h0 : meta_365_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1395 = 9'h16e == _GEN_14606 ? 1'h0 : meta_366_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1396 = 9'h16f == _GEN_14606 ? 1'h0 : meta_367_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1397 = 9'h170 == _GEN_14606 ? 1'h0 : meta_368_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1398 = 9'h171 == _GEN_14606 ? 1'h0 : meta_369_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1399 = 9'h172 == _GEN_14606 ? 1'h0 : meta_370_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1400 = 9'h173 == _GEN_14606 ? 1'h0 : meta_371_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1401 = 9'h174 == _GEN_14606 ? 1'h0 : meta_372_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1402 = 9'h175 == _GEN_14606 ? 1'h0 : meta_373_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1403 = 9'h176 == _GEN_14606 ? 1'h0 : meta_374_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1404 = 9'h177 == _GEN_14606 ? 1'h0 : meta_375_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1405 = 9'h178 == _GEN_14606 ? 1'h0 : meta_376_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1406 = 9'h179 == _GEN_14606 ? 1'h0 : meta_377_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1407 = 9'h17a == _GEN_14606 ? 1'h0 : meta_378_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1408 = 9'h17b == _GEN_14606 ? 1'h0 : meta_379_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1409 = 9'h17c == _GEN_14606 ? 1'h0 : meta_380_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1410 = 9'h17d == _GEN_14606 ? 1'h0 : meta_381_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1411 = 9'h17e == _GEN_14606 ? 1'h0 : meta_382_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1412 = 9'h17f == _GEN_14606 ? 1'h0 : meta_383_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1413 = 9'h180 == _GEN_14606 ? 1'h0 : meta_384_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1414 = 9'h181 == _GEN_14606 ? 1'h0 : meta_385_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1415 = 9'h182 == _GEN_14606 ? 1'h0 : meta_386_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1416 = 9'h183 == _GEN_14606 ? 1'h0 : meta_387_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1417 = 9'h184 == _GEN_14606 ? 1'h0 : meta_388_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1418 = 9'h185 == _GEN_14606 ? 1'h0 : meta_389_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1419 = 9'h186 == _GEN_14606 ? 1'h0 : meta_390_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1420 = 9'h187 == _GEN_14606 ? 1'h0 : meta_391_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1421 = 9'h188 == _GEN_14606 ? 1'h0 : meta_392_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1422 = 9'h189 == _GEN_14606 ? 1'h0 : meta_393_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1423 = 9'h18a == _GEN_14606 ? 1'h0 : meta_394_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1424 = 9'h18b == _GEN_14606 ? 1'h0 : meta_395_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1425 = 9'h18c == _GEN_14606 ? 1'h0 : meta_396_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1426 = 9'h18d == _GEN_14606 ? 1'h0 : meta_397_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1427 = 9'h18e == _GEN_14606 ? 1'h0 : meta_398_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1428 = 9'h18f == _GEN_14606 ? 1'h0 : meta_399_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1429 = 9'h190 == _GEN_14606 ? 1'h0 : meta_400_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1430 = 9'h191 == _GEN_14606 ? 1'h0 : meta_401_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1431 = 9'h192 == _GEN_14606 ? 1'h0 : meta_402_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1432 = 9'h193 == _GEN_14606 ? 1'h0 : meta_403_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1433 = 9'h194 == _GEN_14606 ? 1'h0 : meta_404_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1434 = 9'h195 == _GEN_14606 ? 1'h0 : meta_405_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1435 = 9'h196 == _GEN_14606 ? 1'h0 : meta_406_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1436 = 9'h197 == _GEN_14606 ? 1'h0 : meta_407_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1437 = 9'h198 == _GEN_14606 ? 1'h0 : meta_408_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1438 = 9'h199 == _GEN_14606 ? 1'h0 : meta_409_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1439 = 9'h19a == _GEN_14606 ? 1'h0 : meta_410_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1440 = 9'h19b == _GEN_14606 ? 1'h0 : meta_411_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1441 = 9'h19c == _GEN_14606 ? 1'h0 : meta_412_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1442 = 9'h19d == _GEN_14606 ? 1'h0 : meta_413_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1443 = 9'h19e == _GEN_14606 ? 1'h0 : meta_414_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1444 = 9'h19f == _GEN_14606 ? 1'h0 : meta_415_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1445 = 9'h1a0 == _GEN_14606 ? 1'h0 : meta_416_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1446 = 9'h1a1 == _GEN_14606 ? 1'h0 : meta_417_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1447 = 9'h1a2 == _GEN_14606 ? 1'h0 : meta_418_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1448 = 9'h1a3 == _GEN_14606 ? 1'h0 : meta_419_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1449 = 9'h1a4 == _GEN_14606 ? 1'h0 : meta_420_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1450 = 9'h1a5 == _GEN_14606 ? 1'h0 : meta_421_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1451 = 9'h1a6 == _GEN_14606 ? 1'h0 : meta_422_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1452 = 9'h1a7 == _GEN_14606 ? 1'h0 : meta_423_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1453 = 9'h1a8 == _GEN_14606 ? 1'h0 : meta_424_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1454 = 9'h1a9 == _GEN_14606 ? 1'h0 : meta_425_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1455 = 9'h1aa == _GEN_14606 ? 1'h0 : meta_426_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1456 = 9'h1ab == _GEN_14606 ? 1'h0 : meta_427_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1457 = 9'h1ac == _GEN_14606 ? 1'h0 : meta_428_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1458 = 9'h1ad == _GEN_14606 ? 1'h0 : meta_429_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1459 = 9'h1ae == _GEN_14606 ? 1'h0 : meta_430_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1460 = 9'h1af == _GEN_14606 ? 1'h0 : meta_431_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1461 = 9'h1b0 == _GEN_14606 ? 1'h0 : meta_432_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1462 = 9'h1b1 == _GEN_14606 ? 1'h0 : meta_433_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1463 = 9'h1b2 == _GEN_14606 ? 1'h0 : meta_434_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1464 = 9'h1b3 == _GEN_14606 ? 1'h0 : meta_435_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1465 = 9'h1b4 == _GEN_14606 ? 1'h0 : meta_436_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1466 = 9'h1b5 == _GEN_14606 ? 1'h0 : meta_437_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1467 = 9'h1b6 == _GEN_14606 ? 1'h0 : meta_438_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1468 = 9'h1b7 == _GEN_14606 ? 1'h0 : meta_439_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1469 = 9'h1b8 == _GEN_14606 ? 1'h0 : meta_440_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1470 = 9'h1b9 == _GEN_14606 ? 1'h0 : meta_441_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1471 = 9'h1ba == _GEN_14606 ? 1'h0 : meta_442_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1472 = 9'h1bb == _GEN_14606 ? 1'h0 : meta_443_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1473 = 9'h1bc == _GEN_14606 ? 1'h0 : meta_444_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1474 = 9'h1bd == _GEN_14606 ? 1'h0 : meta_445_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1475 = 9'h1be == _GEN_14606 ? 1'h0 : meta_446_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1476 = 9'h1bf == _GEN_14606 ? 1'h0 : meta_447_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1477 = 9'h1c0 == _GEN_14606 ? 1'h0 : meta_448_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1478 = 9'h1c1 == _GEN_14606 ? 1'h0 : meta_449_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1479 = 9'h1c2 == _GEN_14606 ? 1'h0 : meta_450_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1480 = 9'h1c3 == _GEN_14606 ? 1'h0 : meta_451_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1481 = 9'h1c4 == _GEN_14606 ? 1'h0 : meta_452_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1482 = 9'h1c5 == _GEN_14606 ? 1'h0 : meta_453_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1483 = 9'h1c6 == _GEN_14606 ? 1'h0 : meta_454_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1484 = 9'h1c7 == _GEN_14606 ? 1'h0 : meta_455_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1485 = 9'h1c8 == _GEN_14606 ? 1'h0 : meta_456_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1486 = 9'h1c9 == _GEN_14606 ? 1'h0 : meta_457_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1487 = 9'h1ca == _GEN_14606 ? 1'h0 : meta_458_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1488 = 9'h1cb == _GEN_14606 ? 1'h0 : meta_459_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1489 = 9'h1cc == _GEN_14606 ? 1'h0 : meta_460_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1490 = 9'h1cd == _GEN_14606 ? 1'h0 : meta_461_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1491 = 9'h1ce == _GEN_14606 ? 1'h0 : meta_462_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1492 = 9'h1cf == _GEN_14606 ? 1'h0 : meta_463_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1493 = 9'h1d0 == _GEN_14606 ? 1'h0 : meta_464_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1494 = 9'h1d1 == _GEN_14606 ? 1'h0 : meta_465_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1495 = 9'h1d2 == _GEN_14606 ? 1'h0 : meta_466_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1496 = 9'h1d3 == _GEN_14606 ? 1'h0 : meta_467_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1497 = 9'h1d4 == _GEN_14606 ? 1'h0 : meta_468_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1498 = 9'h1d5 == _GEN_14606 ? 1'h0 : meta_469_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1499 = 9'h1d6 == _GEN_14606 ? 1'h0 : meta_470_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1500 = 9'h1d7 == _GEN_14606 ? 1'h0 : meta_471_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1501 = 9'h1d8 == _GEN_14606 ? 1'h0 : meta_472_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1502 = 9'h1d9 == _GEN_14606 ? 1'h0 : meta_473_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1503 = 9'h1da == _GEN_14606 ? 1'h0 : meta_474_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1504 = 9'h1db == _GEN_14606 ? 1'h0 : meta_475_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1505 = 9'h1dc == _GEN_14606 ? 1'h0 : meta_476_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1506 = 9'h1dd == _GEN_14606 ? 1'h0 : meta_477_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1507 = 9'h1de == _GEN_14606 ? 1'h0 : meta_478_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1508 = 9'h1df == _GEN_14606 ? 1'h0 : meta_479_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1509 = 9'h1e0 == _GEN_14606 ? 1'h0 : meta_480_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1510 = 9'h1e1 == _GEN_14606 ? 1'h0 : meta_481_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1511 = 9'h1e2 == _GEN_14606 ? 1'h0 : meta_482_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1512 = 9'h1e3 == _GEN_14606 ? 1'h0 : meta_483_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1513 = 9'h1e4 == _GEN_14606 ? 1'h0 : meta_484_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1514 = 9'h1e5 == _GEN_14606 ? 1'h0 : meta_485_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1515 = 9'h1e6 == _GEN_14606 ? 1'h0 : meta_486_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1516 = 9'h1e7 == _GEN_14606 ? 1'h0 : meta_487_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1517 = 9'h1e8 == _GEN_14606 ? 1'h0 : meta_488_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1518 = 9'h1e9 == _GEN_14606 ? 1'h0 : meta_489_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1519 = 9'h1ea == _GEN_14606 ? 1'h0 : meta_490_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1520 = 9'h1eb == _GEN_14606 ? 1'h0 : meta_491_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1521 = 9'h1ec == _GEN_14606 ? 1'h0 : meta_492_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1522 = 9'h1ed == _GEN_14606 ? 1'h0 : meta_493_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1523 = 9'h1ee == _GEN_14606 ? 1'h0 : meta_494_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1524 = 9'h1ef == _GEN_14606 ? 1'h0 : meta_495_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1525 = 9'h1f0 == _GEN_14606 ? 1'h0 : meta_496_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1526 = 9'h1f1 == _GEN_14606 ? 1'h0 : meta_497_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1527 = 9'h1f2 == _GEN_14606 ? 1'h0 : meta_498_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1528 = 9'h1f3 == _GEN_14606 ? 1'h0 : meta_499_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1529 = 9'h1f4 == _GEN_14606 ? 1'h0 : meta_500_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1530 = 9'h1f5 == _GEN_14606 ? 1'h0 : meta_501_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1531 = 9'h1f6 == _GEN_14606 ? 1'h0 : meta_502_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1532 = 9'h1f7 == _GEN_14606 ? 1'h0 : meta_503_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1533 = 9'h1f8 == _GEN_14606 ? 1'h0 : meta_504_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1534 = 9'h1f9 == _GEN_14606 ? 1'h0 : meta_505_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1535 = 9'h1fa == _GEN_14606 ? 1'h0 : meta_506_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1536 = 9'h1fb == _GEN_14606 ? 1'h0 : meta_507_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1537 = 9'h1fc == _GEN_14606 ? 1'h0 : meta_508_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1538 = 9'h1fd == _GEN_14606 ? 1'h0 : meta_509_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1539 = 9'h1fe == _GEN_14606 ? 1'h0 : meta_510_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1540 = 9'h1ff == _GEN_14606 ? 1'h0 : meta_511_valid_0; // @[ICache.scala 137:{32,32} 34:21]
  wire  _GEN_1541 = 6'h0 == fence_index ? 1'h0 : meta_0_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1542 = 6'h1 == fence_index ? 1'h0 : meta_1_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1543 = 6'h2 == fence_index ? 1'h0 : meta_2_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1544 = 6'h3 == fence_index ? 1'h0 : meta_3_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1545 = 6'h4 == fence_index ? 1'h0 : meta_4_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1546 = 6'h5 == fence_index ? 1'h0 : meta_5_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1547 = 6'h6 == fence_index ? 1'h0 : meta_6_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1548 = 6'h7 == fence_index ? 1'h0 : meta_7_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1549 = 6'h8 == fence_index ? 1'h0 : meta_8_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1550 = 6'h9 == fence_index ? 1'h0 : meta_9_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1551 = 6'ha == fence_index ? 1'h0 : meta_10_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1552 = 6'hb == fence_index ? 1'h0 : meta_11_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1553 = 6'hc == fence_index ? 1'h0 : meta_12_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1554 = 6'hd == fence_index ? 1'h0 : meta_13_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1555 = 6'he == fence_index ? 1'h0 : meta_14_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1556 = 6'hf == fence_index ? 1'h0 : meta_15_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1557 = 6'h10 == fence_index ? 1'h0 : meta_16_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1558 = 6'h11 == fence_index ? 1'h0 : meta_17_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1559 = 6'h12 == fence_index ? 1'h0 : meta_18_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1560 = 6'h13 == fence_index ? 1'h0 : meta_19_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1561 = 6'h14 == fence_index ? 1'h0 : meta_20_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1562 = 6'h15 == fence_index ? 1'h0 : meta_21_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1563 = 6'h16 == fence_index ? 1'h0 : meta_22_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1564 = 6'h17 == fence_index ? 1'h0 : meta_23_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1565 = 6'h18 == fence_index ? 1'h0 : meta_24_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1566 = 6'h19 == fence_index ? 1'h0 : meta_25_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1567 = 6'h1a == fence_index ? 1'h0 : meta_26_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1568 = 6'h1b == fence_index ? 1'h0 : meta_27_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1569 = 6'h1c == fence_index ? 1'h0 : meta_28_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1570 = 6'h1d == fence_index ? 1'h0 : meta_29_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1571 = 6'h1e == fence_index ? 1'h0 : meta_30_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1572 = 6'h1f == fence_index ? 1'h0 : meta_31_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1573 = 6'h20 == fence_index ? 1'h0 : meta_32_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1574 = 6'h21 == fence_index ? 1'h0 : meta_33_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1575 = 6'h22 == fence_index ? 1'h0 : meta_34_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1576 = 6'h23 == fence_index ? 1'h0 : meta_35_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1577 = 6'h24 == fence_index ? 1'h0 : meta_36_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1578 = 6'h25 == fence_index ? 1'h0 : meta_37_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1579 = 6'h26 == fence_index ? 1'h0 : meta_38_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1580 = 6'h27 == fence_index ? 1'h0 : meta_39_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1581 = 6'h28 == fence_index ? 1'h0 : meta_40_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1582 = 6'h29 == fence_index ? 1'h0 : meta_41_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1583 = 6'h2a == fence_index ? 1'h0 : meta_42_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1584 = 6'h2b == fence_index ? 1'h0 : meta_43_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1585 = 6'h2c == fence_index ? 1'h0 : meta_44_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1586 = 6'h2d == fence_index ? 1'h0 : meta_45_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1587 = 6'h2e == fence_index ? 1'h0 : meta_46_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1588 = 6'h2f == fence_index ? 1'h0 : meta_47_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1589 = 6'h30 == fence_index ? 1'h0 : meta_48_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1590 = 6'h31 == fence_index ? 1'h0 : meta_49_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1591 = 6'h32 == fence_index ? 1'h0 : meta_50_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1592 = 6'h33 == fence_index ? 1'h0 : meta_51_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1593 = 6'h34 == fence_index ? 1'h0 : meta_52_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1594 = 6'h35 == fence_index ? 1'h0 : meta_53_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1595 = 6'h36 == fence_index ? 1'h0 : meta_54_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1596 = 6'h37 == fence_index ? 1'h0 : meta_55_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1597 = 6'h38 == fence_index ? 1'h0 : meta_56_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1598 = 6'h39 == fence_index ? 1'h0 : meta_57_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1599 = 6'h3a == fence_index ? 1'h0 : meta_58_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1600 = 6'h3b == fence_index ? 1'h0 : meta_59_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1601 = 6'h3c == fence_index ? 1'h0 : meta_60_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1602 = 6'h3d == fence_index ? 1'h0 : meta_61_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1603 = 6'h3e == fence_index ? 1'h0 : meta_62_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1604 = 6'h3f == fence_index ? 1'h0 : meta_63_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1605 = 7'h40 == _GEN_14414 ? 1'h0 : meta_64_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1606 = 7'h41 == _GEN_14414 ? 1'h0 : meta_65_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1607 = 7'h42 == _GEN_14414 ? 1'h0 : meta_66_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1608 = 7'h43 == _GEN_14414 ? 1'h0 : meta_67_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1609 = 7'h44 == _GEN_14414 ? 1'h0 : meta_68_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1610 = 7'h45 == _GEN_14414 ? 1'h0 : meta_69_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1611 = 7'h46 == _GEN_14414 ? 1'h0 : meta_70_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1612 = 7'h47 == _GEN_14414 ? 1'h0 : meta_71_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1613 = 7'h48 == _GEN_14414 ? 1'h0 : meta_72_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1614 = 7'h49 == _GEN_14414 ? 1'h0 : meta_73_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1615 = 7'h4a == _GEN_14414 ? 1'h0 : meta_74_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1616 = 7'h4b == _GEN_14414 ? 1'h0 : meta_75_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1617 = 7'h4c == _GEN_14414 ? 1'h0 : meta_76_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1618 = 7'h4d == _GEN_14414 ? 1'h0 : meta_77_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1619 = 7'h4e == _GEN_14414 ? 1'h0 : meta_78_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1620 = 7'h4f == _GEN_14414 ? 1'h0 : meta_79_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1621 = 7'h50 == _GEN_14414 ? 1'h0 : meta_80_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1622 = 7'h51 == _GEN_14414 ? 1'h0 : meta_81_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1623 = 7'h52 == _GEN_14414 ? 1'h0 : meta_82_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1624 = 7'h53 == _GEN_14414 ? 1'h0 : meta_83_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1625 = 7'h54 == _GEN_14414 ? 1'h0 : meta_84_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1626 = 7'h55 == _GEN_14414 ? 1'h0 : meta_85_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1627 = 7'h56 == _GEN_14414 ? 1'h0 : meta_86_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1628 = 7'h57 == _GEN_14414 ? 1'h0 : meta_87_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1629 = 7'h58 == _GEN_14414 ? 1'h0 : meta_88_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1630 = 7'h59 == _GEN_14414 ? 1'h0 : meta_89_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1631 = 7'h5a == _GEN_14414 ? 1'h0 : meta_90_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1632 = 7'h5b == _GEN_14414 ? 1'h0 : meta_91_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1633 = 7'h5c == _GEN_14414 ? 1'h0 : meta_92_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1634 = 7'h5d == _GEN_14414 ? 1'h0 : meta_93_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1635 = 7'h5e == _GEN_14414 ? 1'h0 : meta_94_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1636 = 7'h5f == _GEN_14414 ? 1'h0 : meta_95_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1637 = 7'h60 == _GEN_14414 ? 1'h0 : meta_96_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1638 = 7'h61 == _GEN_14414 ? 1'h0 : meta_97_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1639 = 7'h62 == _GEN_14414 ? 1'h0 : meta_98_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1640 = 7'h63 == _GEN_14414 ? 1'h0 : meta_99_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1641 = 7'h64 == _GEN_14414 ? 1'h0 : meta_100_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1642 = 7'h65 == _GEN_14414 ? 1'h0 : meta_101_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1643 = 7'h66 == _GEN_14414 ? 1'h0 : meta_102_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1644 = 7'h67 == _GEN_14414 ? 1'h0 : meta_103_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1645 = 7'h68 == _GEN_14414 ? 1'h0 : meta_104_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1646 = 7'h69 == _GEN_14414 ? 1'h0 : meta_105_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1647 = 7'h6a == _GEN_14414 ? 1'h0 : meta_106_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1648 = 7'h6b == _GEN_14414 ? 1'h0 : meta_107_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1649 = 7'h6c == _GEN_14414 ? 1'h0 : meta_108_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1650 = 7'h6d == _GEN_14414 ? 1'h0 : meta_109_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1651 = 7'h6e == _GEN_14414 ? 1'h0 : meta_110_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1652 = 7'h6f == _GEN_14414 ? 1'h0 : meta_111_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1653 = 7'h70 == _GEN_14414 ? 1'h0 : meta_112_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1654 = 7'h71 == _GEN_14414 ? 1'h0 : meta_113_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1655 = 7'h72 == _GEN_14414 ? 1'h0 : meta_114_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1656 = 7'h73 == _GEN_14414 ? 1'h0 : meta_115_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1657 = 7'h74 == _GEN_14414 ? 1'h0 : meta_116_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1658 = 7'h75 == _GEN_14414 ? 1'h0 : meta_117_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1659 = 7'h76 == _GEN_14414 ? 1'h0 : meta_118_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1660 = 7'h77 == _GEN_14414 ? 1'h0 : meta_119_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1661 = 7'h78 == _GEN_14414 ? 1'h0 : meta_120_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1662 = 7'h79 == _GEN_14414 ? 1'h0 : meta_121_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1663 = 7'h7a == _GEN_14414 ? 1'h0 : meta_122_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1664 = 7'h7b == _GEN_14414 ? 1'h0 : meta_123_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1665 = 7'h7c == _GEN_14414 ? 1'h0 : meta_124_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1666 = 7'h7d == _GEN_14414 ? 1'h0 : meta_125_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1667 = 7'h7e == _GEN_14414 ? 1'h0 : meta_126_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1668 = 7'h7f == _GEN_14414 ? 1'h0 : meta_127_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1669 = 8'h80 == _GEN_14478 ? 1'h0 : meta_128_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1670 = 8'h81 == _GEN_14478 ? 1'h0 : meta_129_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1671 = 8'h82 == _GEN_14478 ? 1'h0 : meta_130_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1672 = 8'h83 == _GEN_14478 ? 1'h0 : meta_131_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1673 = 8'h84 == _GEN_14478 ? 1'h0 : meta_132_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1674 = 8'h85 == _GEN_14478 ? 1'h0 : meta_133_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1675 = 8'h86 == _GEN_14478 ? 1'h0 : meta_134_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1676 = 8'h87 == _GEN_14478 ? 1'h0 : meta_135_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1677 = 8'h88 == _GEN_14478 ? 1'h0 : meta_136_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1678 = 8'h89 == _GEN_14478 ? 1'h0 : meta_137_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1679 = 8'h8a == _GEN_14478 ? 1'h0 : meta_138_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1680 = 8'h8b == _GEN_14478 ? 1'h0 : meta_139_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1681 = 8'h8c == _GEN_14478 ? 1'h0 : meta_140_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1682 = 8'h8d == _GEN_14478 ? 1'h0 : meta_141_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1683 = 8'h8e == _GEN_14478 ? 1'h0 : meta_142_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1684 = 8'h8f == _GEN_14478 ? 1'h0 : meta_143_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1685 = 8'h90 == _GEN_14478 ? 1'h0 : meta_144_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1686 = 8'h91 == _GEN_14478 ? 1'h0 : meta_145_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1687 = 8'h92 == _GEN_14478 ? 1'h0 : meta_146_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1688 = 8'h93 == _GEN_14478 ? 1'h0 : meta_147_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1689 = 8'h94 == _GEN_14478 ? 1'h0 : meta_148_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1690 = 8'h95 == _GEN_14478 ? 1'h0 : meta_149_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1691 = 8'h96 == _GEN_14478 ? 1'h0 : meta_150_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1692 = 8'h97 == _GEN_14478 ? 1'h0 : meta_151_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1693 = 8'h98 == _GEN_14478 ? 1'h0 : meta_152_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1694 = 8'h99 == _GEN_14478 ? 1'h0 : meta_153_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1695 = 8'h9a == _GEN_14478 ? 1'h0 : meta_154_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1696 = 8'h9b == _GEN_14478 ? 1'h0 : meta_155_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1697 = 8'h9c == _GEN_14478 ? 1'h0 : meta_156_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1698 = 8'h9d == _GEN_14478 ? 1'h0 : meta_157_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1699 = 8'h9e == _GEN_14478 ? 1'h0 : meta_158_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1700 = 8'h9f == _GEN_14478 ? 1'h0 : meta_159_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1701 = 8'ha0 == _GEN_14478 ? 1'h0 : meta_160_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1702 = 8'ha1 == _GEN_14478 ? 1'h0 : meta_161_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1703 = 8'ha2 == _GEN_14478 ? 1'h0 : meta_162_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1704 = 8'ha3 == _GEN_14478 ? 1'h0 : meta_163_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1705 = 8'ha4 == _GEN_14478 ? 1'h0 : meta_164_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1706 = 8'ha5 == _GEN_14478 ? 1'h0 : meta_165_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1707 = 8'ha6 == _GEN_14478 ? 1'h0 : meta_166_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1708 = 8'ha7 == _GEN_14478 ? 1'h0 : meta_167_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1709 = 8'ha8 == _GEN_14478 ? 1'h0 : meta_168_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1710 = 8'ha9 == _GEN_14478 ? 1'h0 : meta_169_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1711 = 8'haa == _GEN_14478 ? 1'h0 : meta_170_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1712 = 8'hab == _GEN_14478 ? 1'h0 : meta_171_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1713 = 8'hac == _GEN_14478 ? 1'h0 : meta_172_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1714 = 8'had == _GEN_14478 ? 1'h0 : meta_173_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1715 = 8'hae == _GEN_14478 ? 1'h0 : meta_174_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1716 = 8'haf == _GEN_14478 ? 1'h0 : meta_175_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1717 = 8'hb0 == _GEN_14478 ? 1'h0 : meta_176_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1718 = 8'hb1 == _GEN_14478 ? 1'h0 : meta_177_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1719 = 8'hb2 == _GEN_14478 ? 1'h0 : meta_178_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1720 = 8'hb3 == _GEN_14478 ? 1'h0 : meta_179_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1721 = 8'hb4 == _GEN_14478 ? 1'h0 : meta_180_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1722 = 8'hb5 == _GEN_14478 ? 1'h0 : meta_181_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1723 = 8'hb6 == _GEN_14478 ? 1'h0 : meta_182_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1724 = 8'hb7 == _GEN_14478 ? 1'h0 : meta_183_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1725 = 8'hb8 == _GEN_14478 ? 1'h0 : meta_184_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1726 = 8'hb9 == _GEN_14478 ? 1'h0 : meta_185_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1727 = 8'hba == _GEN_14478 ? 1'h0 : meta_186_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1728 = 8'hbb == _GEN_14478 ? 1'h0 : meta_187_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1729 = 8'hbc == _GEN_14478 ? 1'h0 : meta_188_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1730 = 8'hbd == _GEN_14478 ? 1'h0 : meta_189_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1731 = 8'hbe == _GEN_14478 ? 1'h0 : meta_190_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1732 = 8'hbf == _GEN_14478 ? 1'h0 : meta_191_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1733 = 8'hc0 == _GEN_14478 ? 1'h0 : meta_192_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1734 = 8'hc1 == _GEN_14478 ? 1'h0 : meta_193_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1735 = 8'hc2 == _GEN_14478 ? 1'h0 : meta_194_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1736 = 8'hc3 == _GEN_14478 ? 1'h0 : meta_195_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1737 = 8'hc4 == _GEN_14478 ? 1'h0 : meta_196_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1738 = 8'hc5 == _GEN_14478 ? 1'h0 : meta_197_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1739 = 8'hc6 == _GEN_14478 ? 1'h0 : meta_198_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1740 = 8'hc7 == _GEN_14478 ? 1'h0 : meta_199_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1741 = 8'hc8 == _GEN_14478 ? 1'h0 : meta_200_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1742 = 8'hc9 == _GEN_14478 ? 1'h0 : meta_201_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1743 = 8'hca == _GEN_14478 ? 1'h0 : meta_202_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1744 = 8'hcb == _GEN_14478 ? 1'h0 : meta_203_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1745 = 8'hcc == _GEN_14478 ? 1'h0 : meta_204_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1746 = 8'hcd == _GEN_14478 ? 1'h0 : meta_205_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1747 = 8'hce == _GEN_14478 ? 1'h0 : meta_206_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1748 = 8'hcf == _GEN_14478 ? 1'h0 : meta_207_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1749 = 8'hd0 == _GEN_14478 ? 1'h0 : meta_208_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1750 = 8'hd1 == _GEN_14478 ? 1'h0 : meta_209_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1751 = 8'hd2 == _GEN_14478 ? 1'h0 : meta_210_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1752 = 8'hd3 == _GEN_14478 ? 1'h0 : meta_211_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1753 = 8'hd4 == _GEN_14478 ? 1'h0 : meta_212_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1754 = 8'hd5 == _GEN_14478 ? 1'h0 : meta_213_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1755 = 8'hd6 == _GEN_14478 ? 1'h0 : meta_214_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1756 = 8'hd7 == _GEN_14478 ? 1'h0 : meta_215_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1757 = 8'hd8 == _GEN_14478 ? 1'h0 : meta_216_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1758 = 8'hd9 == _GEN_14478 ? 1'h0 : meta_217_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1759 = 8'hda == _GEN_14478 ? 1'h0 : meta_218_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1760 = 8'hdb == _GEN_14478 ? 1'h0 : meta_219_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1761 = 8'hdc == _GEN_14478 ? 1'h0 : meta_220_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1762 = 8'hdd == _GEN_14478 ? 1'h0 : meta_221_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1763 = 8'hde == _GEN_14478 ? 1'h0 : meta_222_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1764 = 8'hdf == _GEN_14478 ? 1'h0 : meta_223_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1765 = 8'he0 == _GEN_14478 ? 1'h0 : meta_224_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1766 = 8'he1 == _GEN_14478 ? 1'h0 : meta_225_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1767 = 8'he2 == _GEN_14478 ? 1'h0 : meta_226_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1768 = 8'he3 == _GEN_14478 ? 1'h0 : meta_227_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1769 = 8'he4 == _GEN_14478 ? 1'h0 : meta_228_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1770 = 8'he5 == _GEN_14478 ? 1'h0 : meta_229_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1771 = 8'he6 == _GEN_14478 ? 1'h0 : meta_230_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1772 = 8'he7 == _GEN_14478 ? 1'h0 : meta_231_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1773 = 8'he8 == _GEN_14478 ? 1'h0 : meta_232_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1774 = 8'he9 == _GEN_14478 ? 1'h0 : meta_233_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1775 = 8'hea == _GEN_14478 ? 1'h0 : meta_234_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1776 = 8'heb == _GEN_14478 ? 1'h0 : meta_235_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1777 = 8'hec == _GEN_14478 ? 1'h0 : meta_236_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1778 = 8'hed == _GEN_14478 ? 1'h0 : meta_237_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1779 = 8'hee == _GEN_14478 ? 1'h0 : meta_238_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1780 = 8'hef == _GEN_14478 ? 1'h0 : meta_239_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1781 = 8'hf0 == _GEN_14478 ? 1'h0 : meta_240_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1782 = 8'hf1 == _GEN_14478 ? 1'h0 : meta_241_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1783 = 8'hf2 == _GEN_14478 ? 1'h0 : meta_242_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1784 = 8'hf3 == _GEN_14478 ? 1'h0 : meta_243_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1785 = 8'hf4 == _GEN_14478 ? 1'h0 : meta_244_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1786 = 8'hf5 == _GEN_14478 ? 1'h0 : meta_245_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1787 = 8'hf6 == _GEN_14478 ? 1'h0 : meta_246_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1788 = 8'hf7 == _GEN_14478 ? 1'h0 : meta_247_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1789 = 8'hf8 == _GEN_14478 ? 1'h0 : meta_248_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1790 = 8'hf9 == _GEN_14478 ? 1'h0 : meta_249_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1791 = 8'hfa == _GEN_14478 ? 1'h0 : meta_250_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1792 = 8'hfb == _GEN_14478 ? 1'h0 : meta_251_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1793 = 8'hfc == _GEN_14478 ? 1'h0 : meta_252_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1794 = 8'hfd == _GEN_14478 ? 1'h0 : meta_253_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1795 = 8'hfe == _GEN_14478 ? 1'h0 : meta_254_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1796 = 8'hff == _GEN_14478 ? 1'h0 : meta_255_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1797 = 9'h100 == _GEN_14606 ? 1'h0 : meta_256_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1798 = 9'h101 == _GEN_14606 ? 1'h0 : meta_257_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1799 = 9'h102 == _GEN_14606 ? 1'h0 : meta_258_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1800 = 9'h103 == _GEN_14606 ? 1'h0 : meta_259_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1801 = 9'h104 == _GEN_14606 ? 1'h0 : meta_260_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1802 = 9'h105 == _GEN_14606 ? 1'h0 : meta_261_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1803 = 9'h106 == _GEN_14606 ? 1'h0 : meta_262_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1804 = 9'h107 == _GEN_14606 ? 1'h0 : meta_263_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1805 = 9'h108 == _GEN_14606 ? 1'h0 : meta_264_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1806 = 9'h109 == _GEN_14606 ? 1'h0 : meta_265_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1807 = 9'h10a == _GEN_14606 ? 1'h0 : meta_266_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1808 = 9'h10b == _GEN_14606 ? 1'h0 : meta_267_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1809 = 9'h10c == _GEN_14606 ? 1'h0 : meta_268_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1810 = 9'h10d == _GEN_14606 ? 1'h0 : meta_269_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1811 = 9'h10e == _GEN_14606 ? 1'h0 : meta_270_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1812 = 9'h10f == _GEN_14606 ? 1'h0 : meta_271_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1813 = 9'h110 == _GEN_14606 ? 1'h0 : meta_272_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1814 = 9'h111 == _GEN_14606 ? 1'h0 : meta_273_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1815 = 9'h112 == _GEN_14606 ? 1'h0 : meta_274_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1816 = 9'h113 == _GEN_14606 ? 1'h0 : meta_275_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1817 = 9'h114 == _GEN_14606 ? 1'h0 : meta_276_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1818 = 9'h115 == _GEN_14606 ? 1'h0 : meta_277_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1819 = 9'h116 == _GEN_14606 ? 1'h0 : meta_278_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1820 = 9'h117 == _GEN_14606 ? 1'h0 : meta_279_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1821 = 9'h118 == _GEN_14606 ? 1'h0 : meta_280_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1822 = 9'h119 == _GEN_14606 ? 1'h0 : meta_281_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1823 = 9'h11a == _GEN_14606 ? 1'h0 : meta_282_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1824 = 9'h11b == _GEN_14606 ? 1'h0 : meta_283_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1825 = 9'h11c == _GEN_14606 ? 1'h0 : meta_284_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1826 = 9'h11d == _GEN_14606 ? 1'h0 : meta_285_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1827 = 9'h11e == _GEN_14606 ? 1'h0 : meta_286_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1828 = 9'h11f == _GEN_14606 ? 1'h0 : meta_287_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1829 = 9'h120 == _GEN_14606 ? 1'h0 : meta_288_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1830 = 9'h121 == _GEN_14606 ? 1'h0 : meta_289_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1831 = 9'h122 == _GEN_14606 ? 1'h0 : meta_290_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1832 = 9'h123 == _GEN_14606 ? 1'h0 : meta_291_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1833 = 9'h124 == _GEN_14606 ? 1'h0 : meta_292_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1834 = 9'h125 == _GEN_14606 ? 1'h0 : meta_293_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1835 = 9'h126 == _GEN_14606 ? 1'h0 : meta_294_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1836 = 9'h127 == _GEN_14606 ? 1'h0 : meta_295_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1837 = 9'h128 == _GEN_14606 ? 1'h0 : meta_296_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1838 = 9'h129 == _GEN_14606 ? 1'h0 : meta_297_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1839 = 9'h12a == _GEN_14606 ? 1'h0 : meta_298_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1840 = 9'h12b == _GEN_14606 ? 1'h0 : meta_299_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1841 = 9'h12c == _GEN_14606 ? 1'h0 : meta_300_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1842 = 9'h12d == _GEN_14606 ? 1'h0 : meta_301_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1843 = 9'h12e == _GEN_14606 ? 1'h0 : meta_302_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1844 = 9'h12f == _GEN_14606 ? 1'h0 : meta_303_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1845 = 9'h130 == _GEN_14606 ? 1'h0 : meta_304_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1846 = 9'h131 == _GEN_14606 ? 1'h0 : meta_305_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1847 = 9'h132 == _GEN_14606 ? 1'h0 : meta_306_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1848 = 9'h133 == _GEN_14606 ? 1'h0 : meta_307_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1849 = 9'h134 == _GEN_14606 ? 1'h0 : meta_308_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1850 = 9'h135 == _GEN_14606 ? 1'h0 : meta_309_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1851 = 9'h136 == _GEN_14606 ? 1'h0 : meta_310_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1852 = 9'h137 == _GEN_14606 ? 1'h0 : meta_311_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1853 = 9'h138 == _GEN_14606 ? 1'h0 : meta_312_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1854 = 9'h139 == _GEN_14606 ? 1'h0 : meta_313_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1855 = 9'h13a == _GEN_14606 ? 1'h0 : meta_314_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1856 = 9'h13b == _GEN_14606 ? 1'h0 : meta_315_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1857 = 9'h13c == _GEN_14606 ? 1'h0 : meta_316_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1858 = 9'h13d == _GEN_14606 ? 1'h0 : meta_317_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1859 = 9'h13e == _GEN_14606 ? 1'h0 : meta_318_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1860 = 9'h13f == _GEN_14606 ? 1'h0 : meta_319_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1861 = 9'h140 == _GEN_14606 ? 1'h0 : meta_320_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1862 = 9'h141 == _GEN_14606 ? 1'h0 : meta_321_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1863 = 9'h142 == _GEN_14606 ? 1'h0 : meta_322_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1864 = 9'h143 == _GEN_14606 ? 1'h0 : meta_323_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1865 = 9'h144 == _GEN_14606 ? 1'h0 : meta_324_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1866 = 9'h145 == _GEN_14606 ? 1'h0 : meta_325_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1867 = 9'h146 == _GEN_14606 ? 1'h0 : meta_326_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1868 = 9'h147 == _GEN_14606 ? 1'h0 : meta_327_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1869 = 9'h148 == _GEN_14606 ? 1'h0 : meta_328_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1870 = 9'h149 == _GEN_14606 ? 1'h0 : meta_329_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1871 = 9'h14a == _GEN_14606 ? 1'h0 : meta_330_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1872 = 9'h14b == _GEN_14606 ? 1'h0 : meta_331_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1873 = 9'h14c == _GEN_14606 ? 1'h0 : meta_332_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1874 = 9'h14d == _GEN_14606 ? 1'h0 : meta_333_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1875 = 9'h14e == _GEN_14606 ? 1'h0 : meta_334_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1876 = 9'h14f == _GEN_14606 ? 1'h0 : meta_335_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1877 = 9'h150 == _GEN_14606 ? 1'h0 : meta_336_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1878 = 9'h151 == _GEN_14606 ? 1'h0 : meta_337_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1879 = 9'h152 == _GEN_14606 ? 1'h0 : meta_338_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1880 = 9'h153 == _GEN_14606 ? 1'h0 : meta_339_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1881 = 9'h154 == _GEN_14606 ? 1'h0 : meta_340_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1882 = 9'h155 == _GEN_14606 ? 1'h0 : meta_341_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1883 = 9'h156 == _GEN_14606 ? 1'h0 : meta_342_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1884 = 9'h157 == _GEN_14606 ? 1'h0 : meta_343_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1885 = 9'h158 == _GEN_14606 ? 1'h0 : meta_344_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1886 = 9'h159 == _GEN_14606 ? 1'h0 : meta_345_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1887 = 9'h15a == _GEN_14606 ? 1'h0 : meta_346_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1888 = 9'h15b == _GEN_14606 ? 1'h0 : meta_347_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1889 = 9'h15c == _GEN_14606 ? 1'h0 : meta_348_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1890 = 9'h15d == _GEN_14606 ? 1'h0 : meta_349_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1891 = 9'h15e == _GEN_14606 ? 1'h0 : meta_350_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1892 = 9'h15f == _GEN_14606 ? 1'h0 : meta_351_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1893 = 9'h160 == _GEN_14606 ? 1'h0 : meta_352_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1894 = 9'h161 == _GEN_14606 ? 1'h0 : meta_353_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1895 = 9'h162 == _GEN_14606 ? 1'h0 : meta_354_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1896 = 9'h163 == _GEN_14606 ? 1'h0 : meta_355_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1897 = 9'h164 == _GEN_14606 ? 1'h0 : meta_356_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1898 = 9'h165 == _GEN_14606 ? 1'h0 : meta_357_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1899 = 9'h166 == _GEN_14606 ? 1'h0 : meta_358_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1900 = 9'h167 == _GEN_14606 ? 1'h0 : meta_359_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1901 = 9'h168 == _GEN_14606 ? 1'h0 : meta_360_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1902 = 9'h169 == _GEN_14606 ? 1'h0 : meta_361_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1903 = 9'h16a == _GEN_14606 ? 1'h0 : meta_362_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1904 = 9'h16b == _GEN_14606 ? 1'h0 : meta_363_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1905 = 9'h16c == _GEN_14606 ? 1'h0 : meta_364_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1906 = 9'h16d == _GEN_14606 ? 1'h0 : meta_365_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1907 = 9'h16e == _GEN_14606 ? 1'h0 : meta_366_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1908 = 9'h16f == _GEN_14606 ? 1'h0 : meta_367_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1909 = 9'h170 == _GEN_14606 ? 1'h0 : meta_368_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1910 = 9'h171 == _GEN_14606 ? 1'h0 : meta_369_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1911 = 9'h172 == _GEN_14606 ? 1'h0 : meta_370_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1912 = 9'h173 == _GEN_14606 ? 1'h0 : meta_371_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1913 = 9'h174 == _GEN_14606 ? 1'h0 : meta_372_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1914 = 9'h175 == _GEN_14606 ? 1'h0 : meta_373_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1915 = 9'h176 == _GEN_14606 ? 1'h0 : meta_374_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1916 = 9'h177 == _GEN_14606 ? 1'h0 : meta_375_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1917 = 9'h178 == _GEN_14606 ? 1'h0 : meta_376_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1918 = 9'h179 == _GEN_14606 ? 1'h0 : meta_377_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1919 = 9'h17a == _GEN_14606 ? 1'h0 : meta_378_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1920 = 9'h17b == _GEN_14606 ? 1'h0 : meta_379_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1921 = 9'h17c == _GEN_14606 ? 1'h0 : meta_380_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1922 = 9'h17d == _GEN_14606 ? 1'h0 : meta_381_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1923 = 9'h17e == _GEN_14606 ? 1'h0 : meta_382_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1924 = 9'h17f == _GEN_14606 ? 1'h0 : meta_383_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1925 = 9'h180 == _GEN_14606 ? 1'h0 : meta_384_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1926 = 9'h181 == _GEN_14606 ? 1'h0 : meta_385_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1927 = 9'h182 == _GEN_14606 ? 1'h0 : meta_386_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1928 = 9'h183 == _GEN_14606 ? 1'h0 : meta_387_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1929 = 9'h184 == _GEN_14606 ? 1'h0 : meta_388_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1930 = 9'h185 == _GEN_14606 ? 1'h0 : meta_389_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1931 = 9'h186 == _GEN_14606 ? 1'h0 : meta_390_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1932 = 9'h187 == _GEN_14606 ? 1'h0 : meta_391_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1933 = 9'h188 == _GEN_14606 ? 1'h0 : meta_392_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1934 = 9'h189 == _GEN_14606 ? 1'h0 : meta_393_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1935 = 9'h18a == _GEN_14606 ? 1'h0 : meta_394_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1936 = 9'h18b == _GEN_14606 ? 1'h0 : meta_395_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1937 = 9'h18c == _GEN_14606 ? 1'h0 : meta_396_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1938 = 9'h18d == _GEN_14606 ? 1'h0 : meta_397_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1939 = 9'h18e == _GEN_14606 ? 1'h0 : meta_398_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1940 = 9'h18f == _GEN_14606 ? 1'h0 : meta_399_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1941 = 9'h190 == _GEN_14606 ? 1'h0 : meta_400_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1942 = 9'h191 == _GEN_14606 ? 1'h0 : meta_401_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1943 = 9'h192 == _GEN_14606 ? 1'h0 : meta_402_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1944 = 9'h193 == _GEN_14606 ? 1'h0 : meta_403_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1945 = 9'h194 == _GEN_14606 ? 1'h0 : meta_404_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1946 = 9'h195 == _GEN_14606 ? 1'h0 : meta_405_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1947 = 9'h196 == _GEN_14606 ? 1'h0 : meta_406_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1948 = 9'h197 == _GEN_14606 ? 1'h0 : meta_407_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1949 = 9'h198 == _GEN_14606 ? 1'h0 : meta_408_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1950 = 9'h199 == _GEN_14606 ? 1'h0 : meta_409_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1951 = 9'h19a == _GEN_14606 ? 1'h0 : meta_410_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1952 = 9'h19b == _GEN_14606 ? 1'h0 : meta_411_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1953 = 9'h19c == _GEN_14606 ? 1'h0 : meta_412_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1954 = 9'h19d == _GEN_14606 ? 1'h0 : meta_413_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1955 = 9'h19e == _GEN_14606 ? 1'h0 : meta_414_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1956 = 9'h19f == _GEN_14606 ? 1'h0 : meta_415_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1957 = 9'h1a0 == _GEN_14606 ? 1'h0 : meta_416_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1958 = 9'h1a1 == _GEN_14606 ? 1'h0 : meta_417_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1959 = 9'h1a2 == _GEN_14606 ? 1'h0 : meta_418_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1960 = 9'h1a3 == _GEN_14606 ? 1'h0 : meta_419_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1961 = 9'h1a4 == _GEN_14606 ? 1'h0 : meta_420_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1962 = 9'h1a5 == _GEN_14606 ? 1'h0 : meta_421_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1963 = 9'h1a6 == _GEN_14606 ? 1'h0 : meta_422_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1964 = 9'h1a7 == _GEN_14606 ? 1'h0 : meta_423_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1965 = 9'h1a8 == _GEN_14606 ? 1'h0 : meta_424_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1966 = 9'h1a9 == _GEN_14606 ? 1'h0 : meta_425_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1967 = 9'h1aa == _GEN_14606 ? 1'h0 : meta_426_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1968 = 9'h1ab == _GEN_14606 ? 1'h0 : meta_427_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1969 = 9'h1ac == _GEN_14606 ? 1'h0 : meta_428_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1970 = 9'h1ad == _GEN_14606 ? 1'h0 : meta_429_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1971 = 9'h1ae == _GEN_14606 ? 1'h0 : meta_430_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1972 = 9'h1af == _GEN_14606 ? 1'h0 : meta_431_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1973 = 9'h1b0 == _GEN_14606 ? 1'h0 : meta_432_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1974 = 9'h1b1 == _GEN_14606 ? 1'h0 : meta_433_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1975 = 9'h1b2 == _GEN_14606 ? 1'h0 : meta_434_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1976 = 9'h1b3 == _GEN_14606 ? 1'h0 : meta_435_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1977 = 9'h1b4 == _GEN_14606 ? 1'h0 : meta_436_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1978 = 9'h1b5 == _GEN_14606 ? 1'h0 : meta_437_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1979 = 9'h1b6 == _GEN_14606 ? 1'h0 : meta_438_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1980 = 9'h1b7 == _GEN_14606 ? 1'h0 : meta_439_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1981 = 9'h1b8 == _GEN_14606 ? 1'h0 : meta_440_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1982 = 9'h1b9 == _GEN_14606 ? 1'h0 : meta_441_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1983 = 9'h1ba == _GEN_14606 ? 1'h0 : meta_442_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1984 = 9'h1bb == _GEN_14606 ? 1'h0 : meta_443_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1985 = 9'h1bc == _GEN_14606 ? 1'h0 : meta_444_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1986 = 9'h1bd == _GEN_14606 ? 1'h0 : meta_445_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1987 = 9'h1be == _GEN_14606 ? 1'h0 : meta_446_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1988 = 9'h1bf == _GEN_14606 ? 1'h0 : meta_447_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1989 = 9'h1c0 == _GEN_14606 ? 1'h0 : meta_448_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1990 = 9'h1c1 == _GEN_14606 ? 1'h0 : meta_449_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1991 = 9'h1c2 == _GEN_14606 ? 1'h0 : meta_450_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1992 = 9'h1c3 == _GEN_14606 ? 1'h0 : meta_451_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1993 = 9'h1c4 == _GEN_14606 ? 1'h0 : meta_452_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1994 = 9'h1c5 == _GEN_14606 ? 1'h0 : meta_453_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1995 = 9'h1c6 == _GEN_14606 ? 1'h0 : meta_454_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1996 = 9'h1c7 == _GEN_14606 ? 1'h0 : meta_455_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1997 = 9'h1c8 == _GEN_14606 ? 1'h0 : meta_456_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1998 = 9'h1c9 == _GEN_14606 ? 1'h0 : meta_457_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_1999 = 9'h1ca == _GEN_14606 ? 1'h0 : meta_458_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2000 = 9'h1cb == _GEN_14606 ? 1'h0 : meta_459_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2001 = 9'h1cc == _GEN_14606 ? 1'h0 : meta_460_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2002 = 9'h1cd == _GEN_14606 ? 1'h0 : meta_461_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2003 = 9'h1ce == _GEN_14606 ? 1'h0 : meta_462_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2004 = 9'h1cf == _GEN_14606 ? 1'h0 : meta_463_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2005 = 9'h1d0 == _GEN_14606 ? 1'h0 : meta_464_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2006 = 9'h1d1 == _GEN_14606 ? 1'h0 : meta_465_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2007 = 9'h1d2 == _GEN_14606 ? 1'h0 : meta_466_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2008 = 9'h1d3 == _GEN_14606 ? 1'h0 : meta_467_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2009 = 9'h1d4 == _GEN_14606 ? 1'h0 : meta_468_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2010 = 9'h1d5 == _GEN_14606 ? 1'h0 : meta_469_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2011 = 9'h1d6 == _GEN_14606 ? 1'h0 : meta_470_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2012 = 9'h1d7 == _GEN_14606 ? 1'h0 : meta_471_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2013 = 9'h1d8 == _GEN_14606 ? 1'h0 : meta_472_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2014 = 9'h1d9 == _GEN_14606 ? 1'h0 : meta_473_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2015 = 9'h1da == _GEN_14606 ? 1'h0 : meta_474_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2016 = 9'h1db == _GEN_14606 ? 1'h0 : meta_475_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2017 = 9'h1dc == _GEN_14606 ? 1'h0 : meta_476_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2018 = 9'h1dd == _GEN_14606 ? 1'h0 : meta_477_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2019 = 9'h1de == _GEN_14606 ? 1'h0 : meta_478_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2020 = 9'h1df == _GEN_14606 ? 1'h0 : meta_479_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2021 = 9'h1e0 == _GEN_14606 ? 1'h0 : meta_480_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2022 = 9'h1e1 == _GEN_14606 ? 1'h0 : meta_481_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2023 = 9'h1e2 == _GEN_14606 ? 1'h0 : meta_482_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2024 = 9'h1e3 == _GEN_14606 ? 1'h0 : meta_483_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2025 = 9'h1e4 == _GEN_14606 ? 1'h0 : meta_484_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2026 = 9'h1e5 == _GEN_14606 ? 1'h0 : meta_485_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2027 = 9'h1e6 == _GEN_14606 ? 1'h0 : meta_486_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2028 = 9'h1e7 == _GEN_14606 ? 1'h0 : meta_487_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2029 = 9'h1e8 == _GEN_14606 ? 1'h0 : meta_488_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2030 = 9'h1e9 == _GEN_14606 ? 1'h0 : meta_489_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2031 = 9'h1ea == _GEN_14606 ? 1'h0 : meta_490_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2032 = 9'h1eb == _GEN_14606 ? 1'h0 : meta_491_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2033 = 9'h1ec == _GEN_14606 ? 1'h0 : meta_492_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2034 = 9'h1ed == _GEN_14606 ? 1'h0 : meta_493_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2035 = 9'h1ee == _GEN_14606 ? 1'h0 : meta_494_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2036 = 9'h1ef == _GEN_14606 ? 1'h0 : meta_495_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2037 = 9'h1f0 == _GEN_14606 ? 1'h0 : meta_496_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2038 = 9'h1f1 == _GEN_14606 ? 1'h0 : meta_497_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2039 = 9'h1f2 == _GEN_14606 ? 1'h0 : meta_498_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2040 = 9'h1f3 == _GEN_14606 ? 1'h0 : meta_499_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2041 = 9'h1f4 == _GEN_14606 ? 1'h0 : meta_500_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2042 = 9'h1f5 == _GEN_14606 ? 1'h0 : meta_501_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2043 = 9'h1f6 == _GEN_14606 ? 1'h0 : meta_502_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2044 = 9'h1f7 == _GEN_14606 ? 1'h0 : meta_503_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2045 = 9'h1f8 == _GEN_14606 ? 1'h0 : meta_504_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2046 = 9'h1f9 == _GEN_14606 ? 1'h0 : meta_505_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2047 = 9'h1fa == _GEN_14606 ? 1'h0 : meta_506_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2048 = 9'h1fb == _GEN_14606 ? 1'h0 : meta_507_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2049 = 9'h1fc == _GEN_14606 ? 1'h0 : meta_508_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2050 = 9'h1fd == _GEN_14606 ? 1'h0 : meta_509_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2051 = 9'h1fe == _GEN_14606 ? 1'h0 : meta_510_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2052 = 9'h1ff == _GEN_14606 ? 1'h0 : meta_511_valid_1; // @[ICache.scala 138:{32,32} 34:21]
  wire  _GEN_2053 = io_cpu_fence_value & _T & _T_2 ? _GEN_1029 : meta_0_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2054 = io_cpu_fence_value & _T & _T_2 ? _GEN_1030 : meta_1_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2055 = io_cpu_fence_value & _T & _T_2 ? _GEN_1031 : meta_2_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2056 = io_cpu_fence_value & _T & _T_2 ? _GEN_1032 : meta_3_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2057 = io_cpu_fence_value & _T & _T_2 ? _GEN_1033 : meta_4_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2058 = io_cpu_fence_value & _T & _T_2 ? _GEN_1034 : meta_5_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2059 = io_cpu_fence_value & _T & _T_2 ? _GEN_1035 : meta_6_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2060 = io_cpu_fence_value & _T & _T_2 ? _GEN_1036 : meta_7_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2061 = io_cpu_fence_value & _T & _T_2 ? _GEN_1037 : meta_8_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2062 = io_cpu_fence_value & _T & _T_2 ? _GEN_1038 : meta_9_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2063 = io_cpu_fence_value & _T & _T_2 ? _GEN_1039 : meta_10_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2064 = io_cpu_fence_value & _T & _T_2 ? _GEN_1040 : meta_11_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2065 = io_cpu_fence_value & _T & _T_2 ? _GEN_1041 : meta_12_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2066 = io_cpu_fence_value & _T & _T_2 ? _GEN_1042 : meta_13_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2067 = io_cpu_fence_value & _T & _T_2 ? _GEN_1043 : meta_14_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2068 = io_cpu_fence_value & _T & _T_2 ? _GEN_1044 : meta_15_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2069 = io_cpu_fence_value & _T & _T_2 ? _GEN_1045 : meta_16_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2070 = io_cpu_fence_value & _T & _T_2 ? _GEN_1046 : meta_17_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2071 = io_cpu_fence_value & _T & _T_2 ? _GEN_1047 : meta_18_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2072 = io_cpu_fence_value & _T & _T_2 ? _GEN_1048 : meta_19_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2073 = io_cpu_fence_value & _T & _T_2 ? _GEN_1049 : meta_20_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2074 = io_cpu_fence_value & _T & _T_2 ? _GEN_1050 : meta_21_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2075 = io_cpu_fence_value & _T & _T_2 ? _GEN_1051 : meta_22_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2076 = io_cpu_fence_value & _T & _T_2 ? _GEN_1052 : meta_23_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2077 = io_cpu_fence_value & _T & _T_2 ? _GEN_1053 : meta_24_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2078 = io_cpu_fence_value & _T & _T_2 ? _GEN_1054 : meta_25_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2079 = io_cpu_fence_value & _T & _T_2 ? _GEN_1055 : meta_26_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2080 = io_cpu_fence_value & _T & _T_2 ? _GEN_1056 : meta_27_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2081 = io_cpu_fence_value & _T & _T_2 ? _GEN_1057 : meta_28_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2082 = io_cpu_fence_value & _T & _T_2 ? _GEN_1058 : meta_29_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2083 = io_cpu_fence_value & _T & _T_2 ? _GEN_1059 : meta_30_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2084 = io_cpu_fence_value & _T & _T_2 ? _GEN_1060 : meta_31_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2085 = io_cpu_fence_value & _T & _T_2 ? _GEN_1061 : meta_32_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2086 = io_cpu_fence_value & _T & _T_2 ? _GEN_1062 : meta_33_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2087 = io_cpu_fence_value & _T & _T_2 ? _GEN_1063 : meta_34_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2088 = io_cpu_fence_value & _T & _T_2 ? _GEN_1064 : meta_35_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2089 = io_cpu_fence_value & _T & _T_2 ? _GEN_1065 : meta_36_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2090 = io_cpu_fence_value & _T & _T_2 ? _GEN_1066 : meta_37_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2091 = io_cpu_fence_value & _T & _T_2 ? _GEN_1067 : meta_38_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2092 = io_cpu_fence_value & _T & _T_2 ? _GEN_1068 : meta_39_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2093 = io_cpu_fence_value & _T & _T_2 ? _GEN_1069 : meta_40_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2094 = io_cpu_fence_value & _T & _T_2 ? _GEN_1070 : meta_41_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2095 = io_cpu_fence_value & _T & _T_2 ? _GEN_1071 : meta_42_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2096 = io_cpu_fence_value & _T & _T_2 ? _GEN_1072 : meta_43_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2097 = io_cpu_fence_value & _T & _T_2 ? _GEN_1073 : meta_44_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2098 = io_cpu_fence_value & _T & _T_2 ? _GEN_1074 : meta_45_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2099 = io_cpu_fence_value & _T & _T_2 ? _GEN_1075 : meta_46_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2100 = io_cpu_fence_value & _T & _T_2 ? _GEN_1076 : meta_47_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2101 = io_cpu_fence_value & _T & _T_2 ? _GEN_1077 : meta_48_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2102 = io_cpu_fence_value & _T & _T_2 ? _GEN_1078 : meta_49_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2103 = io_cpu_fence_value & _T & _T_2 ? _GEN_1079 : meta_50_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2104 = io_cpu_fence_value & _T & _T_2 ? _GEN_1080 : meta_51_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2105 = io_cpu_fence_value & _T & _T_2 ? _GEN_1081 : meta_52_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2106 = io_cpu_fence_value & _T & _T_2 ? _GEN_1082 : meta_53_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2107 = io_cpu_fence_value & _T & _T_2 ? _GEN_1083 : meta_54_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2108 = io_cpu_fence_value & _T & _T_2 ? _GEN_1084 : meta_55_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2109 = io_cpu_fence_value & _T & _T_2 ? _GEN_1085 : meta_56_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2110 = io_cpu_fence_value & _T & _T_2 ? _GEN_1086 : meta_57_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2111 = io_cpu_fence_value & _T & _T_2 ? _GEN_1087 : meta_58_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2112 = io_cpu_fence_value & _T & _T_2 ? _GEN_1088 : meta_59_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2113 = io_cpu_fence_value & _T & _T_2 ? _GEN_1089 : meta_60_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2114 = io_cpu_fence_value & _T & _T_2 ? _GEN_1090 : meta_61_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2115 = io_cpu_fence_value & _T & _T_2 ? _GEN_1091 : meta_62_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2116 = io_cpu_fence_value & _T & _T_2 ? _GEN_1092 : meta_63_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2117 = io_cpu_fence_value & _T & _T_2 ? _GEN_1093 : meta_64_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2118 = io_cpu_fence_value & _T & _T_2 ? _GEN_1094 : meta_65_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2119 = io_cpu_fence_value & _T & _T_2 ? _GEN_1095 : meta_66_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2120 = io_cpu_fence_value & _T & _T_2 ? _GEN_1096 : meta_67_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2121 = io_cpu_fence_value & _T & _T_2 ? _GEN_1097 : meta_68_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2122 = io_cpu_fence_value & _T & _T_2 ? _GEN_1098 : meta_69_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2123 = io_cpu_fence_value & _T & _T_2 ? _GEN_1099 : meta_70_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2124 = io_cpu_fence_value & _T & _T_2 ? _GEN_1100 : meta_71_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2125 = io_cpu_fence_value & _T & _T_2 ? _GEN_1101 : meta_72_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2126 = io_cpu_fence_value & _T & _T_2 ? _GEN_1102 : meta_73_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2127 = io_cpu_fence_value & _T & _T_2 ? _GEN_1103 : meta_74_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2128 = io_cpu_fence_value & _T & _T_2 ? _GEN_1104 : meta_75_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2129 = io_cpu_fence_value & _T & _T_2 ? _GEN_1105 : meta_76_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2130 = io_cpu_fence_value & _T & _T_2 ? _GEN_1106 : meta_77_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2131 = io_cpu_fence_value & _T & _T_2 ? _GEN_1107 : meta_78_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2132 = io_cpu_fence_value & _T & _T_2 ? _GEN_1108 : meta_79_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2133 = io_cpu_fence_value & _T & _T_2 ? _GEN_1109 : meta_80_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2134 = io_cpu_fence_value & _T & _T_2 ? _GEN_1110 : meta_81_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2135 = io_cpu_fence_value & _T & _T_2 ? _GEN_1111 : meta_82_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2136 = io_cpu_fence_value & _T & _T_2 ? _GEN_1112 : meta_83_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2137 = io_cpu_fence_value & _T & _T_2 ? _GEN_1113 : meta_84_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2138 = io_cpu_fence_value & _T & _T_2 ? _GEN_1114 : meta_85_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2139 = io_cpu_fence_value & _T & _T_2 ? _GEN_1115 : meta_86_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2140 = io_cpu_fence_value & _T & _T_2 ? _GEN_1116 : meta_87_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2141 = io_cpu_fence_value & _T & _T_2 ? _GEN_1117 : meta_88_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2142 = io_cpu_fence_value & _T & _T_2 ? _GEN_1118 : meta_89_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2143 = io_cpu_fence_value & _T & _T_2 ? _GEN_1119 : meta_90_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2144 = io_cpu_fence_value & _T & _T_2 ? _GEN_1120 : meta_91_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2145 = io_cpu_fence_value & _T & _T_2 ? _GEN_1121 : meta_92_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2146 = io_cpu_fence_value & _T & _T_2 ? _GEN_1122 : meta_93_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2147 = io_cpu_fence_value & _T & _T_2 ? _GEN_1123 : meta_94_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2148 = io_cpu_fence_value & _T & _T_2 ? _GEN_1124 : meta_95_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2149 = io_cpu_fence_value & _T & _T_2 ? _GEN_1125 : meta_96_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2150 = io_cpu_fence_value & _T & _T_2 ? _GEN_1126 : meta_97_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2151 = io_cpu_fence_value & _T & _T_2 ? _GEN_1127 : meta_98_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2152 = io_cpu_fence_value & _T & _T_2 ? _GEN_1128 : meta_99_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2153 = io_cpu_fence_value & _T & _T_2 ? _GEN_1129 : meta_100_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2154 = io_cpu_fence_value & _T & _T_2 ? _GEN_1130 : meta_101_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2155 = io_cpu_fence_value & _T & _T_2 ? _GEN_1131 : meta_102_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2156 = io_cpu_fence_value & _T & _T_2 ? _GEN_1132 : meta_103_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2157 = io_cpu_fence_value & _T & _T_2 ? _GEN_1133 : meta_104_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2158 = io_cpu_fence_value & _T & _T_2 ? _GEN_1134 : meta_105_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2159 = io_cpu_fence_value & _T & _T_2 ? _GEN_1135 : meta_106_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2160 = io_cpu_fence_value & _T & _T_2 ? _GEN_1136 : meta_107_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2161 = io_cpu_fence_value & _T & _T_2 ? _GEN_1137 : meta_108_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2162 = io_cpu_fence_value & _T & _T_2 ? _GEN_1138 : meta_109_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2163 = io_cpu_fence_value & _T & _T_2 ? _GEN_1139 : meta_110_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2164 = io_cpu_fence_value & _T & _T_2 ? _GEN_1140 : meta_111_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2165 = io_cpu_fence_value & _T & _T_2 ? _GEN_1141 : meta_112_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2166 = io_cpu_fence_value & _T & _T_2 ? _GEN_1142 : meta_113_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2167 = io_cpu_fence_value & _T & _T_2 ? _GEN_1143 : meta_114_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2168 = io_cpu_fence_value & _T & _T_2 ? _GEN_1144 : meta_115_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2169 = io_cpu_fence_value & _T & _T_2 ? _GEN_1145 : meta_116_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2170 = io_cpu_fence_value & _T & _T_2 ? _GEN_1146 : meta_117_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2171 = io_cpu_fence_value & _T & _T_2 ? _GEN_1147 : meta_118_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2172 = io_cpu_fence_value & _T & _T_2 ? _GEN_1148 : meta_119_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2173 = io_cpu_fence_value & _T & _T_2 ? _GEN_1149 : meta_120_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2174 = io_cpu_fence_value & _T & _T_2 ? _GEN_1150 : meta_121_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2175 = io_cpu_fence_value & _T & _T_2 ? _GEN_1151 : meta_122_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2176 = io_cpu_fence_value & _T & _T_2 ? _GEN_1152 : meta_123_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2177 = io_cpu_fence_value & _T & _T_2 ? _GEN_1153 : meta_124_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2178 = io_cpu_fence_value & _T & _T_2 ? _GEN_1154 : meta_125_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2179 = io_cpu_fence_value & _T & _T_2 ? _GEN_1155 : meta_126_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2180 = io_cpu_fence_value & _T & _T_2 ? _GEN_1156 : meta_127_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2181 = io_cpu_fence_value & _T & _T_2 ? _GEN_1157 : meta_128_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2182 = io_cpu_fence_value & _T & _T_2 ? _GEN_1158 : meta_129_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2183 = io_cpu_fence_value & _T & _T_2 ? _GEN_1159 : meta_130_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2184 = io_cpu_fence_value & _T & _T_2 ? _GEN_1160 : meta_131_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2185 = io_cpu_fence_value & _T & _T_2 ? _GEN_1161 : meta_132_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2186 = io_cpu_fence_value & _T & _T_2 ? _GEN_1162 : meta_133_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2187 = io_cpu_fence_value & _T & _T_2 ? _GEN_1163 : meta_134_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2188 = io_cpu_fence_value & _T & _T_2 ? _GEN_1164 : meta_135_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2189 = io_cpu_fence_value & _T & _T_2 ? _GEN_1165 : meta_136_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2190 = io_cpu_fence_value & _T & _T_2 ? _GEN_1166 : meta_137_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2191 = io_cpu_fence_value & _T & _T_2 ? _GEN_1167 : meta_138_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2192 = io_cpu_fence_value & _T & _T_2 ? _GEN_1168 : meta_139_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2193 = io_cpu_fence_value & _T & _T_2 ? _GEN_1169 : meta_140_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2194 = io_cpu_fence_value & _T & _T_2 ? _GEN_1170 : meta_141_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2195 = io_cpu_fence_value & _T & _T_2 ? _GEN_1171 : meta_142_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2196 = io_cpu_fence_value & _T & _T_2 ? _GEN_1172 : meta_143_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2197 = io_cpu_fence_value & _T & _T_2 ? _GEN_1173 : meta_144_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2198 = io_cpu_fence_value & _T & _T_2 ? _GEN_1174 : meta_145_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2199 = io_cpu_fence_value & _T & _T_2 ? _GEN_1175 : meta_146_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2200 = io_cpu_fence_value & _T & _T_2 ? _GEN_1176 : meta_147_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2201 = io_cpu_fence_value & _T & _T_2 ? _GEN_1177 : meta_148_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2202 = io_cpu_fence_value & _T & _T_2 ? _GEN_1178 : meta_149_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2203 = io_cpu_fence_value & _T & _T_2 ? _GEN_1179 : meta_150_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2204 = io_cpu_fence_value & _T & _T_2 ? _GEN_1180 : meta_151_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2205 = io_cpu_fence_value & _T & _T_2 ? _GEN_1181 : meta_152_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2206 = io_cpu_fence_value & _T & _T_2 ? _GEN_1182 : meta_153_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2207 = io_cpu_fence_value & _T & _T_2 ? _GEN_1183 : meta_154_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2208 = io_cpu_fence_value & _T & _T_2 ? _GEN_1184 : meta_155_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2209 = io_cpu_fence_value & _T & _T_2 ? _GEN_1185 : meta_156_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2210 = io_cpu_fence_value & _T & _T_2 ? _GEN_1186 : meta_157_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2211 = io_cpu_fence_value & _T & _T_2 ? _GEN_1187 : meta_158_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2212 = io_cpu_fence_value & _T & _T_2 ? _GEN_1188 : meta_159_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2213 = io_cpu_fence_value & _T & _T_2 ? _GEN_1189 : meta_160_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2214 = io_cpu_fence_value & _T & _T_2 ? _GEN_1190 : meta_161_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2215 = io_cpu_fence_value & _T & _T_2 ? _GEN_1191 : meta_162_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2216 = io_cpu_fence_value & _T & _T_2 ? _GEN_1192 : meta_163_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2217 = io_cpu_fence_value & _T & _T_2 ? _GEN_1193 : meta_164_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2218 = io_cpu_fence_value & _T & _T_2 ? _GEN_1194 : meta_165_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2219 = io_cpu_fence_value & _T & _T_2 ? _GEN_1195 : meta_166_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2220 = io_cpu_fence_value & _T & _T_2 ? _GEN_1196 : meta_167_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2221 = io_cpu_fence_value & _T & _T_2 ? _GEN_1197 : meta_168_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2222 = io_cpu_fence_value & _T & _T_2 ? _GEN_1198 : meta_169_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2223 = io_cpu_fence_value & _T & _T_2 ? _GEN_1199 : meta_170_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2224 = io_cpu_fence_value & _T & _T_2 ? _GEN_1200 : meta_171_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2225 = io_cpu_fence_value & _T & _T_2 ? _GEN_1201 : meta_172_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2226 = io_cpu_fence_value & _T & _T_2 ? _GEN_1202 : meta_173_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2227 = io_cpu_fence_value & _T & _T_2 ? _GEN_1203 : meta_174_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2228 = io_cpu_fence_value & _T & _T_2 ? _GEN_1204 : meta_175_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2229 = io_cpu_fence_value & _T & _T_2 ? _GEN_1205 : meta_176_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2230 = io_cpu_fence_value & _T & _T_2 ? _GEN_1206 : meta_177_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2231 = io_cpu_fence_value & _T & _T_2 ? _GEN_1207 : meta_178_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2232 = io_cpu_fence_value & _T & _T_2 ? _GEN_1208 : meta_179_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2233 = io_cpu_fence_value & _T & _T_2 ? _GEN_1209 : meta_180_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2234 = io_cpu_fence_value & _T & _T_2 ? _GEN_1210 : meta_181_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2235 = io_cpu_fence_value & _T & _T_2 ? _GEN_1211 : meta_182_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2236 = io_cpu_fence_value & _T & _T_2 ? _GEN_1212 : meta_183_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2237 = io_cpu_fence_value & _T & _T_2 ? _GEN_1213 : meta_184_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2238 = io_cpu_fence_value & _T & _T_2 ? _GEN_1214 : meta_185_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2239 = io_cpu_fence_value & _T & _T_2 ? _GEN_1215 : meta_186_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2240 = io_cpu_fence_value & _T & _T_2 ? _GEN_1216 : meta_187_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2241 = io_cpu_fence_value & _T & _T_2 ? _GEN_1217 : meta_188_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2242 = io_cpu_fence_value & _T & _T_2 ? _GEN_1218 : meta_189_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2243 = io_cpu_fence_value & _T & _T_2 ? _GEN_1219 : meta_190_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2244 = io_cpu_fence_value & _T & _T_2 ? _GEN_1220 : meta_191_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2245 = io_cpu_fence_value & _T & _T_2 ? _GEN_1221 : meta_192_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2246 = io_cpu_fence_value & _T & _T_2 ? _GEN_1222 : meta_193_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2247 = io_cpu_fence_value & _T & _T_2 ? _GEN_1223 : meta_194_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2248 = io_cpu_fence_value & _T & _T_2 ? _GEN_1224 : meta_195_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2249 = io_cpu_fence_value & _T & _T_2 ? _GEN_1225 : meta_196_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2250 = io_cpu_fence_value & _T & _T_2 ? _GEN_1226 : meta_197_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2251 = io_cpu_fence_value & _T & _T_2 ? _GEN_1227 : meta_198_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2252 = io_cpu_fence_value & _T & _T_2 ? _GEN_1228 : meta_199_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2253 = io_cpu_fence_value & _T & _T_2 ? _GEN_1229 : meta_200_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2254 = io_cpu_fence_value & _T & _T_2 ? _GEN_1230 : meta_201_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2255 = io_cpu_fence_value & _T & _T_2 ? _GEN_1231 : meta_202_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2256 = io_cpu_fence_value & _T & _T_2 ? _GEN_1232 : meta_203_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2257 = io_cpu_fence_value & _T & _T_2 ? _GEN_1233 : meta_204_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2258 = io_cpu_fence_value & _T & _T_2 ? _GEN_1234 : meta_205_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2259 = io_cpu_fence_value & _T & _T_2 ? _GEN_1235 : meta_206_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2260 = io_cpu_fence_value & _T & _T_2 ? _GEN_1236 : meta_207_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2261 = io_cpu_fence_value & _T & _T_2 ? _GEN_1237 : meta_208_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2262 = io_cpu_fence_value & _T & _T_2 ? _GEN_1238 : meta_209_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2263 = io_cpu_fence_value & _T & _T_2 ? _GEN_1239 : meta_210_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2264 = io_cpu_fence_value & _T & _T_2 ? _GEN_1240 : meta_211_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2265 = io_cpu_fence_value & _T & _T_2 ? _GEN_1241 : meta_212_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2266 = io_cpu_fence_value & _T & _T_2 ? _GEN_1242 : meta_213_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2267 = io_cpu_fence_value & _T & _T_2 ? _GEN_1243 : meta_214_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2268 = io_cpu_fence_value & _T & _T_2 ? _GEN_1244 : meta_215_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2269 = io_cpu_fence_value & _T & _T_2 ? _GEN_1245 : meta_216_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2270 = io_cpu_fence_value & _T & _T_2 ? _GEN_1246 : meta_217_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2271 = io_cpu_fence_value & _T & _T_2 ? _GEN_1247 : meta_218_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2272 = io_cpu_fence_value & _T & _T_2 ? _GEN_1248 : meta_219_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2273 = io_cpu_fence_value & _T & _T_2 ? _GEN_1249 : meta_220_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2274 = io_cpu_fence_value & _T & _T_2 ? _GEN_1250 : meta_221_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2275 = io_cpu_fence_value & _T & _T_2 ? _GEN_1251 : meta_222_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2276 = io_cpu_fence_value & _T & _T_2 ? _GEN_1252 : meta_223_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2277 = io_cpu_fence_value & _T & _T_2 ? _GEN_1253 : meta_224_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2278 = io_cpu_fence_value & _T & _T_2 ? _GEN_1254 : meta_225_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2279 = io_cpu_fence_value & _T & _T_2 ? _GEN_1255 : meta_226_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2280 = io_cpu_fence_value & _T & _T_2 ? _GEN_1256 : meta_227_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2281 = io_cpu_fence_value & _T & _T_2 ? _GEN_1257 : meta_228_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2282 = io_cpu_fence_value & _T & _T_2 ? _GEN_1258 : meta_229_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2283 = io_cpu_fence_value & _T & _T_2 ? _GEN_1259 : meta_230_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2284 = io_cpu_fence_value & _T & _T_2 ? _GEN_1260 : meta_231_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2285 = io_cpu_fence_value & _T & _T_2 ? _GEN_1261 : meta_232_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2286 = io_cpu_fence_value & _T & _T_2 ? _GEN_1262 : meta_233_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2287 = io_cpu_fence_value & _T & _T_2 ? _GEN_1263 : meta_234_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2288 = io_cpu_fence_value & _T & _T_2 ? _GEN_1264 : meta_235_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2289 = io_cpu_fence_value & _T & _T_2 ? _GEN_1265 : meta_236_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2290 = io_cpu_fence_value & _T & _T_2 ? _GEN_1266 : meta_237_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2291 = io_cpu_fence_value & _T & _T_2 ? _GEN_1267 : meta_238_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2292 = io_cpu_fence_value & _T & _T_2 ? _GEN_1268 : meta_239_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2293 = io_cpu_fence_value & _T & _T_2 ? _GEN_1269 : meta_240_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2294 = io_cpu_fence_value & _T & _T_2 ? _GEN_1270 : meta_241_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2295 = io_cpu_fence_value & _T & _T_2 ? _GEN_1271 : meta_242_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2296 = io_cpu_fence_value & _T & _T_2 ? _GEN_1272 : meta_243_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2297 = io_cpu_fence_value & _T & _T_2 ? _GEN_1273 : meta_244_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2298 = io_cpu_fence_value & _T & _T_2 ? _GEN_1274 : meta_245_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2299 = io_cpu_fence_value & _T & _T_2 ? _GEN_1275 : meta_246_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2300 = io_cpu_fence_value & _T & _T_2 ? _GEN_1276 : meta_247_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2301 = io_cpu_fence_value & _T & _T_2 ? _GEN_1277 : meta_248_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2302 = io_cpu_fence_value & _T & _T_2 ? _GEN_1278 : meta_249_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2303 = io_cpu_fence_value & _T & _T_2 ? _GEN_1279 : meta_250_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2304 = io_cpu_fence_value & _T & _T_2 ? _GEN_1280 : meta_251_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2305 = io_cpu_fence_value & _T & _T_2 ? _GEN_1281 : meta_252_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2306 = io_cpu_fence_value & _T & _T_2 ? _GEN_1282 : meta_253_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2307 = io_cpu_fence_value & _T & _T_2 ? _GEN_1283 : meta_254_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2308 = io_cpu_fence_value & _T & _T_2 ? _GEN_1284 : meta_255_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2309 = io_cpu_fence_value & _T & _T_2 ? _GEN_1285 : meta_256_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2310 = io_cpu_fence_value & _T & _T_2 ? _GEN_1286 : meta_257_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2311 = io_cpu_fence_value & _T & _T_2 ? _GEN_1287 : meta_258_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2312 = io_cpu_fence_value & _T & _T_2 ? _GEN_1288 : meta_259_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2313 = io_cpu_fence_value & _T & _T_2 ? _GEN_1289 : meta_260_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2314 = io_cpu_fence_value & _T & _T_2 ? _GEN_1290 : meta_261_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2315 = io_cpu_fence_value & _T & _T_2 ? _GEN_1291 : meta_262_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2316 = io_cpu_fence_value & _T & _T_2 ? _GEN_1292 : meta_263_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2317 = io_cpu_fence_value & _T & _T_2 ? _GEN_1293 : meta_264_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2318 = io_cpu_fence_value & _T & _T_2 ? _GEN_1294 : meta_265_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2319 = io_cpu_fence_value & _T & _T_2 ? _GEN_1295 : meta_266_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2320 = io_cpu_fence_value & _T & _T_2 ? _GEN_1296 : meta_267_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2321 = io_cpu_fence_value & _T & _T_2 ? _GEN_1297 : meta_268_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2322 = io_cpu_fence_value & _T & _T_2 ? _GEN_1298 : meta_269_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2323 = io_cpu_fence_value & _T & _T_2 ? _GEN_1299 : meta_270_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2324 = io_cpu_fence_value & _T & _T_2 ? _GEN_1300 : meta_271_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2325 = io_cpu_fence_value & _T & _T_2 ? _GEN_1301 : meta_272_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2326 = io_cpu_fence_value & _T & _T_2 ? _GEN_1302 : meta_273_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2327 = io_cpu_fence_value & _T & _T_2 ? _GEN_1303 : meta_274_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2328 = io_cpu_fence_value & _T & _T_2 ? _GEN_1304 : meta_275_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2329 = io_cpu_fence_value & _T & _T_2 ? _GEN_1305 : meta_276_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2330 = io_cpu_fence_value & _T & _T_2 ? _GEN_1306 : meta_277_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2331 = io_cpu_fence_value & _T & _T_2 ? _GEN_1307 : meta_278_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2332 = io_cpu_fence_value & _T & _T_2 ? _GEN_1308 : meta_279_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2333 = io_cpu_fence_value & _T & _T_2 ? _GEN_1309 : meta_280_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2334 = io_cpu_fence_value & _T & _T_2 ? _GEN_1310 : meta_281_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2335 = io_cpu_fence_value & _T & _T_2 ? _GEN_1311 : meta_282_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2336 = io_cpu_fence_value & _T & _T_2 ? _GEN_1312 : meta_283_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2337 = io_cpu_fence_value & _T & _T_2 ? _GEN_1313 : meta_284_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2338 = io_cpu_fence_value & _T & _T_2 ? _GEN_1314 : meta_285_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2339 = io_cpu_fence_value & _T & _T_2 ? _GEN_1315 : meta_286_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2340 = io_cpu_fence_value & _T & _T_2 ? _GEN_1316 : meta_287_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2341 = io_cpu_fence_value & _T & _T_2 ? _GEN_1317 : meta_288_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2342 = io_cpu_fence_value & _T & _T_2 ? _GEN_1318 : meta_289_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2343 = io_cpu_fence_value & _T & _T_2 ? _GEN_1319 : meta_290_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2344 = io_cpu_fence_value & _T & _T_2 ? _GEN_1320 : meta_291_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2345 = io_cpu_fence_value & _T & _T_2 ? _GEN_1321 : meta_292_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2346 = io_cpu_fence_value & _T & _T_2 ? _GEN_1322 : meta_293_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2347 = io_cpu_fence_value & _T & _T_2 ? _GEN_1323 : meta_294_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2348 = io_cpu_fence_value & _T & _T_2 ? _GEN_1324 : meta_295_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2349 = io_cpu_fence_value & _T & _T_2 ? _GEN_1325 : meta_296_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2350 = io_cpu_fence_value & _T & _T_2 ? _GEN_1326 : meta_297_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2351 = io_cpu_fence_value & _T & _T_2 ? _GEN_1327 : meta_298_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2352 = io_cpu_fence_value & _T & _T_2 ? _GEN_1328 : meta_299_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2353 = io_cpu_fence_value & _T & _T_2 ? _GEN_1329 : meta_300_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2354 = io_cpu_fence_value & _T & _T_2 ? _GEN_1330 : meta_301_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2355 = io_cpu_fence_value & _T & _T_2 ? _GEN_1331 : meta_302_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2356 = io_cpu_fence_value & _T & _T_2 ? _GEN_1332 : meta_303_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2357 = io_cpu_fence_value & _T & _T_2 ? _GEN_1333 : meta_304_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2358 = io_cpu_fence_value & _T & _T_2 ? _GEN_1334 : meta_305_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2359 = io_cpu_fence_value & _T & _T_2 ? _GEN_1335 : meta_306_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2360 = io_cpu_fence_value & _T & _T_2 ? _GEN_1336 : meta_307_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2361 = io_cpu_fence_value & _T & _T_2 ? _GEN_1337 : meta_308_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2362 = io_cpu_fence_value & _T & _T_2 ? _GEN_1338 : meta_309_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2363 = io_cpu_fence_value & _T & _T_2 ? _GEN_1339 : meta_310_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2364 = io_cpu_fence_value & _T & _T_2 ? _GEN_1340 : meta_311_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2365 = io_cpu_fence_value & _T & _T_2 ? _GEN_1341 : meta_312_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2366 = io_cpu_fence_value & _T & _T_2 ? _GEN_1342 : meta_313_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2367 = io_cpu_fence_value & _T & _T_2 ? _GEN_1343 : meta_314_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2368 = io_cpu_fence_value & _T & _T_2 ? _GEN_1344 : meta_315_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2369 = io_cpu_fence_value & _T & _T_2 ? _GEN_1345 : meta_316_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2370 = io_cpu_fence_value & _T & _T_2 ? _GEN_1346 : meta_317_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2371 = io_cpu_fence_value & _T & _T_2 ? _GEN_1347 : meta_318_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2372 = io_cpu_fence_value & _T & _T_2 ? _GEN_1348 : meta_319_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2373 = io_cpu_fence_value & _T & _T_2 ? _GEN_1349 : meta_320_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2374 = io_cpu_fence_value & _T & _T_2 ? _GEN_1350 : meta_321_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2375 = io_cpu_fence_value & _T & _T_2 ? _GEN_1351 : meta_322_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2376 = io_cpu_fence_value & _T & _T_2 ? _GEN_1352 : meta_323_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2377 = io_cpu_fence_value & _T & _T_2 ? _GEN_1353 : meta_324_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2378 = io_cpu_fence_value & _T & _T_2 ? _GEN_1354 : meta_325_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2379 = io_cpu_fence_value & _T & _T_2 ? _GEN_1355 : meta_326_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2380 = io_cpu_fence_value & _T & _T_2 ? _GEN_1356 : meta_327_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2381 = io_cpu_fence_value & _T & _T_2 ? _GEN_1357 : meta_328_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2382 = io_cpu_fence_value & _T & _T_2 ? _GEN_1358 : meta_329_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2383 = io_cpu_fence_value & _T & _T_2 ? _GEN_1359 : meta_330_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2384 = io_cpu_fence_value & _T & _T_2 ? _GEN_1360 : meta_331_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2385 = io_cpu_fence_value & _T & _T_2 ? _GEN_1361 : meta_332_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2386 = io_cpu_fence_value & _T & _T_2 ? _GEN_1362 : meta_333_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2387 = io_cpu_fence_value & _T & _T_2 ? _GEN_1363 : meta_334_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2388 = io_cpu_fence_value & _T & _T_2 ? _GEN_1364 : meta_335_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2389 = io_cpu_fence_value & _T & _T_2 ? _GEN_1365 : meta_336_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2390 = io_cpu_fence_value & _T & _T_2 ? _GEN_1366 : meta_337_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2391 = io_cpu_fence_value & _T & _T_2 ? _GEN_1367 : meta_338_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2392 = io_cpu_fence_value & _T & _T_2 ? _GEN_1368 : meta_339_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2393 = io_cpu_fence_value & _T & _T_2 ? _GEN_1369 : meta_340_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2394 = io_cpu_fence_value & _T & _T_2 ? _GEN_1370 : meta_341_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2395 = io_cpu_fence_value & _T & _T_2 ? _GEN_1371 : meta_342_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2396 = io_cpu_fence_value & _T & _T_2 ? _GEN_1372 : meta_343_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2397 = io_cpu_fence_value & _T & _T_2 ? _GEN_1373 : meta_344_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2398 = io_cpu_fence_value & _T & _T_2 ? _GEN_1374 : meta_345_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2399 = io_cpu_fence_value & _T & _T_2 ? _GEN_1375 : meta_346_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2400 = io_cpu_fence_value & _T & _T_2 ? _GEN_1376 : meta_347_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2401 = io_cpu_fence_value & _T & _T_2 ? _GEN_1377 : meta_348_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2402 = io_cpu_fence_value & _T & _T_2 ? _GEN_1378 : meta_349_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2403 = io_cpu_fence_value & _T & _T_2 ? _GEN_1379 : meta_350_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2404 = io_cpu_fence_value & _T & _T_2 ? _GEN_1380 : meta_351_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2405 = io_cpu_fence_value & _T & _T_2 ? _GEN_1381 : meta_352_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2406 = io_cpu_fence_value & _T & _T_2 ? _GEN_1382 : meta_353_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2407 = io_cpu_fence_value & _T & _T_2 ? _GEN_1383 : meta_354_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2408 = io_cpu_fence_value & _T & _T_2 ? _GEN_1384 : meta_355_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2409 = io_cpu_fence_value & _T & _T_2 ? _GEN_1385 : meta_356_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2410 = io_cpu_fence_value & _T & _T_2 ? _GEN_1386 : meta_357_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2411 = io_cpu_fence_value & _T & _T_2 ? _GEN_1387 : meta_358_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2412 = io_cpu_fence_value & _T & _T_2 ? _GEN_1388 : meta_359_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2413 = io_cpu_fence_value & _T & _T_2 ? _GEN_1389 : meta_360_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2414 = io_cpu_fence_value & _T & _T_2 ? _GEN_1390 : meta_361_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2415 = io_cpu_fence_value & _T & _T_2 ? _GEN_1391 : meta_362_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2416 = io_cpu_fence_value & _T & _T_2 ? _GEN_1392 : meta_363_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2417 = io_cpu_fence_value & _T & _T_2 ? _GEN_1393 : meta_364_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2418 = io_cpu_fence_value & _T & _T_2 ? _GEN_1394 : meta_365_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2419 = io_cpu_fence_value & _T & _T_2 ? _GEN_1395 : meta_366_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2420 = io_cpu_fence_value & _T & _T_2 ? _GEN_1396 : meta_367_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2421 = io_cpu_fence_value & _T & _T_2 ? _GEN_1397 : meta_368_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2422 = io_cpu_fence_value & _T & _T_2 ? _GEN_1398 : meta_369_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2423 = io_cpu_fence_value & _T & _T_2 ? _GEN_1399 : meta_370_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2424 = io_cpu_fence_value & _T & _T_2 ? _GEN_1400 : meta_371_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2425 = io_cpu_fence_value & _T & _T_2 ? _GEN_1401 : meta_372_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2426 = io_cpu_fence_value & _T & _T_2 ? _GEN_1402 : meta_373_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2427 = io_cpu_fence_value & _T & _T_2 ? _GEN_1403 : meta_374_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2428 = io_cpu_fence_value & _T & _T_2 ? _GEN_1404 : meta_375_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2429 = io_cpu_fence_value & _T & _T_2 ? _GEN_1405 : meta_376_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2430 = io_cpu_fence_value & _T & _T_2 ? _GEN_1406 : meta_377_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2431 = io_cpu_fence_value & _T & _T_2 ? _GEN_1407 : meta_378_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2432 = io_cpu_fence_value & _T & _T_2 ? _GEN_1408 : meta_379_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2433 = io_cpu_fence_value & _T & _T_2 ? _GEN_1409 : meta_380_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2434 = io_cpu_fence_value & _T & _T_2 ? _GEN_1410 : meta_381_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2435 = io_cpu_fence_value & _T & _T_2 ? _GEN_1411 : meta_382_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2436 = io_cpu_fence_value & _T & _T_2 ? _GEN_1412 : meta_383_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2437 = io_cpu_fence_value & _T & _T_2 ? _GEN_1413 : meta_384_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2438 = io_cpu_fence_value & _T & _T_2 ? _GEN_1414 : meta_385_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2439 = io_cpu_fence_value & _T & _T_2 ? _GEN_1415 : meta_386_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2440 = io_cpu_fence_value & _T & _T_2 ? _GEN_1416 : meta_387_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2441 = io_cpu_fence_value & _T & _T_2 ? _GEN_1417 : meta_388_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2442 = io_cpu_fence_value & _T & _T_2 ? _GEN_1418 : meta_389_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2443 = io_cpu_fence_value & _T & _T_2 ? _GEN_1419 : meta_390_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2444 = io_cpu_fence_value & _T & _T_2 ? _GEN_1420 : meta_391_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2445 = io_cpu_fence_value & _T & _T_2 ? _GEN_1421 : meta_392_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2446 = io_cpu_fence_value & _T & _T_2 ? _GEN_1422 : meta_393_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2447 = io_cpu_fence_value & _T & _T_2 ? _GEN_1423 : meta_394_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2448 = io_cpu_fence_value & _T & _T_2 ? _GEN_1424 : meta_395_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2449 = io_cpu_fence_value & _T & _T_2 ? _GEN_1425 : meta_396_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2450 = io_cpu_fence_value & _T & _T_2 ? _GEN_1426 : meta_397_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2451 = io_cpu_fence_value & _T & _T_2 ? _GEN_1427 : meta_398_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2452 = io_cpu_fence_value & _T & _T_2 ? _GEN_1428 : meta_399_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2453 = io_cpu_fence_value & _T & _T_2 ? _GEN_1429 : meta_400_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2454 = io_cpu_fence_value & _T & _T_2 ? _GEN_1430 : meta_401_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2455 = io_cpu_fence_value & _T & _T_2 ? _GEN_1431 : meta_402_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2456 = io_cpu_fence_value & _T & _T_2 ? _GEN_1432 : meta_403_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2457 = io_cpu_fence_value & _T & _T_2 ? _GEN_1433 : meta_404_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2458 = io_cpu_fence_value & _T & _T_2 ? _GEN_1434 : meta_405_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2459 = io_cpu_fence_value & _T & _T_2 ? _GEN_1435 : meta_406_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2460 = io_cpu_fence_value & _T & _T_2 ? _GEN_1436 : meta_407_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2461 = io_cpu_fence_value & _T & _T_2 ? _GEN_1437 : meta_408_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2462 = io_cpu_fence_value & _T & _T_2 ? _GEN_1438 : meta_409_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2463 = io_cpu_fence_value & _T & _T_2 ? _GEN_1439 : meta_410_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2464 = io_cpu_fence_value & _T & _T_2 ? _GEN_1440 : meta_411_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2465 = io_cpu_fence_value & _T & _T_2 ? _GEN_1441 : meta_412_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2466 = io_cpu_fence_value & _T & _T_2 ? _GEN_1442 : meta_413_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2467 = io_cpu_fence_value & _T & _T_2 ? _GEN_1443 : meta_414_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2468 = io_cpu_fence_value & _T & _T_2 ? _GEN_1444 : meta_415_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2469 = io_cpu_fence_value & _T & _T_2 ? _GEN_1445 : meta_416_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2470 = io_cpu_fence_value & _T & _T_2 ? _GEN_1446 : meta_417_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2471 = io_cpu_fence_value & _T & _T_2 ? _GEN_1447 : meta_418_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2472 = io_cpu_fence_value & _T & _T_2 ? _GEN_1448 : meta_419_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2473 = io_cpu_fence_value & _T & _T_2 ? _GEN_1449 : meta_420_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2474 = io_cpu_fence_value & _T & _T_2 ? _GEN_1450 : meta_421_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2475 = io_cpu_fence_value & _T & _T_2 ? _GEN_1451 : meta_422_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2476 = io_cpu_fence_value & _T & _T_2 ? _GEN_1452 : meta_423_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2477 = io_cpu_fence_value & _T & _T_2 ? _GEN_1453 : meta_424_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2478 = io_cpu_fence_value & _T & _T_2 ? _GEN_1454 : meta_425_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2479 = io_cpu_fence_value & _T & _T_2 ? _GEN_1455 : meta_426_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2480 = io_cpu_fence_value & _T & _T_2 ? _GEN_1456 : meta_427_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2481 = io_cpu_fence_value & _T & _T_2 ? _GEN_1457 : meta_428_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2482 = io_cpu_fence_value & _T & _T_2 ? _GEN_1458 : meta_429_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2483 = io_cpu_fence_value & _T & _T_2 ? _GEN_1459 : meta_430_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2484 = io_cpu_fence_value & _T & _T_2 ? _GEN_1460 : meta_431_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2485 = io_cpu_fence_value & _T & _T_2 ? _GEN_1461 : meta_432_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2486 = io_cpu_fence_value & _T & _T_2 ? _GEN_1462 : meta_433_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2487 = io_cpu_fence_value & _T & _T_2 ? _GEN_1463 : meta_434_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2488 = io_cpu_fence_value & _T & _T_2 ? _GEN_1464 : meta_435_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2489 = io_cpu_fence_value & _T & _T_2 ? _GEN_1465 : meta_436_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2490 = io_cpu_fence_value & _T & _T_2 ? _GEN_1466 : meta_437_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2491 = io_cpu_fence_value & _T & _T_2 ? _GEN_1467 : meta_438_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2492 = io_cpu_fence_value & _T & _T_2 ? _GEN_1468 : meta_439_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2493 = io_cpu_fence_value & _T & _T_2 ? _GEN_1469 : meta_440_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2494 = io_cpu_fence_value & _T & _T_2 ? _GEN_1470 : meta_441_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2495 = io_cpu_fence_value & _T & _T_2 ? _GEN_1471 : meta_442_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2496 = io_cpu_fence_value & _T & _T_2 ? _GEN_1472 : meta_443_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2497 = io_cpu_fence_value & _T & _T_2 ? _GEN_1473 : meta_444_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2498 = io_cpu_fence_value & _T & _T_2 ? _GEN_1474 : meta_445_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2499 = io_cpu_fence_value & _T & _T_2 ? _GEN_1475 : meta_446_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2500 = io_cpu_fence_value & _T & _T_2 ? _GEN_1476 : meta_447_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2501 = io_cpu_fence_value & _T & _T_2 ? _GEN_1477 : meta_448_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2502 = io_cpu_fence_value & _T & _T_2 ? _GEN_1478 : meta_449_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2503 = io_cpu_fence_value & _T & _T_2 ? _GEN_1479 : meta_450_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2504 = io_cpu_fence_value & _T & _T_2 ? _GEN_1480 : meta_451_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2505 = io_cpu_fence_value & _T & _T_2 ? _GEN_1481 : meta_452_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2506 = io_cpu_fence_value & _T & _T_2 ? _GEN_1482 : meta_453_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2507 = io_cpu_fence_value & _T & _T_2 ? _GEN_1483 : meta_454_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2508 = io_cpu_fence_value & _T & _T_2 ? _GEN_1484 : meta_455_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2509 = io_cpu_fence_value & _T & _T_2 ? _GEN_1485 : meta_456_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2510 = io_cpu_fence_value & _T & _T_2 ? _GEN_1486 : meta_457_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2511 = io_cpu_fence_value & _T & _T_2 ? _GEN_1487 : meta_458_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2512 = io_cpu_fence_value & _T & _T_2 ? _GEN_1488 : meta_459_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2513 = io_cpu_fence_value & _T & _T_2 ? _GEN_1489 : meta_460_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2514 = io_cpu_fence_value & _T & _T_2 ? _GEN_1490 : meta_461_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2515 = io_cpu_fence_value & _T & _T_2 ? _GEN_1491 : meta_462_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2516 = io_cpu_fence_value & _T & _T_2 ? _GEN_1492 : meta_463_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2517 = io_cpu_fence_value & _T & _T_2 ? _GEN_1493 : meta_464_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2518 = io_cpu_fence_value & _T & _T_2 ? _GEN_1494 : meta_465_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2519 = io_cpu_fence_value & _T & _T_2 ? _GEN_1495 : meta_466_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2520 = io_cpu_fence_value & _T & _T_2 ? _GEN_1496 : meta_467_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2521 = io_cpu_fence_value & _T & _T_2 ? _GEN_1497 : meta_468_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2522 = io_cpu_fence_value & _T & _T_2 ? _GEN_1498 : meta_469_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2523 = io_cpu_fence_value & _T & _T_2 ? _GEN_1499 : meta_470_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2524 = io_cpu_fence_value & _T & _T_2 ? _GEN_1500 : meta_471_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2525 = io_cpu_fence_value & _T & _T_2 ? _GEN_1501 : meta_472_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2526 = io_cpu_fence_value & _T & _T_2 ? _GEN_1502 : meta_473_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2527 = io_cpu_fence_value & _T & _T_2 ? _GEN_1503 : meta_474_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2528 = io_cpu_fence_value & _T & _T_2 ? _GEN_1504 : meta_475_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2529 = io_cpu_fence_value & _T & _T_2 ? _GEN_1505 : meta_476_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2530 = io_cpu_fence_value & _T & _T_2 ? _GEN_1506 : meta_477_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2531 = io_cpu_fence_value & _T & _T_2 ? _GEN_1507 : meta_478_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2532 = io_cpu_fence_value & _T & _T_2 ? _GEN_1508 : meta_479_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2533 = io_cpu_fence_value & _T & _T_2 ? _GEN_1509 : meta_480_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2534 = io_cpu_fence_value & _T & _T_2 ? _GEN_1510 : meta_481_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2535 = io_cpu_fence_value & _T & _T_2 ? _GEN_1511 : meta_482_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2536 = io_cpu_fence_value & _T & _T_2 ? _GEN_1512 : meta_483_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2537 = io_cpu_fence_value & _T & _T_2 ? _GEN_1513 : meta_484_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2538 = io_cpu_fence_value & _T & _T_2 ? _GEN_1514 : meta_485_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2539 = io_cpu_fence_value & _T & _T_2 ? _GEN_1515 : meta_486_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2540 = io_cpu_fence_value & _T & _T_2 ? _GEN_1516 : meta_487_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2541 = io_cpu_fence_value & _T & _T_2 ? _GEN_1517 : meta_488_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2542 = io_cpu_fence_value & _T & _T_2 ? _GEN_1518 : meta_489_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2543 = io_cpu_fence_value & _T & _T_2 ? _GEN_1519 : meta_490_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2544 = io_cpu_fence_value & _T & _T_2 ? _GEN_1520 : meta_491_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2545 = io_cpu_fence_value & _T & _T_2 ? _GEN_1521 : meta_492_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2546 = io_cpu_fence_value & _T & _T_2 ? _GEN_1522 : meta_493_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2547 = io_cpu_fence_value & _T & _T_2 ? _GEN_1523 : meta_494_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2548 = io_cpu_fence_value & _T & _T_2 ? _GEN_1524 : meta_495_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2549 = io_cpu_fence_value & _T & _T_2 ? _GEN_1525 : meta_496_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2550 = io_cpu_fence_value & _T & _T_2 ? _GEN_1526 : meta_497_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2551 = io_cpu_fence_value & _T & _T_2 ? _GEN_1527 : meta_498_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2552 = io_cpu_fence_value & _T & _T_2 ? _GEN_1528 : meta_499_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2553 = io_cpu_fence_value & _T & _T_2 ? _GEN_1529 : meta_500_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2554 = io_cpu_fence_value & _T & _T_2 ? _GEN_1530 : meta_501_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2555 = io_cpu_fence_value & _T & _T_2 ? _GEN_1531 : meta_502_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2556 = io_cpu_fence_value & _T & _T_2 ? _GEN_1532 : meta_503_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2557 = io_cpu_fence_value & _T & _T_2 ? _GEN_1533 : meta_504_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2558 = io_cpu_fence_value & _T & _T_2 ? _GEN_1534 : meta_505_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2559 = io_cpu_fence_value & _T & _T_2 ? _GEN_1535 : meta_506_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2560 = io_cpu_fence_value & _T & _T_2 ? _GEN_1536 : meta_507_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2561 = io_cpu_fence_value & _T & _T_2 ? _GEN_1537 : meta_508_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2562 = io_cpu_fence_value & _T & _T_2 ? _GEN_1538 : meta_509_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2563 = io_cpu_fence_value & _T & _T_2 ? _GEN_1539 : meta_510_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2564 = io_cpu_fence_value & _T & _T_2 ? _GEN_1540 : meta_511_valid_0; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2565 = io_cpu_fence_value & _T & _T_2 ? _GEN_1541 : meta_0_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2566 = io_cpu_fence_value & _T & _T_2 ? _GEN_1542 : meta_1_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2567 = io_cpu_fence_value & _T & _T_2 ? _GEN_1543 : meta_2_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2568 = io_cpu_fence_value & _T & _T_2 ? _GEN_1544 : meta_3_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2569 = io_cpu_fence_value & _T & _T_2 ? _GEN_1545 : meta_4_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2570 = io_cpu_fence_value & _T & _T_2 ? _GEN_1546 : meta_5_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2571 = io_cpu_fence_value & _T & _T_2 ? _GEN_1547 : meta_6_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2572 = io_cpu_fence_value & _T & _T_2 ? _GEN_1548 : meta_7_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2573 = io_cpu_fence_value & _T & _T_2 ? _GEN_1549 : meta_8_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2574 = io_cpu_fence_value & _T & _T_2 ? _GEN_1550 : meta_9_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2575 = io_cpu_fence_value & _T & _T_2 ? _GEN_1551 : meta_10_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2576 = io_cpu_fence_value & _T & _T_2 ? _GEN_1552 : meta_11_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2577 = io_cpu_fence_value & _T & _T_2 ? _GEN_1553 : meta_12_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2578 = io_cpu_fence_value & _T & _T_2 ? _GEN_1554 : meta_13_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2579 = io_cpu_fence_value & _T & _T_2 ? _GEN_1555 : meta_14_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2580 = io_cpu_fence_value & _T & _T_2 ? _GEN_1556 : meta_15_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2581 = io_cpu_fence_value & _T & _T_2 ? _GEN_1557 : meta_16_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2582 = io_cpu_fence_value & _T & _T_2 ? _GEN_1558 : meta_17_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2583 = io_cpu_fence_value & _T & _T_2 ? _GEN_1559 : meta_18_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2584 = io_cpu_fence_value & _T & _T_2 ? _GEN_1560 : meta_19_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2585 = io_cpu_fence_value & _T & _T_2 ? _GEN_1561 : meta_20_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2586 = io_cpu_fence_value & _T & _T_2 ? _GEN_1562 : meta_21_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2587 = io_cpu_fence_value & _T & _T_2 ? _GEN_1563 : meta_22_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2588 = io_cpu_fence_value & _T & _T_2 ? _GEN_1564 : meta_23_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2589 = io_cpu_fence_value & _T & _T_2 ? _GEN_1565 : meta_24_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2590 = io_cpu_fence_value & _T & _T_2 ? _GEN_1566 : meta_25_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2591 = io_cpu_fence_value & _T & _T_2 ? _GEN_1567 : meta_26_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2592 = io_cpu_fence_value & _T & _T_2 ? _GEN_1568 : meta_27_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2593 = io_cpu_fence_value & _T & _T_2 ? _GEN_1569 : meta_28_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2594 = io_cpu_fence_value & _T & _T_2 ? _GEN_1570 : meta_29_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2595 = io_cpu_fence_value & _T & _T_2 ? _GEN_1571 : meta_30_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2596 = io_cpu_fence_value & _T & _T_2 ? _GEN_1572 : meta_31_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2597 = io_cpu_fence_value & _T & _T_2 ? _GEN_1573 : meta_32_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2598 = io_cpu_fence_value & _T & _T_2 ? _GEN_1574 : meta_33_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2599 = io_cpu_fence_value & _T & _T_2 ? _GEN_1575 : meta_34_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2600 = io_cpu_fence_value & _T & _T_2 ? _GEN_1576 : meta_35_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2601 = io_cpu_fence_value & _T & _T_2 ? _GEN_1577 : meta_36_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2602 = io_cpu_fence_value & _T & _T_2 ? _GEN_1578 : meta_37_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2603 = io_cpu_fence_value & _T & _T_2 ? _GEN_1579 : meta_38_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2604 = io_cpu_fence_value & _T & _T_2 ? _GEN_1580 : meta_39_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2605 = io_cpu_fence_value & _T & _T_2 ? _GEN_1581 : meta_40_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2606 = io_cpu_fence_value & _T & _T_2 ? _GEN_1582 : meta_41_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2607 = io_cpu_fence_value & _T & _T_2 ? _GEN_1583 : meta_42_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2608 = io_cpu_fence_value & _T & _T_2 ? _GEN_1584 : meta_43_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2609 = io_cpu_fence_value & _T & _T_2 ? _GEN_1585 : meta_44_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2610 = io_cpu_fence_value & _T & _T_2 ? _GEN_1586 : meta_45_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2611 = io_cpu_fence_value & _T & _T_2 ? _GEN_1587 : meta_46_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2612 = io_cpu_fence_value & _T & _T_2 ? _GEN_1588 : meta_47_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2613 = io_cpu_fence_value & _T & _T_2 ? _GEN_1589 : meta_48_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2614 = io_cpu_fence_value & _T & _T_2 ? _GEN_1590 : meta_49_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2615 = io_cpu_fence_value & _T & _T_2 ? _GEN_1591 : meta_50_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2616 = io_cpu_fence_value & _T & _T_2 ? _GEN_1592 : meta_51_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2617 = io_cpu_fence_value & _T & _T_2 ? _GEN_1593 : meta_52_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2618 = io_cpu_fence_value & _T & _T_2 ? _GEN_1594 : meta_53_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2619 = io_cpu_fence_value & _T & _T_2 ? _GEN_1595 : meta_54_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2620 = io_cpu_fence_value & _T & _T_2 ? _GEN_1596 : meta_55_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2621 = io_cpu_fence_value & _T & _T_2 ? _GEN_1597 : meta_56_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2622 = io_cpu_fence_value & _T & _T_2 ? _GEN_1598 : meta_57_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2623 = io_cpu_fence_value & _T & _T_2 ? _GEN_1599 : meta_58_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2624 = io_cpu_fence_value & _T & _T_2 ? _GEN_1600 : meta_59_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2625 = io_cpu_fence_value & _T & _T_2 ? _GEN_1601 : meta_60_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2626 = io_cpu_fence_value & _T & _T_2 ? _GEN_1602 : meta_61_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2627 = io_cpu_fence_value & _T & _T_2 ? _GEN_1603 : meta_62_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2628 = io_cpu_fence_value & _T & _T_2 ? _GEN_1604 : meta_63_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2629 = io_cpu_fence_value & _T & _T_2 ? _GEN_1605 : meta_64_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2630 = io_cpu_fence_value & _T & _T_2 ? _GEN_1606 : meta_65_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2631 = io_cpu_fence_value & _T & _T_2 ? _GEN_1607 : meta_66_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2632 = io_cpu_fence_value & _T & _T_2 ? _GEN_1608 : meta_67_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2633 = io_cpu_fence_value & _T & _T_2 ? _GEN_1609 : meta_68_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2634 = io_cpu_fence_value & _T & _T_2 ? _GEN_1610 : meta_69_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2635 = io_cpu_fence_value & _T & _T_2 ? _GEN_1611 : meta_70_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2636 = io_cpu_fence_value & _T & _T_2 ? _GEN_1612 : meta_71_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2637 = io_cpu_fence_value & _T & _T_2 ? _GEN_1613 : meta_72_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2638 = io_cpu_fence_value & _T & _T_2 ? _GEN_1614 : meta_73_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2639 = io_cpu_fence_value & _T & _T_2 ? _GEN_1615 : meta_74_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2640 = io_cpu_fence_value & _T & _T_2 ? _GEN_1616 : meta_75_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2641 = io_cpu_fence_value & _T & _T_2 ? _GEN_1617 : meta_76_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2642 = io_cpu_fence_value & _T & _T_2 ? _GEN_1618 : meta_77_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2643 = io_cpu_fence_value & _T & _T_2 ? _GEN_1619 : meta_78_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2644 = io_cpu_fence_value & _T & _T_2 ? _GEN_1620 : meta_79_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2645 = io_cpu_fence_value & _T & _T_2 ? _GEN_1621 : meta_80_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2646 = io_cpu_fence_value & _T & _T_2 ? _GEN_1622 : meta_81_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2647 = io_cpu_fence_value & _T & _T_2 ? _GEN_1623 : meta_82_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2648 = io_cpu_fence_value & _T & _T_2 ? _GEN_1624 : meta_83_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2649 = io_cpu_fence_value & _T & _T_2 ? _GEN_1625 : meta_84_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2650 = io_cpu_fence_value & _T & _T_2 ? _GEN_1626 : meta_85_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2651 = io_cpu_fence_value & _T & _T_2 ? _GEN_1627 : meta_86_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2652 = io_cpu_fence_value & _T & _T_2 ? _GEN_1628 : meta_87_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2653 = io_cpu_fence_value & _T & _T_2 ? _GEN_1629 : meta_88_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2654 = io_cpu_fence_value & _T & _T_2 ? _GEN_1630 : meta_89_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2655 = io_cpu_fence_value & _T & _T_2 ? _GEN_1631 : meta_90_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2656 = io_cpu_fence_value & _T & _T_2 ? _GEN_1632 : meta_91_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2657 = io_cpu_fence_value & _T & _T_2 ? _GEN_1633 : meta_92_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2658 = io_cpu_fence_value & _T & _T_2 ? _GEN_1634 : meta_93_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2659 = io_cpu_fence_value & _T & _T_2 ? _GEN_1635 : meta_94_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2660 = io_cpu_fence_value & _T & _T_2 ? _GEN_1636 : meta_95_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2661 = io_cpu_fence_value & _T & _T_2 ? _GEN_1637 : meta_96_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2662 = io_cpu_fence_value & _T & _T_2 ? _GEN_1638 : meta_97_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2663 = io_cpu_fence_value & _T & _T_2 ? _GEN_1639 : meta_98_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2664 = io_cpu_fence_value & _T & _T_2 ? _GEN_1640 : meta_99_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2665 = io_cpu_fence_value & _T & _T_2 ? _GEN_1641 : meta_100_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2666 = io_cpu_fence_value & _T & _T_2 ? _GEN_1642 : meta_101_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2667 = io_cpu_fence_value & _T & _T_2 ? _GEN_1643 : meta_102_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2668 = io_cpu_fence_value & _T & _T_2 ? _GEN_1644 : meta_103_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2669 = io_cpu_fence_value & _T & _T_2 ? _GEN_1645 : meta_104_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2670 = io_cpu_fence_value & _T & _T_2 ? _GEN_1646 : meta_105_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2671 = io_cpu_fence_value & _T & _T_2 ? _GEN_1647 : meta_106_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2672 = io_cpu_fence_value & _T & _T_2 ? _GEN_1648 : meta_107_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2673 = io_cpu_fence_value & _T & _T_2 ? _GEN_1649 : meta_108_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2674 = io_cpu_fence_value & _T & _T_2 ? _GEN_1650 : meta_109_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2675 = io_cpu_fence_value & _T & _T_2 ? _GEN_1651 : meta_110_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2676 = io_cpu_fence_value & _T & _T_2 ? _GEN_1652 : meta_111_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2677 = io_cpu_fence_value & _T & _T_2 ? _GEN_1653 : meta_112_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2678 = io_cpu_fence_value & _T & _T_2 ? _GEN_1654 : meta_113_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2679 = io_cpu_fence_value & _T & _T_2 ? _GEN_1655 : meta_114_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2680 = io_cpu_fence_value & _T & _T_2 ? _GEN_1656 : meta_115_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2681 = io_cpu_fence_value & _T & _T_2 ? _GEN_1657 : meta_116_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2682 = io_cpu_fence_value & _T & _T_2 ? _GEN_1658 : meta_117_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2683 = io_cpu_fence_value & _T & _T_2 ? _GEN_1659 : meta_118_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2684 = io_cpu_fence_value & _T & _T_2 ? _GEN_1660 : meta_119_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2685 = io_cpu_fence_value & _T & _T_2 ? _GEN_1661 : meta_120_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2686 = io_cpu_fence_value & _T & _T_2 ? _GEN_1662 : meta_121_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2687 = io_cpu_fence_value & _T & _T_2 ? _GEN_1663 : meta_122_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2688 = io_cpu_fence_value & _T & _T_2 ? _GEN_1664 : meta_123_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2689 = io_cpu_fence_value & _T & _T_2 ? _GEN_1665 : meta_124_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2690 = io_cpu_fence_value & _T & _T_2 ? _GEN_1666 : meta_125_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2691 = io_cpu_fence_value & _T & _T_2 ? _GEN_1667 : meta_126_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2692 = io_cpu_fence_value & _T & _T_2 ? _GEN_1668 : meta_127_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2693 = io_cpu_fence_value & _T & _T_2 ? _GEN_1669 : meta_128_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2694 = io_cpu_fence_value & _T & _T_2 ? _GEN_1670 : meta_129_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2695 = io_cpu_fence_value & _T & _T_2 ? _GEN_1671 : meta_130_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2696 = io_cpu_fence_value & _T & _T_2 ? _GEN_1672 : meta_131_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2697 = io_cpu_fence_value & _T & _T_2 ? _GEN_1673 : meta_132_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2698 = io_cpu_fence_value & _T & _T_2 ? _GEN_1674 : meta_133_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2699 = io_cpu_fence_value & _T & _T_2 ? _GEN_1675 : meta_134_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2700 = io_cpu_fence_value & _T & _T_2 ? _GEN_1676 : meta_135_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2701 = io_cpu_fence_value & _T & _T_2 ? _GEN_1677 : meta_136_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2702 = io_cpu_fence_value & _T & _T_2 ? _GEN_1678 : meta_137_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2703 = io_cpu_fence_value & _T & _T_2 ? _GEN_1679 : meta_138_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2704 = io_cpu_fence_value & _T & _T_2 ? _GEN_1680 : meta_139_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2705 = io_cpu_fence_value & _T & _T_2 ? _GEN_1681 : meta_140_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2706 = io_cpu_fence_value & _T & _T_2 ? _GEN_1682 : meta_141_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2707 = io_cpu_fence_value & _T & _T_2 ? _GEN_1683 : meta_142_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2708 = io_cpu_fence_value & _T & _T_2 ? _GEN_1684 : meta_143_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2709 = io_cpu_fence_value & _T & _T_2 ? _GEN_1685 : meta_144_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2710 = io_cpu_fence_value & _T & _T_2 ? _GEN_1686 : meta_145_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2711 = io_cpu_fence_value & _T & _T_2 ? _GEN_1687 : meta_146_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2712 = io_cpu_fence_value & _T & _T_2 ? _GEN_1688 : meta_147_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2713 = io_cpu_fence_value & _T & _T_2 ? _GEN_1689 : meta_148_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2714 = io_cpu_fence_value & _T & _T_2 ? _GEN_1690 : meta_149_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2715 = io_cpu_fence_value & _T & _T_2 ? _GEN_1691 : meta_150_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2716 = io_cpu_fence_value & _T & _T_2 ? _GEN_1692 : meta_151_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2717 = io_cpu_fence_value & _T & _T_2 ? _GEN_1693 : meta_152_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2718 = io_cpu_fence_value & _T & _T_2 ? _GEN_1694 : meta_153_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2719 = io_cpu_fence_value & _T & _T_2 ? _GEN_1695 : meta_154_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2720 = io_cpu_fence_value & _T & _T_2 ? _GEN_1696 : meta_155_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2721 = io_cpu_fence_value & _T & _T_2 ? _GEN_1697 : meta_156_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2722 = io_cpu_fence_value & _T & _T_2 ? _GEN_1698 : meta_157_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2723 = io_cpu_fence_value & _T & _T_2 ? _GEN_1699 : meta_158_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2724 = io_cpu_fence_value & _T & _T_2 ? _GEN_1700 : meta_159_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2725 = io_cpu_fence_value & _T & _T_2 ? _GEN_1701 : meta_160_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2726 = io_cpu_fence_value & _T & _T_2 ? _GEN_1702 : meta_161_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2727 = io_cpu_fence_value & _T & _T_2 ? _GEN_1703 : meta_162_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2728 = io_cpu_fence_value & _T & _T_2 ? _GEN_1704 : meta_163_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2729 = io_cpu_fence_value & _T & _T_2 ? _GEN_1705 : meta_164_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2730 = io_cpu_fence_value & _T & _T_2 ? _GEN_1706 : meta_165_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2731 = io_cpu_fence_value & _T & _T_2 ? _GEN_1707 : meta_166_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2732 = io_cpu_fence_value & _T & _T_2 ? _GEN_1708 : meta_167_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2733 = io_cpu_fence_value & _T & _T_2 ? _GEN_1709 : meta_168_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2734 = io_cpu_fence_value & _T & _T_2 ? _GEN_1710 : meta_169_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2735 = io_cpu_fence_value & _T & _T_2 ? _GEN_1711 : meta_170_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2736 = io_cpu_fence_value & _T & _T_2 ? _GEN_1712 : meta_171_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2737 = io_cpu_fence_value & _T & _T_2 ? _GEN_1713 : meta_172_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2738 = io_cpu_fence_value & _T & _T_2 ? _GEN_1714 : meta_173_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2739 = io_cpu_fence_value & _T & _T_2 ? _GEN_1715 : meta_174_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2740 = io_cpu_fence_value & _T & _T_2 ? _GEN_1716 : meta_175_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2741 = io_cpu_fence_value & _T & _T_2 ? _GEN_1717 : meta_176_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2742 = io_cpu_fence_value & _T & _T_2 ? _GEN_1718 : meta_177_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2743 = io_cpu_fence_value & _T & _T_2 ? _GEN_1719 : meta_178_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2744 = io_cpu_fence_value & _T & _T_2 ? _GEN_1720 : meta_179_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2745 = io_cpu_fence_value & _T & _T_2 ? _GEN_1721 : meta_180_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2746 = io_cpu_fence_value & _T & _T_2 ? _GEN_1722 : meta_181_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2747 = io_cpu_fence_value & _T & _T_2 ? _GEN_1723 : meta_182_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2748 = io_cpu_fence_value & _T & _T_2 ? _GEN_1724 : meta_183_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2749 = io_cpu_fence_value & _T & _T_2 ? _GEN_1725 : meta_184_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2750 = io_cpu_fence_value & _T & _T_2 ? _GEN_1726 : meta_185_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2751 = io_cpu_fence_value & _T & _T_2 ? _GEN_1727 : meta_186_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2752 = io_cpu_fence_value & _T & _T_2 ? _GEN_1728 : meta_187_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2753 = io_cpu_fence_value & _T & _T_2 ? _GEN_1729 : meta_188_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2754 = io_cpu_fence_value & _T & _T_2 ? _GEN_1730 : meta_189_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2755 = io_cpu_fence_value & _T & _T_2 ? _GEN_1731 : meta_190_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2756 = io_cpu_fence_value & _T & _T_2 ? _GEN_1732 : meta_191_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2757 = io_cpu_fence_value & _T & _T_2 ? _GEN_1733 : meta_192_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2758 = io_cpu_fence_value & _T & _T_2 ? _GEN_1734 : meta_193_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2759 = io_cpu_fence_value & _T & _T_2 ? _GEN_1735 : meta_194_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2760 = io_cpu_fence_value & _T & _T_2 ? _GEN_1736 : meta_195_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2761 = io_cpu_fence_value & _T & _T_2 ? _GEN_1737 : meta_196_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2762 = io_cpu_fence_value & _T & _T_2 ? _GEN_1738 : meta_197_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2763 = io_cpu_fence_value & _T & _T_2 ? _GEN_1739 : meta_198_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2764 = io_cpu_fence_value & _T & _T_2 ? _GEN_1740 : meta_199_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2765 = io_cpu_fence_value & _T & _T_2 ? _GEN_1741 : meta_200_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2766 = io_cpu_fence_value & _T & _T_2 ? _GEN_1742 : meta_201_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2767 = io_cpu_fence_value & _T & _T_2 ? _GEN_1743 : meta_202_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2768 = io_cpu_fence_value & _T & _T_2 ? _GEN_1744 : meta_203_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2769 = io_cpu_fence_value & _T & _T_2 ? _GEN_1745 : meta_204_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2770 = io_cpu_fence_value & _T & _T_2 ? _GEN_1746 : meta_205_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2771 = io_cpu_fence_value & _T & _T_2 ? _GEN_1747 : meta_206_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2772 = io_cpu_fence_value & _T & _T_2 ? _GEN_1748 : meta_207_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2773 = io_cpu_fence_value & _T & _T_2 ? _GEN_1749 : meta_208_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2774 = io_cpu_fence_value & _T & _T_2 ? _GEN_1750 : meta_209_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2775 = io_cpu_fence_value & _T & _T_2 ? _GEN_1751 : meta_210_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2776 = io_cpu_fence_value & _T & _T_2 ? _GEN_1752 : meta_211_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2777 = io_cpu_fence_value & _T & _T_2 ? _GEN_1753 : meta_212_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2778 = io_cpu_fence_value & _T & _T_2 ? _GEN_1754 : meta_213_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2779 = io_cpu_fence_value & _T & _T_2 ? _GEN_1755 : meta_214_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2780 = io_cpu_fence_value & _T & _T_2 ? _GEN_1756 : meta_215_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2781 = io_cpu_fence_value & _T & _T_2 ? _GEN_1757 : meta_216_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2782 = io_cpu_fence_value & _T & _T_2 ? _GEN_1758 : meta_217_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2783 = io_cpu_fence_value & _T & _T_2 ? _GEN_1759 : meta_218_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2784 = io_cpu_fence_value & _T & _T_2 ? _GEN_1760 : meta_219_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2785 = io_cpu_fence_value & _T & _T_2 ? _GEN_1761 : meta_220_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2786 = io_cpu_fence_value & _T & _T_2 ? _GEN_1762 : meta_221_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2787 = io_cpu_fence_value & _T & _T_2 ? _GEN_1763 : meta_222_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2788 = io_cpu_fence_value & _T & _T_2 ? _GEN_1764 : meta_223_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2789 = io_cpu_fence_value & _T & _T_2 ? _GEN_1765 : meta_224_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2790 = io_cpu_fence_value & _T & _T_2 ? _GEN_1766 : meta_225_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2791 = io_cpu_fence_value & _T & _T_2 ? _GEN_1767 : meta_226_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2792 = io_cpu_fence_value & _T & _T_2 ? _GEN_1768 : meta_227_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2793 = io_cpu_fence_value & _T & _T_2 ? _GEN_1769 : meta_228_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2794 = io_cpu_fence_value & _T & _T_2 ? _GEN_1770 : meta_229_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2795 = io_cpu_fence_value & _T & _T_2 ? _GEN_1771 : meta_230_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2796 = io_cpu_fence_value & _T & _T_2 ? _GEN_1772 : meta_231_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2797 = io_cpu_fence_value & _T & _T_2 ? _GEN_1773 : meta_232_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2798 = io_cpu_fence_value & _T & _T_2 ? _GEN_1774 : meta_233_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2799 = io_cpu_fence_value & _T & _T_2 ? _GEN_1775 : meta_234_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2800 = io_cpu_fence_value & _T & _T_2 ? _GEN_1776 : meta_235_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2801 = io_cpu_fence_value & _T & _T_2 ? _GEN_1777 : meta_236_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2802 = io_cpu_fence_value & _T & _T_2 ? _GEN_1778 : meta_237_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2803 = io_cpu_fence_value & _T & _T_2 ? _GEN_1779 : meta_238_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2804 = io_cpu_fence_value & _T & _T_2 ? _GEN_1780 : meta_239_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2805 = io_cpu_fence_value & _T & _T_2 ? _GEN_1781 : meta_240_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2806 = io_cpu_fence_value & _T & _T_2 ? _GEN_1782 : meta_241_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2807 = io_cpu_fence_value & _T & _T_2 ? _GEN_1783 : meta_242_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2808 = io_cpu_fence_value & _T & _T_2 ? _GEN_1784 : meta_243_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2809 = io_cpu_fence_value & _T & _T_2 ? _GEN_1785 : meta_244_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2810 = io_cpu_fence_value & _T & _T_2 ? _GEN_1786 : meta_245_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2811 = io_cpu_fence_value & _T & _T_2 ? _GEN_1787 : meta_246_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2812 = io_cpu_fence_value & _T & _T_2 ? _GEN_1788 : meta_247_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2813 = io_cpu_fence_value & _T & _T_2 ? _GEN_1789 : meta_248_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2814 = io_cpu_fence_value & _T & _T_2 ? _GEN_1790 : meta_249_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2815 = io_cpu_fence_value & _T & _T_2 ? _GEN_1791 : meta_250_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2816 = io_cpu_fence_value & _T & _T_2 ? _GEN_1792 : meta_251_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2817 = io_cpu_fence_value & _T & _T_2 ? _GEN_1793 : meta_252_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2818 = io_cpu_fence_value & _T & _T_2 ? _GEN_1794 : meta_253_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2819 = io_cpu_fence_value & _T & _T_2 ? _GEN_1795 : meta_254_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2820 = io_cpu_fence_value & _T & _T_2 ? _GEN_1796 : meta_255_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2821 = io_cpu_fence_value & _T & _T_2 ? _GEN_1797 : meta_256_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2822 = io_cpu_fence_value & _T & _T_2 ? _GEN_1798 : meta_257_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2823 = io_cpu_fence_value & _T & _T_2 ? _GEN_1799 : meta_258_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2824 = io_cpu_fence_value & _T & _T_2 ? _GEN_1800 : meta_259_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2825 = io_cpu_fence_value & _T & _T_2 ? _GEN_1801 : meta_260_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2826 = io_cpu_fence_value & _T & _T_2 ? _GEN_1802 : meta_261_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2827 = io_cpu_fence_value & _T & _T_2 ? _GEN_1803 : meta_262_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2828 = io_cpu_fence_value & _T & _T_2 ? _GEN_1804 : meta_263_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2829 = io_cpu_fence_value & _T & _T_2 ? _GEN_1805 : meta_264_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2830 = io_cpu_fence_value & _T & _T_2 ? _GEN_1806 : meta_265_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2831 = io_cpu_fence_value & _T & _T_2 ? _GEN_1807 : meta_266_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2832 = io_cpu_fence_value & _T & _T_2 ? _GEN_1808 : meta_267_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2833 = io_cpu_fence_value & _T & _T_2 ? _GEN_1809 : meta_268_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2834 = io_cpu_fence_value & _T & _T_2 ? _GEN_1810 : meta_269_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2835 = io_cpu_fence_value & _T & _T_2 ? _GEN_1811 : meta_270_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2836 = io_cpu_fence_value & _T & _T_2 ? _GEN_1812 : meta_271_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2837 = io_cpu_fence_value & _T & _T_2 ? _GEN_1813 : meta_272_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2838 = io_cpu_fence_value & _T & _T_2 ? _GEN_1814 : meta_273_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2839 = io_cpu_fence_value & _T & _T_2 ? _GEN_1815 : meta_274_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2840 = io_cpu_fence_value & _T & _T_2 ? _GEN_1816 : meta_275_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2841 = io_cpu_fence_value & _T & _T_2 ? _GEN_1817 : meta_276_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2842 = io_cpu_fence_value & _T & _T_2 ? _GEN_1818 : meta_277_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2843 = io_cpu_fence_value & _T & _T_2 ? _GEN_1819 : meta_278_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2844 = io_cpu_fence_value & _T & _T_2 ? _GEN_1820 : meta_279_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2845 = io_cpu_fence_value & _T & _T_2 ? _GEN_1821 : meta_280_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2846 = io_cpu_fence_value & _T & _T_2 ? _GEN_1822 : meta_281_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2847 = io_cpu_fence_value & _T & _T_2 ? _GEN_1823 : meta_282_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2848 = io_cpu_fence_value & _T & _T_2 ? _GEN_1824 : meta_283_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2849 = io_cpu_fence_value & _T & _T_2 ? _GEN_1825 : meta_284_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2850 = io_cpu_fence_value & _T & _T_2 ? _GEN_1826 : meta_285_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2851 = io_cpu_fence_value & _T & _T_2 ? _GEN_1827 : meta_286_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2852 = io_cpu_fence_value & _T & _T_2 ? _GEN_1828 : meta_287_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2853 = io_cpu_fence_value & _T & _T_2 ? _GEN_1829 : meta_288_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2854 = io_cpu_fence_value & _T & _T_2 ? _GEN_1830 : meta_289_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2855 = io_cpu_fence_value & _T & _T_2 ? _GEN_1831 : meta_290_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2856 = io_cpu_fence_value & _T & _T_2 ? _GEN_1832 : meta_291_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2857 = io_cpu_fence_value & _T & _T_2 ? _GEN_1833 : meta_292_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2858 = io_cpu_fence_value & _T & _T_2 ? _GEN_1834 : meta_293_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2859 = io_cpu_fence_value & _T & _T_2 ? _GEN_1835 : meta_294_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2860 = io_cpu_fence_value & _T & _T_2 ? _GEN_1836 : meta_295_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2861 = io_cpu_fence_value & _T & _T_2 ? _GEN_1837 : meta_296_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2862 = io_cpu_fence_value & _T & _T_2 ? _GEN_1838 : meta_297_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2863 = io_cpu_fence_value & _T & _T_2 ? _GEN_1839 : meta_298_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2864 = io_cpu_fence_value & _T & _T_2 ? _GEN_1840 : meta_299_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2865 = io_cpu_fence_value & _T & _T_2 ? _GEN_1841 : meta_300_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2866 = io_cpu_fence_value & _T & _T_2 ? _GEN_1842 : meta_301_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2867 = io_cpu_fence_value & _T & _T_2 ? _GEN_1843 : meta_302_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2868 = io_cpu_fence_value & _T & _T_2 ? _GEN_1844 : meta_303_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2869 = io_cpu_fence_value & _T & _T_2 ? _GEN_1845 : meta_304_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2870 = io_cpu_fence_value & _T & _T_2 ? _GEN_1846 : meta_305_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2871 = io_cpu_fence_value & _T & _T_2 ? _GEN_1847 : meta_306_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2872 = io_cpu_fence_value & _T & _T_2 ? _GEN_1848 : meta_307_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2873 = io_cpu_fence_value & _T & _T_2 ? _GEN_1849 : meta_308_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2874 = io_cpu_fence_value & _T & _T_2 ? _GEN_1850 : meta_309_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2875 = io_cpu_fence_value & _T & _T_2 ? _GEN_1851 : meta_310_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2876 = io_cpu_fence_value & _T & _T_2 ? _GEN_1852 : meta_311_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2877 = io_cpu_fence_value & _T & _T_2 ? _GEN_1853 : meta_312_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2878 = io_cpu_fence_value & _T & _T_2 ? _GEN_1854 : meta_313_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2879 = io_cpu_fence_value & _T & _T_2 ? _GEN_1855 : meta_314_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2880 = io_cpu_fence_value & _T & _T_2 ? _GEN_1856 : meta_315_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2881 = io_cpu_fence_value & _T & _T_2 ? _GEN_1857 : meta_316_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2882 = io_cpu_fence_value & _T & _T_2 ? _GEN_1858 : meta_317_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2883 = io_cpu_fence_value & _T & _T_2 ? _GEN_1859 : meta_318_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2884 = io_cpu_fence_value & _T & _T_2 ? _GEN_1860 : meta_319_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2885 = io_cpu_fence_value & _T & _T_2 ? _GEN_1861 : meta_320_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2886 = io_cpu_fence_value & _T & _T_2 ? _GEN_1862 : meta_321_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2887 = io_cpu_fence_value & _T & _T_2 ? _GEN_1863 : meta_322_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2888 = io_cpu_fence_value & _T & _T_2 ? _GEN_1864 : meta_323_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2889 = io_cpu_fence_value & _T & _T_2 ? _GEN_1865 : meta_324_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2890 = io_cpu_fence_value & _T & _T_2 ? _GEN_1866 : meta_325_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2891 = io_cpu_fence_value & _T & _T_2 ? _GEN_1867 : meta_326_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2892 = io_cpu_fence_value & _T & _T_2 ? _GEN_1868 : meta_327_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2893 = io_cpu_fence_value & _T & _T_2 ? _GEN_1869 : meta_328_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2894 = io_cpu_fence_value & _T & _T_2 ? _GEN_1870 : meta_329_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2895 = io_cpu_fence_value & _T & _T_2 ? _GEN_1871 : meta_330_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2896 = io_cpu_fence_value & _T & _T_2 ? _GEN_1872 : meta_331_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2897 = io_cpu_fence_value & _T & _T_2 ? _GEN_1873 : meta_332_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2898 = io_cpu_fence_value & _T & _T_2 ? _GEN_1874 : meta_333_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2899 = io_cpu_fence_value & _T & _T_2 ? _GEN_1875 : meta_334_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2900 = io_cpu_fence_value & _T & _T_2 ? _GEN_1876 : meta_335_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2901 = io_cpu_fence_value & _T & _T_2 ? _GEN_1877 : meta_336_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2902 = io_cpu_fence_value & _T & _T_2 ? _GEN_1878 : meta_337_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2903 = io_cpu_fence_value & _T & _T_2 ? _GEN_1879 : meta_338_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2904 = io_cpu_fence_value & _T & _T_2 ? _GEN_1880 : meta_339_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2905 = io_cpu_fence_value & _T & _T_2 ? _GEN_1881 : meta_340_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2906 = io_cpu_fence_value & _T & _T_2 ? _GEN_1882 : meta_341_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2907 = io_cpu_fence_value & _T & _T_2 ? _GEN_1883 : meta_342_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2908 = io_cpu_fence_value & _T & _T_2 ? _GEN_1884 : meta_343_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2909 = io_cpu_fence_value & _T & _T_2 ? _GEN_1885 : meta_344_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2910 = io_cpu_fence_value & _T & _T_2 ? _GEN_1886 : meta_345_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2911 = io_cpu_fence_value & _T & _T_2 ? _GEN_1887 : meta_346_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2912 = io_cpu_fence_value & _T & _T_2 ? _GEN_1888 : meta_347_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2913 = io_cpu_fence_value & _T & _T_2 ? _GEN_1889 : meta_348_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2914 = io_cpu_fence_value & _T & _T_2 ? _GEN_1890 : meta_349_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2915 = io_cpu_fence_value & _T & _T_2 ? _GEN_1891 : meta_350_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2916 = io_cpu_fence_value & _T & _T_2 ? _GEN_1892 : meta_351_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2917 = io_cpu_fence_value & _T & _T_2 ? _GEN_1893 : meta_352_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2918 = io_cpu_fence_value & _T & _T_2 ? _GEN_1894 : meta_353_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2919 = io_cpu_fence_value & _T & _T_2 ? _GEN_1895 : meta_354_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2920 = io_cpu_fence_value & _T & _T_2 ? _GEN_1896 : meta_355_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2921 = io_cpu_fence_value & _T & _T_2 ? _GEN_1897 : meta_356_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2922 = io_cpu_fence_value & _T & _T_2 ? _GEN_1898 : meta_357_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2923 = io_cpu_fence_value & _T & _T_2 ? _GEN_1899 : meta_358_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2924 = io_cpu_fence_value & _T & _T_2 ? _GEN_1900 : meta_359_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2925 = io_cpu_fence_value & _T & _T_2 ? _GEN_1901 : meta_360_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2926 = io_cpu_fence_value & _T & _T_2 ? _GEN_1902 : meta_361_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2927 = io_cpu_fence_value & _T & _T_2 ? _GEN_1903 : meta_362_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2928 = io_cpu_fence_value & _T & _T_2 ? _GEN_1904 : meta_363_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2929 = io_cpu_fence_value & _T & _T_2 ? _GEN_1905 : meta_364_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2930 = io_cpu_fence_value & _T & _T_2 ? _GEN_1906 : meta_365_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2931 = io_cpu_fence_value & _T & _T_2 ? _GEN_1907 : meta_366_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2932 = io_cpu_fence_value & _T & _T_2 ? _GEN_1908 : meta_367_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2933 = io_cpu_fence_value & _T & _T_2 ? _GEN_1909 : meta_368_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2934 = io_cpu_fence_value & _T & _T_2 ? _GEN_1910 : meta_369_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2935 = io_cpu_fence_value & _T & _T_2 ? _GEN_1911 : meta_370_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2936 = io_cpu_fence_value & _T & _T_2 ? _GEN_1912 : meta_371_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2937 = io_cpu_fence_value & _T & _T_2 ? _GEN_1913 : meta_372_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2938 = io_cpu_fence_value & _T & _T_2 ? _GEN_1914 : meta_373_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2939 = io_cpu_fence_value & _T & _T_2 ? _GEN_1915 : meta_374_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2940 = io_cpu_fence_value & _T & _T_2 ? _GEN_1916 : meta_375_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2941 = io_cpu_fence_value & _T & _T_2 ? _GEN_1917 : meta_376_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2942 = io_cpu_fence_value & _T & _T_2 ? _GEN_1918 : meta_377_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2943 = io_cpu_fence_value & _T & _T_2 ? _GEN_1919 : meta_378_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2944 = io_cpu_fence_value & _T & _T_2 ? _GEN_1920 : meta_379_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2945 = io_cpu_fence_value & _T & _T_2 ? _GEN_1921 : meta_380_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2946 = io_cpu_fence_value & _T & _T_2 ? _GEN_1922 : meta_381_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2947 = io_cpu_fence_value & _T & _T_2 ? _GEN_1923 : meta_382_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2948 = io_cpu_fence_value & _T & _T_2 ? _GEN_1924 : meta_383_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2949 = io_cpu_fence_value & _T & _T_2 ? _GEN_1925 : meta_384_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2950 = io_cpu_fence_value & _T & _T_2 ? _GEN_1926 : meta_385_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2951 = io_cpu_fence_value & _T & _T_2 ? _GEN_1927 : meta_386_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2952 = io_cpu_fence_value & _T & _T_2 ? _GEN_1928 : meta_387_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2953 = io_cpu_fence_value & _T & _T_2 ? _GEN_1929 : meta_388_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2954 = io_cpu_fence_value & _T & _T_2 ? _GEN_1930 : meta_389_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2955 = io_cpu_fence_value & _T & _T_2 ? _GEN_1931 : meta_390_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2956 = io_cpu_fence_value & _T & _T_2 ? _GEN_1932 : meta_391_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2957 = io_cpu_fence_value & _T & _T_2 ? _GEN_1933 : meta_392_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2958 = io_cpu_fence_value & _T & _T_2 ? _GEN_1934 : meta_393_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2959 = io_cpu_fence_value & _T & _T_2 ? _GEN_1935 : meta_394_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2960 = io_cpu_fence_value & _T & _T_2 ? _GEN_1936 : meta_395_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2961 = io_cpu_fence_value & _T & _T_2 ? _GEN_1937 : meta_396_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2962 = io_cpu_fence_value & _T & _T_2 ? _GEN_1938 : meta_397_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2963 = io_cpu_fence_value & _T & _T_2 ? _GEN_1939 : meta_398_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2964 = io_cpu_fence_value & _T & _T_2 ? _GEN_1940 : meta_399_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2965 = io_cpu_fence_value & _T & _T_2 ? _GEN_1941 : meta_400_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2966 = io_cpu_fence_value & _T & _T_2 ? _GEN_1942 : meta_401_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2967 = io_cpu_fence_value & _T & _T_2 ? _GEN_1943 : meta_402_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2968 = io_cpu_fence_value & _T & _T_2 ? _GEN_1944 : meta_403_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2969 = io_cpu_fence_value & _T & _T_2 ? _GEN_1945 : meta_404_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2970 = io_cpu_fence_value & _T & _T_2 ? _GEN_1946 : meta_405_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2971 = io_cpu_fence_value & _T & _T_2 ? _GEN_1947 : meta_406_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2972 = io_cpu_fence_value & _T & _T_2 ? _GEN_1948 : meta_407_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2973 = io_cpu_fence_value & _T & _T_2 ? _GEN_1949 : meta_408_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2974 = io_cpu_fence_value & _T & _T_2 ? _GEN_1950 : meta_409_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2975 = io_cpu_fence_value & _T & _T_2 ? _GEN_1951 : meta_410_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2976 = io_cpu_fence_value & _T & _T_2 ? _GEN_1952 : meta_411_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2977 = io_cpu_fence_value & _T & _T_2 ? _GEN_1953 : meta_412_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2978 = io_cpu_fence_value & _T & _T_2 ? _GEN_1954 : meta_413_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2979 = io_cpu_fence_value & _T & _T_2 ? _GEN_1955 : meta_414_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2980 = io_cpu_fence_value & _T & _T_2 ? _GEN_1956 : meta_415_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2981 = io_cpu_fence_value & _T & _T_2 ? _GEN_1957 : meta_416_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2982 = io_cpu_fence_value & _T & _T_2 ? _GEN_1958 : meta_417_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2983 = io_cpu_fence_value & _T & _T_2 ? _GEN_1959 : meta_418_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2984 = io_cpu_fence_value & _T & _T_2 ? _GEN_1960 : meta_419_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2985 = io_cpu_fence_value & _T & _T_2 ? _GEN_1961 : meta_420_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2986 = io_cpu_fence_value & _T & _T_2 ? _GEN_1962 : meta_421_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2987 = io_cpu_fence_value & _T & _T_2 ? _GEN_1963 : meta_422_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2988 = io_cpu_fence_value & _T & _T_2 ? _GEN_1964 : meta_423_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2989 = io_cpu_fence_value & _T & _T_2 ? _GEN_1965 : meta_424_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2990 = io_cpu_fence_value & _T & _T_2 ? _GEN_1966 : meta_425_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2991 = io_cpu_fence_value & _T & _T_2 ? _GEN_1967 : meta_426_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2992 = io_cpu_fence_value & _T & _T_2 ? _GEN_1968 : meta_427_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2993 = io_cpu_fence_value & _T & _T_2 ? _GEN_1969 : meta_428_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2994 = io_cpu_fence_value & _T & _T_2 ? _GEN_1970 : meta_429_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2995 = io_cpu_fence_value & _T & _T_2 ? _GEN_1971 : meta_430_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2996 = io_cpu_fence_value & _T & _T_2 ? _GEN_1972 : meta_431_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2997 = io_cpu_fence_value & _T & _T_2 ? _GEN_1973 : meta_432_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2998 = io_cpu_fence_value & _T & _T_2 ? _GEN_1974 : meta_433_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_2999 = io_cpu_fence_value & _T & _T_2 ? _GEN_1975 : meta_434_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3000 = io_cpu_fence_value & _T & _T_2 ? _GEN_1976 : meta_435_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3001 = io_cpu_fence_value & _T & _T_2 ? _GEN_1977 : meta_436_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3002 = io_cpu_fence_value & _T & _T_2 ? _GEN_1978 : meta_437_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3003 = io_cpu_fence_value & _T & _T_2 ? _GEN_1979 : meta_438_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3004 = io_cpu_fence_value & _T & _T_2 ? _GEN_1980 : meta_439_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3005 = io_cpu_fence_value & _T & _T_2 ? _GEN_1981 : meta_440_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3006 = io_cpu_fence_value & _T & _T_2 ? _GEN_1982 : meta_441_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3007 = io_cpu_fence_value & _T & _T_2 ? _GEN_1983 : meta_442_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3008 = io_cpu_fence_value & _T & _T_2 ? _GEN_1984 : meta_443_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3009 = io_cpu_fence_value & _T & _T_2 ? _GEN_1985 : meta_444_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3010 = io_cpu_fence_value & _T & _T_2 ? _GEN_1986 : meta_445_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3011 = io_cpu_fence_value & _T & _T_2 ? _GEN_1987 : meta_446_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3012 = io_cpu_fence_value & _T & _T_2 ? _GEN_1988 : meta_447_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3013 = io_cpu_fence_value & _T & _T_2 ? _GEN_1989 : meta_448_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3014 = io_cpu_fence_value & _T & _T_2 ? _GEN_1990 : meta_449_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3015 = io_cpu_fence_value & _T & _T_2 ? _GEN_1991 : meta_450_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3016 = io_cpu_fence_value & _T & _T_2 ? _GEN_1992 : meta_451_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3017 = io_cpu_fence_value & _T & _T_2 ? _GEN_1993 : meta_452_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3018 = io_cpu_fence_value & _T & _T_2 ? _GEN_1994 : meta_453_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3019 = io_cpu_fence_value & _T & _T_2 ? _GEN_1995 : meta_454_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3020 = io_cpu_fence_value & _T & _T_2 ? _GEN_1996 : meta_455_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3021 = io_cpu_fence_value & _T & _T_2 ? _GEN_1997 : meta_456_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3022 = io_cpu_fence_value & _T & _T_2 ? _GEN_1998 : meta_457_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3023 = io_cpu_fence_value & _T & _T_2 ? _GEN_1999 : meta_458_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3024 = io_cpu_fence_value & _T & _T_2 ? _GEN_2000 : meta_459_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3025 = io_cpu_fence_value & _T & _T_2 ? _GEN_2001 : meta_460_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3026 = io_cpu_fence_value & _T & _T_2 ? _GEN_2002 : meta_461_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3027 = io_cpu_fence_value & _T & _T_2 ? _GEN_2003 : meta_462_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3028 = io_cpu_fence_value & _T & _T_2 ? _GEN_2004 : meta_463_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3029 = io_cpu_fence_value & _T & _T_2 ? _GEN_2005 : meta_464_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3030 = io_cpu_fence_value & _T & _T_2 ? _GEN_2006 : meta_465_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3031 = io_cpu_fence_value & _T & _T_2 ? _GEN_2007 : meta_466_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3032 = io_cpu_fence_value & _T & _T_2 ? _GEN_2008 : meta_467_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3033 = io_cpu_fence_value & _T & _T_2 ? _GEN_2009 : meta_468_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3034 = io_cpu_fence_value & _T & _T_2 ? _GEN_2010 : meta_469_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3035 = io_cpu_fence_value & _T & _T_2 ? _GEN_2011 : meta_470_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3036 = io_cpu_fence_value & _T & _T_2 ? _GEN_2012 : meta_471_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3037 = io_cpu_fence_value & _T & _T_2 ? _GEN_2013 : meta_472_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3038 = io_cpu_fence_value & _T & _T_2 ? _GEN_2014 : meta_473_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3039 = io_cpu_fence_value & _T & _T_2 ? _GEN_2015 : meta_474_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3040 = io_cpu_fence_value & _T & _T_2 ? _GEN_2016 : meta_475_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3041 = io_cpu_fence_value & _T & _T_2 ? _GEN_2017 : meta_476_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3042 = io_cpu_fence_value & _T & _T_2 ? _GEN_2018 : meta_477_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3043 = io_cpu_fence_value & _T & _T_2 ? _GEN_2019 : meta_478_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3044 = io_cpu_fence_value & _T & _T_2 ? _GEN_2020 : meta_479_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3045 = io_cpu_fence_value & _T & _T_2 ? _GEN_2021 : meta_480_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3046 = io_cpu_fence_value & _T & _T_2 ? _GEN_2022 : meta_481_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3047 = io_cpu_fence_value & _T & _T_2 ? _GEN_2023 : meta_482_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3048 = io_cpu_fence_value & _T & _T_2 ? _GEN_2024 : meta_483_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3049 = io_cpu_fence_value & _T & _T_2 ? _GEN_2025 : meta_484_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3050 = io_cpu_fence_value & _T & _T_2 ? _GEN_2026 : meta_485_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3051 = io_cpu_fence_value & _T & _T_2 ? _GEN_2027 : meta_486_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3052 = io_cpu_fence_value & _T & _T_2 ? _GEN_2028 : meta_487_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3053 = io_cpu_fence_value & _T & _T_2 ? _GEN_2029 : meta_488_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3054 = io_cpu_fence_value & _T & _T_2 ? _GEN_2030 : meta_489_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3055 = io_cpu_fence_value & _T & _T_2 ? _GEN_2031 : meta_490_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3056 = io_cpu_fence_value & _T & _T_2 ? _GEN_2032 : meta_491_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3057 = io_cpu_fence_value & _T & _T_2 ? _GEN_2033 : meta_492_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3058 = io_cpu_fence_value & _T & _T_2 ? _GEN_2034 : meta_493_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3059 = io_cpu_fence_value & _T & _T_2 ? _GEN_2035 : meta_494_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3060 = io_cpu_fence_value & _T & _T_2 ? _GEN_2036 : meta_495_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3061 = io_cpu_fence_value & _T & _T_2 ? _GEN_2037 : meta_496_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3062 = io_cpu_fence_value & _T & _T_2 ? _GEN_2038 : meta_497_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3063 = io_cpu_fence_value & _T & _T_2 ? _GEN_2039 : meta_498_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3064 = io_cpu_fence_value & _T & _T_2 ? _GEN_2040 : meta_499_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3065 = io_cpu_fence_value & _T & _T_2 ? _GEN_2041 : meta_500_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3066 = io_cpu_fence_value & _T & _T_2 ? _GEN_2042 : meta_501_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3067 = io_cpu_fence_value & _T & _T_2 ? _GEN_2043 : meta_502_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3068 = io_cpu_fence_value & _T & _T_2 ? _GEN_2044 : meta_503_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3069 = io_cpu_fence_value & _T & _T_2 ? _GEN_2045 : meta_504_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3070 = io_cpu_fence_value & _T & _T_2 ? _GEN_2046 : meta_505_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3071 = io_cpu_fence_value & _T & _T_2 ? _GEN_2047 : meta_506_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3072 = io_cpu_fence_value & _T & _T_2 ? _GEN_2048 : meta_507_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3073 = io_cpu_fence_value & _T & _T_2 ? _GEN_2049 : meta_508_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3074 = io_cpu_fence_value & _T & _T_2 ? _GEN_2050 : meta_509_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3075 = io_cpu_fence_value & _T & _T_2 ? _GEN_2051 : meta_510_valid_1; // @[ICache.scala 136:73 34:21]
  wire  _GEN_3076 = io_cpu_fence_value & _T & _T_2 ? _GEN_2052 : meta_511_valid_1; // @[ICache.scala 136:73 34:21]
  reg [31:0] ar_addr; // @[ICache.scala 141:24]
  reg [7:0] ar_len; // @[ICache.scala 141:24]
  reg [2:0] ar_size; // @[ICache.scala 141:24]
  reg  arvalid; // @[ICache.scala 142:24]
  reg  rready; // @[ICache.scala 147:23]
  reg  tlb1_invalid; // @[ICache.scala 151:21]
  wire [31:0] _ar_addr_T_1 = {inst_pa[31:6],6'h0}; // @[Cat.scala 33:92]
  wire  _GEN_3078 = 6'h1 == va_line_addr ? meta_1_lru : meta_0_lru; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3079 = 6'h2 == va_line_addr ? meta_2_lru : _GEN_3078; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3080 = 6'h3 == va_line_addr ? meta_3_lru : _GEN_3079; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3081 = 6'h4 == va_line_addr ? meta_4_lru : _GEN_3080; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3082 = 6'h5 == va_line_addr ? meta_5_lru : _GEN_3081; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3083 = 6'h6 == va_line_addr ? meta_6_lru : _GEN_3082; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3084 = 6'h7 == va_line_addr ? meta_7_lru : _GEN_3083; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3085 = 6'h8 == va_line_addr ? meta_8_lru : _GEN_3084; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3086 = 6'h9 == va_line_addr ? meta_9_lru : _GEN_3085; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3087 = 6'ha == va_line_addr ? meta_10_lru : _GEN_3086; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3088 = 6'hb == va_line_addr ? meta_11_lru : _GEN_3087; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3089 = 6'hc == va_line_addr ? meta_12_lru : _GEN_3088; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3090 = 6'hd == va_line_addr ? meta_13_lru : _GEN_3089; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3091 = 6'he == va_line_addr ? meta_14_lru : _GEN_3090; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3092 = 6'hf == va_line_addr ? meta_15_lru : _GEN_3091; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3093 = 6'h10 == va_line_addr ? meta_16_lru : _GEN_3092; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3094 = 6'h11 == va_line_addr ? meta_17_lru : _GEN_3093; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3095 = 6'h12 == va_line_addr ? meta_18_lru : _GEN_3094; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3096 = 6'h13 == va_line_addr ? meta_19_lru : _GEN_3095; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3097 = 6'h14 == va_line_addr ? meta_20_lru : _GEN_3096; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3098 = 6'h15 == va_line_addr ? meta_21_lru : _GEN_3097; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3099 = 6'h16 == va_line_addr ? meta_22_lru : _GEN_3098; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3100 = 6'h17 == va_line_addr ? meta_23_lru : _GEN_3099; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3101 = 6'h18 == va_line_addr ? meta_24_lru : _GEN_3100; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3102 = 6'h19 == va_line_addr ? meta_25_lru : _GEN_3101; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3103 = 6'h1a == va_line_addr ? meta_26_lru : _GEN_3102; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3104 = 6'h1b == va_line_addr ? meta_27_lru : _GEN_3103; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3105 = 6'h1c == va_line_addr ? meta_28_lru : _GEN_3104; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3106 = 6'h1d == va_line_addr ? meta_29_lru : _GEN_3105; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3107 = 6'h1e == va_line_addr ? meta_30_lru : _GEN_3106; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3108 = 6'h1f == va_line_addr ? meta_31_lru : _GEN_3107; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3109 = 6'h20 == va_line_addr ? meta_32_lru : _GEN_3108; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3110 = 6'h21 == va_line_addr ? meta_33_lru : _GEN_3109; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3111 = 6'h22 == va_line_addr ? meta_34_lru : _GEN_3110; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3112 = 6'h23 == va_line_addr ? meta_35_lru : _GEN_3111; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3113 = 6'h24 == va_line_addr ? meta_36_lru : _GEN_3112; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3114 = 6'h25 == va_line_addr ? meta_37_lru : _GEN_3113; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3115 = 6'h26 == va_line_addr ? meta_38_lru : _GEN_3114; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3116 = 6'h27 == va_line_addr ? meta_39_lru : _GEN_3115; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3117 = 6'h28 == va_line_addr ? meta_40_lru : _GEN_3116; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3118 = 6'h29 == va_line_addr ? meta_41_lru : _GEN_3117; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3119 = 6'h2a == va_line_addr ? meta_42_lru : _GEN_3118; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3120 = 6'h2b == va_line_addr ? meta_43_lru : _GEN_3119; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3121 = 6'h2c == va_line_addr ? meta_44_lru : _GEN_3120; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3122 = 6'h2d == va_line_addr ? meta_45_lru : _GEN_3121; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3123 = 6'h2e == va_line_addr ? meta_46_lru : _GEN_3122; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3124 = 6'h2f == va_line_addr ? meta_47_lru : _GEN_3123; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3125 = 6'h30 == va_line_addr ? meta_48_lru : _GEN_3124; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3126 = 6'h31 == va_line_addr ? meta_49_lru : _GEN_3125; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3127 = 6'h32 == va_line_addr ? meta_50_lru : _GEN_3126; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3128 = 6'h33 == va_line_addr ? meta_51_lru : _GEN_3127; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3129 = 6'h34 == va_line_addr ? meta_52_lru : _GEN_3128; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3130 = 6'h35 == va_line_addr ? meta_53_lru : _GEN_3129; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3131 = 6'h36 == va_line_addr ? meta_54_lru : _GEN_3130; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3132 = 6'h37 == va_line_addr ? meta_55_lru : _GEN_3131; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3133 = 6'h38 == va_line_addr ? meta_56_lru : _GEN_3132; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3134 = 6'h39 == va_line_addr ? meta_57_lru : _GEN_3133; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3135 = 6'h3a == va_line_addr ? meta_58_lru : _GEN_3134; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3136 = 6'h3b == va_line_addr ? meta_59_lru : _GEN_3135; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3137 = 6'h3c == va_line_addr ? meta_60_lru : _GEN_3136; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3138 = 6'h3d == va_line_addr ? meta_61_lru : _GEN_3137; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3139 = 6'h3e == va_line_addr ? meta_62_lru : _GEN_3138; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3140 = 6'h3f == va_line_addr ? meta_63_lru : _GEN_3139; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3141 = 7'h40 == _GEN_13517 ? meta_64_lru : _GEN_3140; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3142 = 7'h41 == _GEN_13517 ? meta_65_lru : _GEN_3141; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3143 = 7'h42 == _GEN_13517 ? meta_66_lru : _GEN_3142; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3144 = 7'h43 == _GEN_13517 ? meta_67_lru : _GEN_3143; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3145 = 7'h44 == _GEN_13517 ? meta_68_lru : _GEN_3144; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3146 = 7'h45 == _GEN_13517 ? meta_69_lru : _GEN_3145; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3147 = 7'h46 == _GEN_13517 ? meta_70_lru : _GEN_3146; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3148 = 7'h47 == _GEN_13517 ? meta_71_lru : _GEN_3147; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3149 = 7'h48 == _GEN_13517 ? meta_72_lru : _GEN_3148; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3150 = 7'h49 == _GEN_13517 ? meta_73_lru : _GEN_3149; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3151 = 7'h4a == _GEN_13517 ? meta_74_lru : _GEN_3150; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3152 = 7'h4b == _GEN_13517 ? meta_75_lru : _GEN_3151; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3153 = 7'h4c == _GEN_13517 ? meta_76_lru : _GEN_3152; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3154 = 7'h4d == _GEN_13517 ? meta_77_lru : _GEN_3153; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3155 = 7'h4e == _GEN_13517 ? meta_78_lru : _GEN_3154; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3156 = 7'h4f == _GEN_13517 ? meta_79_lru : _GEN_3155; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3157 = 7'h50 == _GEN_13517 ? meta_80_lru : _GEN_3156; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3158 = 7'h51 == _GEN_13517 ? meta_81_lru : _GEN_3157; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3159 = 7'h52 == _GEN_13517 ? meta_82_lru : _GEN_3158; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3160 = 7'h53 == _GEN_13517 ? meta_83_lru : _GEN_3159; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3161 = 7'h54 == _GEN_13517 ? meta_84_lru : _GEN_3160; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3162 = 7'h55 == _GEN_13517 ? meta_85_lru : _GEN_3161; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3163 = 7'h56 == _GEN_13517 ? meta_86_lru : _GEN_3162; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3164 = 7'h57 == _GEN_13517 ? meta_87_lru : _GEN_3163; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3165 = 7'h58 == _GEN_13517 ? meta_88_lru : _GEN_3164; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3166 = 7'h59 == _GEN_13517 ? meta_89_lru : _GEN_3165; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3167 = 7'h5a == _GEN_13517 ? meta_90_lru : _GEN_3166; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3168 = 7'h5b == _GEN_13517 ? meta_91_lru : _GEN_3167; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3169 = 7'h5c == _GEN_13517 ? meta_92_lru : _GEN_3168; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3170 = 7'h5d == _GEN_13517 ? meta_93_lru : _GEN_3169; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3171 = 7'h5e == _GEN_13517 ? meta_94_lru : _GEN_3170; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3172 = 7'h5f == _GEN_13517 ? meta_95_lru : _GEN_3171; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3173 = 7'h60 == _GEN_13517 ? meta_96_lru : _GEN_3172; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3174 = 7'h61 == _GEN_13517 ? meta_97_lru : _GEN_3173; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3175 = 7'h62 == _GEN_13517 ? meta_98_lru : _GEN_3174; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3176 = 7'h63 == _GEN_13517 ? meta_99_lru : _GEN_3175; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3177 = 7'h64 == _GEN_13517 ? meta_100_lru : _GEN_3176; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3178 = 7'h65 == _GEN_13517 ? meta_101_lru : _GEN_3177; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3179 = 7'h66 == _GEN_13517 ? meta_102_lru : _GEN_3178; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3180 = 7'h67 == _GEN_13517 ? meta_103_lru : _GEN_3179; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3181 = 7'h68 == _GEN_13517 ? meta_104_lru : _GEN_3180; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3182 = 7'h69 == _GEN_13517 ? meta_105_lru : _GEN_3181; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3183 = 7'h6a == _GEN_13517 ? meta_106_lru : _GEN_3182; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3184 = 7'h6b == _GEN_13517 ? meta_107_lru : _GEN_3183; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3185 = 7'h6c == _GEN_13517 ? meta_108_lru : _GEN_3184; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3186 = 7'h6d == _GEN_13517 ? meta_109_lru : _GEN_3185; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3187 = 7'h6e == _GEN_13517 ? meta_110_lru : _GEN_3186; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3188 = 7'h6f == _GEN_13517 ? meta_111_lru : _GEN_3187; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3189 = 7'h70 == _GEN_13517 ? meta_112_lru : _GEN_3188; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3190 = 7'h71 == _GEN_13517 ? meta_113_lru : _GEN_3189; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3191 = 7'h72 == _GEN_13517 ? meta_114_lru : _GEN_3190; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3192 = 7'h73 == _GEN_13517 ? meta_115_lru : _GEN_3191; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3193 = 7'h74 == _GEN_13517 ? meta_116_lru : _GEN_3192; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3194 = 7'h75 == _GEN_13517 ? meta_117_lru : _GEN_3193; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3195 = 7'h76 == _GEN_13517 ? meta_118_lru : _GEN_3194; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3196 = 7'h77 == _GEN_13517 ? meta_119_lru : _GEN_3195; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3197 = 7'h78 == _GEN_13517 ? meta_120_lru : _GEN_3196; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3198 = 7'h79 == _GEN_13517 ? meta_121_lru : _GEN_3197; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3199 = 7'h7a == _GEN_13517 ? meta_122_lru : _GEN_3198; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3200 = 7'h7b == _GEN_13517 ? meta_123_lru : _GEN_3199; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3201 = 7'h7c == _GEN_13517 ? meta_124_lru : _GEN_3200; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3202 = 7'h7d == _GEN_13517 ? meta_125_lru : _GEN_3201; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3203 = 7'h7e == _GEN_13517 ? meta_126_lru : _GEN_3202; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3204 = 7'h7f == _GEN_13517 ? meta_127_lru : _GEN_3203; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3205 = 8'h80 == _GEN_13581 ? meta_128_lru : _GEN_3204; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3206 = 8'h81 == _GEN_13581 ? meta_129_lru : _GEN_3205; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3207 = 8'h82 == _GEN_13581 ? meta_130_lru : _GEN_3206; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3208 = 8'h83 == _GEN_13581 ? meta_131_lru : _GEN_3207; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3209 = 8'h84 == _GEN_13581 ? meta_132_lru : _GEN_3208; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3210 = 8'h85 == _GEN_13581 ? meta_133_lru : _GEN_3209; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3211 = 8'h86 == _GEN_13581 ? meta_134_lru : _GEN_3210; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3212 = 8'h87 == _GEN_13581 ? meta_135_lru : _GEN_3211; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3213 = 8'h88 == _GEN_13581 ? meta_136_lru : _GEN_3212; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3214 = 8'h89 == _GEN_13581 ? meta_137_lru : _GEN_3213; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3215 = 8'h8a == _GEN_13581 ? meta_138_lru : _GEN_3214; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3216 = 8'h8b == _GEN_13581 ? meta_139_lru : _GEN_3215; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3217 = 8'h8c == _GEN_13581 ? meta_140_lru : _GEN_3216; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3218 = 8'h8d == _GEN_13581 ? meta_141_lru : _GEN_3217; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3219 = 8'h8e == _GEN_13581 ? meta_142_lru : _GEN_3218; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3220 = 8'h8f == _GEN_13581 ? meta_143_lru : _GEN_3219; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3221 = 8'h90 == _GEN_13581 ? meta_144_lru : _GEN_3220; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3222 = 8'h91 == _GEN_13581 ? meta_145_lru : _GEN_3221; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3223 = 8'h92 == _GEN_13581 ? meta_146_lru : _GEN_3222; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3224 = 8'h93 == _GEN_13581 ? meta_147_lru : _GEN_3223; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3225 = 8'h94 == _GEN_13581 ? meta_148_lru : _GEN_3224; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3226 = 8'h95 == _GEN_13581 ? meta_149_lru : _GEN_3225; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3227 = 8'h96 == _GEN_13581 ? meta_150_lru : _GEN_3226; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3228 = 8'h97 == _GEN_13581 ? meta_151_lru : _GEN_3227; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3229 = 8'h98 == _GEN_13581 ? meta_152_lru : _GEN_3228; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3230 = 8'h99 == _GEN_13581 ? meta_153_lru : _GEN_3229; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3231 = 8'h9a == _GEN_13581 ? meta_154_lru : _GEN_3230; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3232 = 8'h9b == _GEN_13581 ? meta_155_lru : _GEN_3231; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3233 = 8'h9c == _GEN_13581 ? meta_156_lru : _GEN_3232; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3234 = 8'h9d == _GEN_13581 ? meta_157_lru : _GEN_3233; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3235 = 8'h9e == _GEN_13581 ? meta_158_lru : _GEN_3234; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3236 = 8'h9f == _GEN_13581 ? meta_159_lru : _GEN_3235; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3237 = 8'ha0 == _GEN_13581 ? meta_160_lru : _GEN_3236; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3238 = 8'ha1 == _GEN_13581 ? meta_161_lru : _GEN_3237; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3239 = 8'ha2 == _GEN_13581 ? meta_162_lru : _GEN_3238; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3240 = 8'ha3 == _GEN_13581 ? meta_163_lru : _GEN_3239; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3241 = 8'ha4 == _GEN_13581 ? meta_164_lru : _GEN_3240; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3242 = 8'ha5 == _GEN_13581 ? meta_165_lru : _GEN_3241; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3243 = 8'ha6 == _GEN_13581 ? meta_166_lru : _GEN_3242; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3244 = 8'ha7 == _GEN_13581 ? meta_167_lru : _GEN_3243; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3245 = 8'ha8 == _GEN_13581 ? meta_168_lru : _GEN_3244; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3246 = 8'ha9 == _GEN_13581 ? meta_169_lru : _GEN_3245; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3247 = 8'haa == _GEN_13581 ? meta_170_lru : _GEN_3246; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3248 = 8'hab == _GEN_13581 ? meta_171_lru : _GEN_3247; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3249 = 8'hac == _GEN_13581 ? meta_172_lru : _GEN_3248; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3250 = 8'had == _GEN_13581 ? meta_173_lru : _GEN_3249; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3251 = 8'hae == _GEN_13581 ? meta_174_lru : _GEN_3250; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3252 = 8'haf == _GEN_13581 ? meta_175_lru : _GEN_3251; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3253 = 8'hb0 == _GEN_13581 ? meta_176_lru : _GEN_3252; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3254 = 8'hb1 == _GEN_13581 ? meta_177_lru : _GEN_3253; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3255 = 8'hb2 == _GEN_13581 ? meta_178_lru : _GEN_3254; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3256 = 8'hb3 == _GEN_13581 ? meta_179_lru : _GEN_3255; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3257 = 8'hb4 == _GEN_13581 ? meta_180_lru : _GEN_3256; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3258 = 8'hb5 == _GEN_13581 ? meta_181_lru : _GEN_3257; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3259 = 8'hb6 == _GEN_13581 ? meta_182_lru : _GEN_3258; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3260 = 8'hb7 == _GEN_13581 ? meta_183_lru : _GEN_3259; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3261 = 8'hb8 == _GEN_13581 ? meta_184_lru : _GEN_3260; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3262 = 8'hb9 == _GEN_13581 ? meta_185_lru : _GEN_3261; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3263 = 8'hba == _GEN_13581 ? meta_186_lru : _GEN_3262; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3264 = 8'hbb == _GEN_13581 ? meta_187_lru : _GEN_3263; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3265 = 8'hbc == _GEN_13581 ? meta_188_lru : _GEN_3264; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3266 = 8'hbd == _GEN_13581 ? meta_189_lru : _GEN_3265; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3267 = 8'hbe == _GEN_13581 ? meta_190_lru : _GEN_3266; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3268 = 8'hbf == _GEN_13581 ? meta_191_lru : _GEN_3267; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3269 = 8'hc0 == _GEN_13581 ? meta_192_lru : _GEN_3268; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3270 = 8'hc1 == _GEN_13581 ? meta_193_lru : _GEN_3269; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3271 = 8'hc2 == _GEN_13581 ? meta_194_lru : _GEN_3270; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3272 = 8'hc3 == _GEN_13581 ? meta_195_lru : _GEN_3271; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3273 = 8'hc4 == _GEN_13581 ? meta_196_lru : _GEN_3272; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3274 = 8'hc5 == _GEN_13581 ? meta_197_lru : _GEN_3273; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3275 = 8'hc6 == _GEN_13581 ? meta_198_lru : _GEN_3274; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3276 = 8'hc7 == _GEN_13581 ? meta_199_lru : _GEN_3275; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3277 = 8'hc8 == _GEN_13581 ? meta_200_lru : _GEN_3276; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3278 = 8'hc9 == _GEN_13581 ? meta_201_lru : _GEN_3277; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3279 = 8'hca == _GEN_13581 ? meta_202_lru : _GEN_3278; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3280 = 8'hcb == _GEN_13581 ? meta_203_lru : _GEN_3279; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3281 = 8'hcc == _GEN_13581 ? meta_204_lru : _GEN_3280; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3282 = 8'hcd == _GEN_13581 ? meta_205_lru : _GEN_3281; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3283 = 8'hce == _GEN_13581 ? meta_206_lru : _GEN_3282; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3284 = 8'hcf == _GEN_13581 ? meta_207_lru : _GEN_3283; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3285 = 8'hd0 == _GEN_13581 ? meta_208_lru : _GEN_3284; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3286 = 8'hd1 == _GEN_13581 ? meta_209_lru : _GEN_3285; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3287 = 8'hd2 == _GEN_13581 ? meta_210_lru : _GEN_3286; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3288 = 8'hd3 == _GEN_13581 ? meta_211_lru : _GEN_3287; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3289 = 8'hd4 == _GEN_13581 ? meta_212_lru : _GEN_3288; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3290 = 8'hd5 == _GEN_13581 ? meta_213_lru : _GEN_3289; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3291 = 8'hd6 == _GEN_13581 ? meta_214_lru : _GEN_3290; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3292 = 8'hd7 == _GEN_13581 ? meta_215_lru : _GEN_3291; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3293 = 8'hd8 == _GEN_13581 ? meta_216_lru : _GEN_3292; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3294 = 8'hd9 == _GEN_13581 ? meta_217_lru : _GEN_3293; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3295 = 8'hda == _GEN_13581 ? meta_218_lru : _GEN_3294; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3296 = 8'hdb == _GEN_13581 ? meta_219_lru : _GEN_3295; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3297 = 8'hdc == _GEN_13581 ? meta_220_lru : _GEN_3296; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3298 = 8'hdd == _GEN_13581 ? meta_221_lru : _GEN_3297; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3299 = 8'hde == _GEN_13581 ? meta_222_lru : _GEN_3298; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3300 = 8'hdf == _GEN_13581 ? meta_223_lru : _GEN_3299; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3301 = 8'he0 == _GEN_13581 ? meta_224_lru : _GEN_3300; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3302 = 8'he1 == _GEN_13581 ? meta_225_lru : _GEN_3301; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3303 = 8'he2 == _GEN_13581 ? meta_226_lru : _GEN_3302; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3304 = 8'he3 == _GEN_13581 ? meta_227_lru : _GEN_3303; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3305 = 8'he4 == _GEN_13581 ? meta_228_lru : _GEN_3304; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3306 = 8'he5 == _GEN_13581 ? meta_229_lru : _GEN_3305; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3307 = 8'he6 == _GEN_13581 ? meta_230_lru : _GEN_3306; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3308 = 8'he7 == _GEN_13581 ? meta_231_lru : _GEN_3307; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3309 = 8'he8 == _GEN_13581 ? meta_232_lru : _GEN_3308; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3310 = 8'he9 == _GEN_13581 ? meta_233_lru : _GEN_3309; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3311 = 8'hea == _GEN_13581 ? meta_234_lru : _GEN_3310; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3312 = 8'heb == _GEN_13581 ? meta_235_lru : _GEN_3311; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3313 = 8'hec == _GEN_13581 ? meta_236_lru : _GEN_3312; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3314 = 8'hed == _GEN_13581 ? meta_237_lru : _GEN_3313; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3315 = 8'hee == _GEN_13581 ? meta_238_lru : _GEN_3314; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3316 = 8'hef == _GEN_13581 ? meta_239_lru : _GEN_3315; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3317 = 8'hf0 == _GEN_13581 ? meta_240_lru : _GEN_3316; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3318 = 8'hf1 == _GEN_13581 ? meta_241_lru : _GEN_3317; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3319 = 8'hf2 == _GEN_13581 ? meta_242_lru : _GEN_3318; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3320 = 8'hf3 == _GEN_13581 ? meta_243_lru : _GEN_3319; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3321 = 8'hf4 == _GEN_13581 ? meta_244_lru : _GEN_3320; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3322 = 8'hf5 == _GEN_13581 ? meta_245_lru : _GEN_3321; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3323 = 8'hf6 == _GEN_13581 ? meta_246_lru : _GEN_3322; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3324 = 8'hf7 == _GEN_13581 ? meta_247_lru : _GEN_3323; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3325 = 8'hf8 == _GEN_13581 ? meta_248_lru : _GEN_3324; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3326 = 8'hf9 == _GEN_13581 ? meta_249_lru : _GEN_3325; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3327 = 8'hfa == _GEN_13581 ? meta_250_lru : _GEN_3326; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3328 = 8'hfb == _GEN_13581 ? meta_251_lru : _GEN_3327; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3329 = 8'hfc == _GEN_13581 ? meta_252_lru : _GEN_3328; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3330 = 8'hfd == _GEN_13581 ? meta_253_lru : _GEN_3329; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3331 = 8'hfe == _GEN_13581 ? meta_254_lru : _GEN_3330; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3332 = 8'hff == _GEN_13581 ? meta_255_lru : _GEN_3331; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3333 = 9'h100 == _GEN_13709 ? meta_256_lru : _GEN_3332; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3334 = 9'h101 == _GEN_13709 ? meta_257_lru : _GEN_3333; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3335 = 9'h102 == _GEN_13709 ? meta_258_lru : _GEN_3334; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3336 = 9'h103 == _GEN_13709 ? meta_259_lru : _GEN_3335; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3337 = 9'h104 == _GEN_13709 ? meta_260_lru : _GEN_3336; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3338 = 9'h105 == _GEN_13709 ? meta_261_lru : _GEN_3337; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3339 = 9'h106 == _GEN_13709 ? meta_262_lru : _GEN_3338; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3340 = 9'h107 == _GEN_13709 ? meta_263_lru : _GEN_3339; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3341 = 9'h108 == _GEN_13709 ? meta_264_lru : _GEN_3340; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3342 = 9'h109 == _GEN_13709 ? meta_265_lru : _GEN_3341; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3343 = 9'h10a == _GEN_13709 ? meta_266_lru : _GEN_3342; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3344 = 9'h10b == _GEN_13709 ? meta_267_lru : _GEN_3343; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3345 = 9'h10c == _GEN_13709 ? meta_268_lru : _GEN_3344; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3346 = 9'h10d == _GEN_13709 ? meta_269_lru : _GEN_3345; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3347 = 9'h10e == _GEN_13709 ? meta_270_lru : _GEN_3346; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3348 = 9'h10f == _GEN_13709 ? meta_271_lru : _GEN_3347; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3349 = 9'h110 == _GEN_13709 ? meta_272_lru : _GEN_3348; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3350 = 9'h111 == _GEN_13709 ? meta_273_lru : _GEN_3349; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3351 = 9'h112 == _GEN_13709 ? meta_274_lru : _GEN_3350; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3352 = 9'h113 == _GEN_13709 ? meta_275_lru : _GEN_3351; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3353 = 9'h114 == _GEN_13709 ? meta_276_lru : _GEN_3352; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3354 = 9'h115 == _GEN_13709 ? meta_277_lru : _GEN_3353; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3355 = 9'h116 == _GEN_13709 ? meta_278_lru : _GEN_3354; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3356 = 9'h117 == _GEN_13709 ? meta_279_lru : _GEN_3355; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3357 = 9'h118 == _GEN_13709 ? meta_280_lru : _GEN_3356; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3358 = 9'h119 == _GEN_13709 ? meta_281_lru : _GEN_3357; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3359 = 9'h11a == _GEN_13709 ? meta_282_lru : _GEN_3358; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3360 = 9'h11b == _GEN_13709 ? meta_283_lru : _GEN_3359; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3361 = 9'h11c == _GEN_13709 ? meta_284_lru : _GEN_3360; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3362 = 9'h11d == _GEN_13709 ? meta_285_lru : _GEN_3361; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3363 = 9'h11e == _GEN_13709 ? meta_286_lru : _GEN_3362; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3364 = 9'h11f == _GEN_13709 ? meta_287_lru : _GEN_3363; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3365 = 9'h120 == _GEN_13709 ? meta_288_lru : _GEN_3364; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3366 = 9'h121 == _GEN_13709 ? meta_289_lru : _GEN_3365; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3367 = 9'h122 == _GEN_13709 ? meta_290_lru : _GEN_3366; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3368 = 9'h123 == _GEN_13709 ? meta_291_lru : _GEN_3367; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3369 = 9'h124 == _GEN_13709 ? meta_292_lru : _GEN_3368; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3370 = 9'h125 == _GEN_13709 ? meta_293_lru : _GEN_3369; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3371 = 9'h126 == _GEN_13709 ? meta_294_lru : _GEN_3370; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3372 = 9'h127 == _GEN_13709 ? meta_295_lru : _GEN_3371; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3373 = 9'h128 == _GEN_13709 ? meta_296_lru : _GEN_3372; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3374 = 9'h129 == _GEN_13709 ? meta_297_lru : _GEN_3373; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3375 = 9'h12a == _GEN_13709 ? meta_298_lru : _GEN_3374; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3376 = 9'h12b == _GEN_13709 ? meta_299_lru : _GEN_3375; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3377 = 9'h12c == _GEN_13709 ? meta_300_lru : _GEN_3376; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3378 = 9'h12d == _GEN_13709 ? meta_301_lru : _GEN_3377; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3379 = 9'h12e == _GEN_13709 ? meta_302_lru : _GEN_3378; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3380 = 9'h12f == _GEN_13709 ? meta_303_lru : _GEN_3379; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3381 = 9'h130 == _GEN_13709 ? meta_304_lru : _GEN_3380; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3382 = 9'h131 == _GEN_13709 ? meta_305_lru : _GEN_3381; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3383 = 9'h132 == _GEN_13709 ? meta_306_lru : _GEN_3382; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3384 = 9'h133 == _GEN_13709 ? meta_307_lru : _GEN_3383; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3385 = 9'h134 == _GEN_13709 ? meta_308_lru : _GEN_3384; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3386 = 9'h135 == _GEN_13709 ? meta_309_lru : _GEN_3385; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3387 = 9'h136 == _GEN_13709 ? meta_310_lru : _GEN_3386; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3388 = 9'h137 == _GEN_13709 ? meta_311_lru : _GEN_3387; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3389 = 9'h138 == _GEN_13709 ? meta_312_lru : _GEN_3388; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3390 = 9'h139 == _GEN_13709 ? meta_313_lru : _GEN_3389; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3391 = 9'h13a == _GEN_13709 ? meta_314_lru : _GEN_3390; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3392 = 9'h13b == _GEN_13709 ? meta_315_lru : _GEN_3391; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3393 = 9'h13c == _GEN_13709 ? meta_316_lru : _GEN_3392; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3394 = 9'h13d == _GEN_13709 ? meta_317_lru : _GEN_3393; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3395 = 9'h13e == _GEN_13709 ? meta_318_lru : _GEN_3394; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3396 = 9'h13f == _GEN_13709 ? meta_319_lru : _GEN_3395; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3397 = 9'h140 == _GEN_13709 ? meta_320_lru : _GEN_3396; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3398 = 9'h141 == _GEN_13709 ? meta_321_lru : _GEN_3397; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3399 = 9'h142 == _GEN_13709 ? meta_322_lru : _GEN_3398; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3400 = 9'h143 == _GEN_13709 ? meta_323_lru : _GEN_3399; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3401 = 9'h144 == _GEN_13709 ? meta_324_lru : _GEN_3400; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3402 = 9'h145 == _GEN_13709 ? meta_325_lru : _GEN_3401; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3403 = 9'h146 == _GEN_13709 ? meta_326_lru : _GEN_3402; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3404 = 9'h147 == _GEN_13709 ? meta_327_lru : _GEN_3403; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3405 = 9'h148 == _GEN_13709 ? meta_328_lru : _GEN_3404; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3406 = 9'h149 == _GEN_13709 ? meta_329_lru : _GEN_3405; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3407 = 9'h14a == _GEN_13709 ? meta_330_lru : _GEN_3406; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3408 = 9'h14b == _GEN_13709 ? meta_331_lru : _GEN_3407; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3409 = 9'h14c == _GEN_13709 ? meta_332_lru : _GEN_3408; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3410 = 9'h14d == _GEN_13709 ? meta_333_lru : _GEN_3409; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3411 = 9'h14e == _GEN_13709 ? meta_334_lru : _GEN_3410; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3412 = 9'h14f == _GEN_13709 ? meta_335_lru : _GEN_3411; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3413 = 9'h150 == _GEN_13709 ? meta_336_lru : _GEN_3412; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3414 = 9'h151 == _GEN_13709 ? meta_337_lru : _GEN_3413; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3415 = 9'h152 == _GEN_13709 ? meta_338_lru : _GEN_3414; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3416 = 9'h153 == _GEN_13709 ? meta_339_lru : _GEN_3415; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3417 = 9'h154 == _GEN_13709 ? meta_340_lru : _GEN_3416; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3418 = 9'h155 == _GEN_13709 ? meta_341_lru : _GEN_3417; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3419 = 9'h156 == _GEN_13709 ? meta_342_lru : _GEN_3418; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3420 = 9'h157 == _GEN_13709 ? meta_343_lru : _GEN_3419; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3421 = 9'h158 == _GEN_13709 ? meta_344_lru : _GEN_3420; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3422 = 9'h159 == _GEN_13709 ? meta_345_lru : _GEN_3421; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3423 = 9'h15a == _GEN_13709 ? meta_346_lru : _GEN_3422; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3424 = 9'h15b == _GEN_13709 ? meta_347_lru : _GEN_3423; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3425 = 9'h15c == _GEN_13709 ? meta_348_lru : _GEN_3424; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3426 = 9'h15d == _GEN_13709 ? meta_349_lru : _GEN_3425; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3427 = 9'h15e == _GEN_13709 ? meta_350_lru : _GEN_3426; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3428 = 9'h15f == _GEN_13709 ? meta_351_lru : _GEN_3427; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3429 = 9'h160 == _GEN_13709 ? meta_352_lru : _GEN_3428; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3430 = 9'h161 == _GEN_13709 ? meta_353_lru : _GEN_3429; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3431 = 9'h162 == _GEN_13709 ? meta_354_lru : _GEN_3430; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3432 = 9'h163 == _GEN_13709 ? meta_355_lru : _GEN_3431; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3433 = 9'h164 == _GEN_13709 ? meta_356_lru : _GEN_3432; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3434 = 9'h165 == _GEN_13709 ? meta_357_lru : _GEN_3433; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3435 = 9'h166 == _GEN_13709 ? meta_358_lru : _GEN_3434; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3436 = 9'h167 == _GEN_13709 ? meta_359_lru : _GEN_3435; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3437 = 9'h168 == _GEN_13709 ? meta_360_lru : _GEN_3436; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3438 = 9'h169 == _GEN_13709 ? meta_361_lru : _GEN_3437; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3439 = 9'h16a == _GEN_13709 ? meta_362_lru : _GEN_3438; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3440 = 9'h16b == _GEN_13709 ? meta_363_lru : _GEN_3439; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3441 = 9'h16c == _GEN_13709 ? meta_364_lru : _GEN_3440; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3442 = 9'h16d == _GEN_13709 ? meta_365_lru : _GEN_3441; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3443 = 9'h16e == _GEN_13709 ? meta_366_lru : _GEN_3442; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3444 = 9'h16f == _GEN_13709 ? meta_367_lru : _GEN_3443; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3445 = 9'h170 == _GEN_13709 ? meta_368_lru : _GEN_3444; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3446 = 9'h171 == _GEN_13709 ? meta_369_lru : _GEN_3445; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3447 = 9'h172 == _GEN_13709 ? meta_370_lru : _GEN_3446; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3448 = 9'h173 == _GEN_13709 ? meta_371_lru : _GEN_3447; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3449 = 9'h174 == _GEN_13709 ? meta_372_lru : _GEN_3448; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3450 = 9'h175 == _GEN_13709 ? meta_373_lru : _GEN_3449; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3451 = 9'h176 == _GEN_13709 ? meta_374_lru : _GEN_3450; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3452 = 9'h177 == _GEN_13709 ? meta_375_lru : _GEN_3451; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3453 = 9'h178 == _GEN_13709 ? meta_376_lru : _GEN_3452; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3454 = 9'h179 == _GEN_13709 ? meta_377_lru : _GEN_3453; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3455 = 9'h17a == _GEN_13709 ? meta_378_lru : _GEN_3454; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3456 = 9'h17b == _GEN_13709 ? meta_379_lru : _GEN_3455; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3457 = 9'h17c == _GEN_13709 ? meta_380_lru : _GEN_3456; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3458 = 9'h17d == _GEN_13709 ? meta_381_lru : _GEN_3457; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3459 = 9'h17e == _GEN_13709 ? meta_382_lru : _GEN_3458; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3460 = 9'h17f == _GEN_13709 ? meta_383_lru : _GEN_3459; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3461 = 9'h180 == _GEN_13709 ? meta_384_lru : _GEN_3460; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3462 = 9'h181 == _GEN_13709 ? meta_385_lru : _GEN_3461; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3463 = 9'h182 == _GEN_13709 ? meta_386_lru : _GEN_3462; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3464 = 9'h183 == _GEN_13709 ? meta_387_lru : _GEN_3463; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3465 = 9'h184 == _GEN_13709 ? meta_388_lru : _GEN_3464; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3466 = 9'h185 == _GEN_13709 ? meta_389_lru : _GEN_3465; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3467 = 9'h186 == _GEN_13709 ? meta_390_lru : _GEN_3466; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3468 = 9'h187 == _GEN_13709 ? meta_391_lru : _GEN_3467; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3469 = 9'h188 == _GEN_13709 ? meta_392_lru : _GEN_3468; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3470 = 9'h189 == _GEN_13709 ? meta_393_lru : _GEN_3469; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3471 = 9'h18a == _GEN_13709 ? meta_394_lru : _GEN_3470; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3472 = 9'h18b == _GEN_13709 ? meta_395_lru : _GEN_3471; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3473 = 9'h18c == _GEN_13709 ? meta_396_lru : _GEN_3472; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3474 = 9'h18d == _GEN_13709 ? meta_397_lru : _GEN_3473; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3475 = 9'h18e == _GEN_13709 ? meta_398_lru : _GEN_3474; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3476 = 9'h18f == _GEN_13709 ? meta_399_lru : _GEN_3475; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3477 = 9'h190 == _GEN_13709 ? meta_400_lru : _GEN_3476; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3478 = 9'h191 == _GEN_13709 ? meta_401_lru : _GEN_3477; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3479 = 9'h192 == _GEN_13709 ? meta_402_lru : _GEN_3478; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3480 = 9'h193 == _GEN_13709 ? meta_403_lru : _GEN_3479; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3481 = 9'h194 == _GEN_13709 ? meta_404_lru : _GEN_3480; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3482 = 9'h195 == _GEN_13709 ? meta_405_lru : _GEN_3481; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3483 = 9'h196 == _GEN_13709 ? meta_406_lru : _GEN_3482; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3484 = 9'h197 == _GEN_13709 ? meta_407_lru : _GEN_3483; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3485 = 9'h198 == _GEN_13709 ? meta_408_lru : _GEN_3484; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3486 = 9'h199 == _GEN_13709 ? meta_409_lru : _GEN_3485; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3487 = 9'h19a == _GEN_13709 ? meta_410_lru : _GEN_3486; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3488 = 9'h19b == _GEN_13709 ? meta_411_lru : _GEN_3487; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3489 = 9'h19c == _GEN_13709 ? meta_412_lru : _GEN_3488; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3490 = 9'h19d == _GEN_13709 ? meta_413_lru : _GEN_3489; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3491 = 9'h19e == _GEN_13709 ? meta_414_lru : _GEN_3490; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3492 = 9'h19f == _GEN_13709 ? meta_415_lru : _GEN_3491; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3493 = 9'h1a0 == _GEN_13709 ? meta_416_lru : _GEN_3492; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3494 = 9'h1a1 == _GEN_13709 ? meta_417_lru : _GEN_3493; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3495 = 9'h1a2 == _GEN_13709 ? meta_418_lru : _GEN_3494; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3496 = 9'h1a3 == _GEN_13709 ? meta_419_lru : _GEN_3495; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3497 = 9'h1a4 == _GEN_13709 ? meta_420_lru : _GEN_3496; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3498 = 9'h1a5 == _GEN_13709 ? meta_421_lru : _GEN_3497; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3499 = 9'h1a6 == _GEN_13709 ? meta_422_lru : _GEN_3498; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3500 = 9'h1a7 == _GEN_13709 ? meta_423_lru : _GEN_3499; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3501 = 9'h1a8 == _GEN_13709 ? meta_424_lru : _GEN_3500; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3502 = 9'h1a9 == _GEN_13709 ? meta_425_lru : _GEN_3501; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3503 = 9'h1aa == _GEN_13709 ? meta_426_lru : _GEN_3502; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3504 = 9'h1ab == _GEN_13709 ? meta_427_lru : _GEN_3503; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3505 = 9'h1ac == _GEN_13709 ? meta_428_lru : _GEN_3504; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3506 = 9'h1ad == _GEN_13709 ? meta_429_lru : _GEN_3505; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3507 = 9'h1ae == _GEN_13709 ? meta_430_lru : _GEN_3506; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3508 = 9'h1af == _GEN_13709 ? meta_431_lru : _GEN_3507; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3509 = 9'h1b0 == _GEN_13709 ? meta_432_lru : _GEN_3508; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3510 = 9'h1b1 == _GEN_13709 ? meta_433_lru : _GEN_3509; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3511 = 9'h1b2 == _GEN_13709 ? meta_434_lru : _GEN_3510; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3512 = 9'h1b3 == _GEN_13709 ? meta_435_lru : _GEN_3511; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3513 = 9'h1b4 == _GEN_13709 ? meta_436_lru : _GEN_3512; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3514 = 9'h1b5 == _GEN_13709 ? meta_437_lru : _GEN_3513; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3515 = 9'h1b6 == _GEN_13709 ? meta_438_lru : _GEN_3514; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3516 = 9'h1b7 == _GEN_13709 ? meta_439_lru : _GEN_3515; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3517 = 9'h1b8 == _GEN_13709 ? meta_440_lru : _GEN_3516; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3518 = 9'h1b9 == _GEN_13709 ? meta_441_lru : _GEN_3517; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3519 = 9'h1ba == _GEN_13709 ? meta_442_lru : _GEN_3518; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3520 = 9'h1bb == _GEN_13709 ? meta_443_lru : _GEN_3519; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3521 = 9'h1bc == _GEN_13709 ? meta_444_lru : _GEN_3520; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3522 = 9'h1bd == _GEN_13709 ? meta_445_lru : _GEN_3521; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3523 = 9'h1be == _GEN_13709 ? meta_446_lru : _GEN_3522; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3524 = 9'h1bf == _GEN_13709 ? meta_447_lru : _GEN_3523; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3525 = 9'h1c0 == _GEN_13709 ? meta_448_lru : _GEN_3524; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3526 = 9'h1c1 == _GEN_13709 ? meta_449_lru : _GEN_3525; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3527 = 9'h1c2 == _GEN_13709 ? meta_450_lru : _GEN_3526; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3528 = 9'h1c3 == _GEN_13709 ? meta_451_lru : _GEN_3527; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3529 = 9'h1c4 == _GEN_13709 ? meta_452_lru : _GEN_3528; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3530 = 9'h1c5 == _GEN_13709 ? meta_453_lru : _GEN_3529; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3531 = 9'h1c6 == _GEN_13709 ? meta_454_lru : _GEN_3530; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3532 = 9'h1c7 == _GEN_13709 ? meta_455_lru : _GEN_3531; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3533 = 9'h1c8 == _GEN_13709 ? meta_456_lru : _GEN_3532; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3534 = 9'h1c9 == _GEN_13709 ? meta_457_lru : _GEN_3533; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3535 = 9'h1ca == _GEN_13709 ? meta_458_lru : _GEN_3534; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3536 = 9'h1cb == _GEN_13709 ? meta_459_lru : _GEN_3535; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3537 = 9'h1cc == _GEN_13709 ? meta_460_lru : _GEN_3536; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3538 = 9'h1cd == _GEN_13709 ? meta_461_lru : _GEN_3537; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3539 = 9'h1ce == _GEN_13709 ? meta_462_lru : _GEN_3538; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3540 = 9'h1cf == _GEN_13709 ? meta_463_lru : _GEN_3539; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3541 = 9'h1d0 == _GEN_13709 ? meta_464_lru : _GEN_3540; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3542 = 9'h1d1 == _GEN_13709 ? meta_465_lru : _GEN_3541; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3543 = 9'h1d2 == _GEN_13709 ? meta_466_lru : _GEN_3542; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3544 = 9'h1d3 == _GEN_13709 ? meta_467_lru : _GEN_3543; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3545 = 9'h1d4 == _GEN_13709 ? meta_468_lru : _GEN_3544; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3546 = 9'h1d5 == _GEN_13709 ? meta_469_lru : _GEN_3545; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3547 = 9'h1d6 == _GEN_13709 ? meta_470_lru : _GEN_3546; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3548 = 9'h1d7 == _GEN_13709 ? meta_471_lru : _GEN_3547; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3549 = 9'h1d8 == _GEN_13709 ? meta_472_lru : _GEN_3548; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3550 = 9'h1d9 == _GEN_13709 ? meta_473_lru : _GEN_3549; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3551 = 9'h1da == _GEN_13709 ? meta_474_lru : _GEN_3550; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3552 = 9'h1db == _GEN_13709 ? meta_475_lru : _GEN_3551; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3553 = 9'h1dc == _GEN_13709 ? meta_476_lru : _GEN_3552; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3554 = 9'h1dd == _GEN_13709 ? meta_477_lru : _GEN_3553; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3555 = 9'h1de == _GEN_13709 ? meta_478_lru : _GEN_3554; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3556 = 9'h1df == _GEN_13709 ? meta_479_lru : _GEN_3555; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3557 = 9'h1e0 == _GEN_13709 ? meta_480_lru : _GEN_3556; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3558 = 9'h1e1 == _GEN_13709 ? meta_481_lru : _GEN_3557; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3559 = 9'h1e2 == _GEN_13709 ? meta_482_lru : _GEN_3558; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3560 = 9'h1e3 == _GEN_13709 ? meta_483_lru : _GEN_3559; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3561 = 9'h1e4 == _GEN_13709 ? meta_484_lru : _GEN_3560; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3562 = 9'h1e5 == _GEN_13709 ? meta_485_lru : _GEN_3561; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3563 = 9'h1e6 == _GEN_13709 ? meta_486_lru : _GEN_3562; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3564 = 9'h1e7 == _GEN_13709 ? meta_487_lru : _GEN_3563; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3565 = 9'h1e8 == _GEN_13709 ? meta_488_lru : _GEN_3564; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3566 = 9'h1e9 == _GEN_13709 ? meta_489_lru : _GEN_3565; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3567 = 9'h1ea == _GEN_13709 ? meta_490_lru : _GEN_3566; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3568 = 9'h1eb == _GEN_13709 ? meta_491_lru : _GEN_3567; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3569 = 9'h1ec == _GEN_13709 ? meta_492_lru : _GEN_3568; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3570 = 9'h1ed == _GEN_13709 ? meta_493_lru : _GEN_3569; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3571 = 9'h1ee == _GEN_13709 ? meta_494_lru : _GEN_3570; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3572 = 9'h1ef == _GEN_13709 ? meta_495_lru : _GEN_3571; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3573 = 9'h1f0 == _GEN_13709 ? meta_496_lru : _GEN_3572; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3574 = 9'h1f1 == _GEN_13709 ? meta_497_lru : _GEN_3573; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3575 = 9'h1f2 == _GEN_13709 ? meta_498_lru : _GEN_3574; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3576 = 9'h1f3 == _GEN_13709 ? meta_499_lru : _GEN_3575; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3577 = 9'h1f4 == _GEN_13709 ? meta_500_lru : _GEN_3576; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3578 = 9'h1f5 == _GEN_13709 ? meta_501_lru : _GEN_3577; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3579 = 9'h1f6 == _GEN_13709 ? meta_502_lru : _GEN_3578; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3580 = 9'h1f7 == _GEN_13709 ? meta_503_lru : _GEN_3579; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3581 = 9'h1f8 == _GEN_13709 ? meta_504_lru : _GEN_3580; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3582 = 9'h1f9 == _GEN_13709 ? meta_505_lru : _GEN_3581; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3583 = 9'h1fa == _GEN_13709 ? meta_506_lru : _GEN_3582; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3584 = 9'h1fb == _GEN_13709 ? meta_507_lru : _GEN_3583; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3585 = 9'h1fc == _GEN_13709 ? meta_508_lru : _GEN_3584; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3586 = 9'h1fd == _GEN_13709 ? meta_509_lru : _GEN_3585; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3587 = 9'h1fe == _GEN_13709 ? meta_510_lru : _GEN_3586; // @[ICache.scala 183:{60,60}]
  wire  _GEN_3588 = 9'h1ff == _GEN_13709 ? meta_511_lru : _GEN_3587; // @[ICache.scala 183:{60,60}]
  wire [7:0] _GEN_3589 = ~_GEN_3588 ? 8'hf : data_wen_0; // @[ICache.scala 183:{60,60} 66:30]
  wire [7:0] _GEN_3590 = _GEN_3588 ? 8'hf : data_wen_1; // @[ICache.scala 183:{60,60} 66:30]
  wire  _GEN_15758 = ~_GEN_3588; // @[ICache.scala 184:{60,60} 67:30]
  wire  _GEN_3591 = ~_GEN_3588 | tag_wen_0; // @[ICache.scala 184:{60,60} 67:30]
  wire  _GEN_3592 = _GEN_3588 | tag_wen_1; // @[ICache.scala 184:{60,60} 67:30]
  wire  _GEN_3593 = 6'h0 == va_line_addr & _GEN_15758 | _GEN_2053; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3594 = 6'h0 == va_line_addr & _GEN_3588 | _GEN_2565; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3595 = 6'h1 == va_line_addr & _GEN_15758 | _GEN_2054; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3596 = 6'h1 == va_line_addr & _GEN_3588 | _GEN_2566; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3597 = 6'h2 == va_line_addr & _GEN_15758 | _GEN_2055; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3598 = 6'h2 == va_line_addr & _GEN_3588 | _GEN_2567; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3599 = 6'h3 == va_line_addr & _GEN_15758 | _GEN_2056; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3600 = 6'h3 == va_line_addr & _GEN_3588 | _GEN_2568; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3601 = 6'h4 == va_line_addr & _GEN_15758 | _GEN_2057; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3602 = 6'h4 == va_line_addr & _GEN_3588 | _GEN_2569; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3603 = 6'h5 == va_line_addr & _GEN_15758 | _GEN_2058; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3604 = 6'h5 == va_line_addr & _GEN_3588 | _GEN_2570; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3605 = 6'h6 == va_line_addr & _GEN_15758 | _GEN_2059; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3606 = 6'h6 == va_line_addr & _GEN_3588 | _GEN_2571; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3607 = 6'h7 == va_line_addr & _GEN_15758 | _GEN_2060; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3608 = 6'h7 == va_line_addr & _GEN_3588 | _GEN_2572; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3609 = 6'h8 == va_line_addr & _GEN_15758 | _GEN_2061; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3610 = 6'h8 == va_line_addr & _GEN_3588 | _GEN_2573; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3611 = 6'h9 == va_line_addr & _GEN_15758 | _GEN_2062; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3612 = 6'h9 == va_line_addr & _GEN_3588 | _GEN_2574; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3613 = 6'ha == va_line_addr & _GEN_15758 | _GEN_2063; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3614 = 6'ha == va_line_addr & _GEN_3588 | _GEN_2575; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3615 = 6'hb == va_line_addr & _GEN_15758 | _GEN_2064; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3616 = 6'hb == va_line_addr & _GEN_3588 | _GEN_2576; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3617 = 6'hc == va_line_addr & _GEN_15758 | _GEN_2065; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3618 = 6'hc == va_line_addr & _GEN_3588 | _GEN_2577; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3619 = 6'hd == va_line_addr & _GEN_15758 | _GEN_2066; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3620 = 6'hd == va_line_addr & _GEN_3588 | _GEN_2578; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3621 = 6'he == va_line_addr & _GEN_15758 | _GEN_2067; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3622 = 6'he == va_line_addr & _GEN_3588 | _GEN_2579; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3623 = 6'hf == va_line_addr & _GEN_15758 | _GEN_2068; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3624 = 6'hf == va_line_addr & _GEN_3588 | _GEN_2580; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3625 = 6'h10 == va_line_addr & _GEN_15758 | _GEN_2069; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3626 = 6'h10 == va_line_addr & _GEN_3588 | _GEN_2581; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3627 = 6'h11 == va_line_addr & _GEN_15758 | _GEN_2070; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3628 = 6'h11 == va_line_addr & _GEN_3588 | _GEN_2582; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3629 = 6'h12 == va_line_addr & _GEN_15758 | _GEN_2071; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3630 = 6'h12 == va_line_addr & _GEN_3588 | _GEN_2583; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3631 = 6'h13 == va_line_addr & _GEN_15758 | _GEN_2072; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3632 = 6'h13 == va_line_addr & _GEN_3588 | _GEN_2584; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3633 = 6'h14 == va_line_addr & _GEN_15758 | _GEN_2073; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3634 = 6'h14 == va_line_addr & _GEN_3588 | _GEN_2585; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3635 = 6'h15 == va_line_addr & _GEN_15758 | _GEN_2074; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3636 = 6'h15 == va_line_addr & _GEN_3588 | _GEN_2586; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3637 = 6'h16 == va_line_addr & _GEN_15758 | _GEN_2075; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3638 = 6'h16 == va_line_addr & _GEN_3588 | _GEN_2587; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3639 = 6'h17 == va_line_addr & _GEN_15758 | _GEN_2076; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3640 = 6'h17 == va_line_addr & _GEN_3588 | _GEN_2588; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3641 = 6'h18 == va_line_addr & _GEN_15758 | _GEN_2077; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3642 = 6'h18 == va_line_addr & _GEN_3588 | _GEN_2589; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3643 = 6'h19 == va_line_addr & _GEN_15758 | _GEN_2078; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3644 = 6'h19 == va_line_addr & _GEN_3588 | _GEN_2590; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3645 = 6'h1a == va_line_addr & _GEN_15758 | _GEN_2079; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3646 = 6'h1a == va_line_addr & _GEN_3588 | _GEN_2591; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3647 = 6'h1b == va_line_addr & _GEN_15758 | _GEN_2080; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3648 = 6'h1b == va_line_addr & _GEN_3588 | _GEN_2592; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3649 = 6'h1c == va_line_addr & _GEN_15758 | _GEN_2081; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3650 = 6'h1c == va_line_addr & _GEN_3588 | _GEN_2593; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3651 = 6'h1d == va_line_addr & _GEN_15758 | _GEN_2082; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3652 = 6'h1d == va_line_addr & _GEN_3588 | _GEN_2594; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3653 = 6'h1e == va_line_addr & _GEN_15758 | _GEN_2083; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3654 = 6'h1e == va_line_addr & _GEN_3588 | _GEN_2595; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3655 = 6'h1f == va_line_addr & _GEN_15758 | _GEN_2084; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3656 = 6'h1f == va_line_addr & _GEN_3588 | _GEN_2596; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3657 = 6'h20 == va_line_addr & _GEN_15758 | _GEN_2085; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3658 = 6'h20 == va_line_addr & _GEN_3588 | _GEN_2597; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3659 = 6'h21 == va_line_addr & _GEN_15758 | _GEN_2086; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3660 = 6'h21 == va_line_addr & _GEN_3588 | _GEN_2598; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3661 = 6'h22 == va_line_addr & _GEN_15758 | _GEN_2087; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3662 = 6'h22 == va_line_addr & _GEN_3588 | _GEN_2599; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3663 = 6'h23 == va_line_addr & _GEN_15758 | _GEN_2088; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3664 = 6'h23 == va_line_addr & _GEN_3588 | _GEN_2600; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3665 = 6'h24 == va_line_addr & _GEN_15758 | _GEN_2089; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3666 = 6'h24 == va_line_addr & _GEN_3588 | _GEN_2601; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3667 = 6'h25 == va_line_addr & _GEN_15758 | _GEN_2090; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3668 = 6'h25 == va_line_addr & _GEN_3588 | _GEN_2602; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3669 = 6'h26 == va_line_addr & _GEN_15758 | _GEN_2091; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3670 = 6'h26 == va_line_addr & _GEN_3588 | _GEN_2603; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3671 = 6'h27 == va_line_addr & _GEN_15758 | _GEN_2092; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3672 = 6'h27 == va_line_addr & _GEN_3588 | _GEN_2604; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3673 = 6'h28 == va_line_addr & _GEN_15758 | _GEN_2093; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3674 = 6'h28 == va_line_addr & _GEN_3588 | _GEN_2605; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3675 = 6'h29 == va_line_addr & _GEN_15758 | _GEN_2094; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3676 = 6'h29 == va_line_addr & _GEN_3588 | _GEN_2606; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3677 = 6'h2a == va_line_addr & _GEN_15758 | _GEN_2095; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3678 = 6'h2a == va_line_addr & _GEN_3588 | _GEN_2607; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3679 = 6'h2b == va_line_addr & _GEN_15758 | _GEN_2096; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3680 = 6'h2b == va_line_addr & _GEN_3588 | _GEN_2608; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3681 = 6'h2c == va_line_addr & _GEN_15758 | _GEN_2097; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3682 = 6'h2c == va_line_addr & _GEN_3588 | _GEN_2609; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3683 = 6'h2d == va_line_addr & _GEN_15758 | _GEN_2098; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3684 = 6'h2d == va_line_addr & _GEN_3588 | _GEN_2610; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3685 = 6'h2e == va_line_addr & _GEN_15758 | _GEN_2099; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3686 = 6'h2e == va_line_addr & _GEN_3588 | _GEN_2611; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3687 = 6'h2f == va_line_addr & _GEN_15758 | _GEN_2100; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3688 = 6'h2f == va_line_addr & _GEN_3588 | _GEN_2612; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3689 = 6'h30 == va_line_addr & _GEN_15758 | _GEN_2101; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3690 = 6'h30 == va_line_addr & _GEN_3588 | _GEN_2613; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3691 = 6'h31 == va_line_addr & _GEN_15758 | _GEN_2102; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3692 = 6'h31 == va_line_addr & _GEN_3588 | _GEN_2614; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3693 = 6'h32 == va_line_addr & _GEN_15758 | _GEN_2103; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3694 = 6'h32 == va_line_addr & _GEN_3588 | _GEN_2615; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3695 = 6'h33 == va_line_addr & _GEN_15758 | _GEN_2104; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3696 = 6'h33 == va_line_addr & _GEN_3588 | _GEN_2616; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3697 = 6'h34 == va_line_addr & _GEN_15758 | _GEN_2105; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3698 = 6'h34 == va_line_addr & _GEN_3588 | _GEN_2617; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3699 = 6'h35 == va_line_addr & _GEN_15758 | _GEN_2106; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3700 = 6'h35 == va_line_addr & _GEN_3588 | _GEN_2618; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3701 = 6'h36 == va_line_addr & _GEN_15758 | _GEN_2107; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3702 = 6'h36 == va_line_addr & _GEN_3588 | _GEN_2619; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3703 = 6'h37 == va_line_addr & _GEN_15758 | _GEN_2108; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3704 = 6'h37 == va_line_addr & _GEN_3588 | _GEN_2620; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3705 = 6'h38 == va_line_addr & _GEN_15758 | _GEN_2109; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3706 = 6'h38 == va_line_addr & _GEN_3588 | _GEN_2621; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3707 = 6'h39 == va_line_addr & _GEN_15758 | _GEN_2110; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3708 = 6'h39 == va_line_addr & _GEN_3588 | _GEN_2622; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3709 = 6'h3a == va_line_addr & _GEN_15758 | _GEN_2111; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3710 = 6'h3a == va_line_addr & _GEN_3588 | _GEN_2623; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3711 = 6'h3b == va_line_addr & _GEN_15758 | _GEN_2112; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3712 = 6'h3b == va_line_addr & _GEN_3588 | _GEN_2624; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3713 = 6'h3c == va_line_addr & _GEN_15758 | _GEN_2113; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3714 = 6'h3c == va_line_addr & _GEN_3588 | _GEN_2625; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3715 = 6'h3d == va_line_addr & _GEN_15758 | _GEN_2114; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3716 = 6'h3d == va_line_addr & _GEN_3588 | _GEN_2626; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3717 = 6'h3e == va_line_addr & _GEN_15758 | _GEN_2115; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3718 = 6'h3e == va_line_addr & _GEN_3588 | _GEN_2627; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3719 = 6'h3f == va_line_addr & _GEN_15758 | _GEN_2116; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3720 = 6'h3f == va_line_addr & _GEN_3588 | _GEN_2628; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3721 = 7'h40 == _GEN_13517 & _GEN_15758 | _GEN_2117; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3722 = 7'h40 == _GEN_13517 & _GEN_3588 | _GEN_2629; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3723 = 7'h41 == _GEN_13517 & _GEN_15758 | _GEN_2118; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3724 = 7'h41 == _GEN_13517 & _GEN_3588 | _GEN_2630; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3725 = 7'h42 == _GEN_13517 & _GEN_15758 | _GEN_2119; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3726 = 7'h42 == _GEN_13517 & _GEN_3588 | _GEN_2631; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3727 = 7'h43 == _GEN_13517 & _GEN_15758 | _GEN_2120; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3728 = 7'h43 == _GEN_13517 & _GEN_3588 | _GEN_2632; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3729 = 7'h44 == _GEN_13517 & _GEN_15758 | _GEN_2121; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3730 = 7'h44 == _GEN_13517 & _GEN_3588 | _GEN_2633; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3731 = 7'h45 == _GEN_13517 & _GEN_15758 | _GEN_2122; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3732 = 7'h45 == _GEN_13517 & _GEN_3588 | _GEN_2634; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3733 = 7'h46 == _GEN_13517 & _GEN_15758 | _GEN_2123; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3734 = 7'h46 == _GEN_13517 & _GEN_3588 | _GEN_2635; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3735 = 7'h47 == _GEN_13517 & _GEN_15758 | _GEN_2124; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3736 = 7'h47 == _GEN_13517 & _GEN_3588 | _GEN_2636; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3737 = 7'h48 == _GEN_13517 & _GEN_15758 | _GEN_2125; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3738 = 7'h48 == _GEN_13517 & _GEN_3588 | _GEN_2637; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3739 = 7'h49 == _GEN_13517 & _GEN_15758 | _GEN_2126; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3740 = 7'h49 == _GEN_13517 & _GEN_3588 | _GEN_2638; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3741 = 7'h4a == _GEN_13517 & _GEN_15758 | _GEN_2127; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3742 = 7'h4a == _GEN_13517 & _GEN_3588 | _GEN_2639; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3743 = 7'h4b == _GEN_13517 & _GEN_15758 | _GEN_2128; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3744 = 7'h4b == _GEN_13517 & _GEN_3588 | _GEN_2640; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3745 = 7'h4c == _GEN_13517 & _GEN_15758 | _GEN_2129; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3746 = 7'h4c == _GEN_13517 & _GEN_3588 | _GEN_2641; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3747 = 7'h4d == _GEN_13517 & _GEN_15758 | _GEN_2130; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3748 = 7'h4d == _GEN_13517 & _GEN_3588 | _GEN_2642; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3749 = 7'h4e == _GEN_13517 & _GEN_15758 | _GEN_2131; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3750 = 7'h4e == _GEN_13517 & _GEN_3588 | _GEN_2643; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3751 = 7'h4f == _GEN_13517 & _GEN_15758 | _GEN_2132; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3752 = 7'h4f == _GEN_13517 & _GEN_3588 | _GEN_2644; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3753 = 7'h50 == _GEN_13517 & _GEN_15758 | _GEN_2133; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3754 = 7'h50 == _GEN_13517 & _GEN_3588 | _GEN_2645; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3755 = 7'h51 == _GEN_13517 & _GEN_15758 | _GEN_2134; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3756 = 7'h51 == _GEN_13517 & _GEN_3588 | _GEN_2646; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3757 = 7'h52 == _GEN_13517 & _GEN_15758 | _GEN_2135; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3758 = 7'h52 == _GEN_13517 & _GEN_3588 | _GEN_2647; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3759 = 7'h53 == _GEN_13517 & _GEN_15758 | _GEN_2136; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3760 = 7'h53 == _GEN_13517 & _GEN_3588 | _GEN_2648; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3761 = 7'h54 == _GEN_13517 & _GEN_15758 | _GEN_2137; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3762 = 7'h54 == _GEN_13517 & _GEN_3588 | _GEN_2649; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3763 = 7'h55 == _GEN_13517 & _GEN_15758 | _GEN_2138; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3764 = 7'h55 == _GEN_13517 & _GEN_3588 | _GEN_2650; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3765 = 7'h56 == _GEN_13517 & _GEN_15758 | _GEN_2139; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3766 = 7'h56 == _GEN_13517 & _GEN_3588 | _GEN_2651; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3767 = 7'h57 == _GEN_13517 & _GEN_15758 | _GEN_2140; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3768 = 7'h57 == _GEN_13517 & _GEN_3588 | _GEN_2652; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3769 = 7'h58 == _GEN_13517 & _GEN_15758 | _GEN_2141; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3770 = 7'h58 == _GEN_13517 & _GEN_3588 | _GEN_2653; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3771 = 7'h59 == _GEN_13517 & _GEN_15758 | _GEN_2142; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3772 = 7'h59 == _GEN_13517 & _GEN_3588 | _GEN_2654; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3773 = 7'h5a == _GEN_13517 & _GEN_15758 | _GEN_2143; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3774 = 7'h5a == _GEN_13517 & _GEN_3588 | _GEN_2655; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3775 = 7'h5b == _GEN_13517 & _GEN_15758 | _GEN_2144; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3776 = 7'h5b == _GEN_13517 & _GEN_3588 | _GEN_2656; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3777 = 7'h5c == _GEN_13517 & _GEN_15758 | _GEN_2145; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3778 = 7'h5c == _GEN_13517 & _GEN_3588 | _GEN_2657; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3779 = 7'h5d == _GEN_13517 & _GEN_15758 | _GEN_2146; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3780 = 7'h5d == _GEN_13517 & _GEN_3588 | _GEN_2658; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3781 = 7'h5e == _GEN_13517 & _GEN_15758 | _GEN_2147; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3782 = 7'h5e == _GEN_13517 & _GEN_3588 | _GEN_2659; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3783 = 7'h5f == _GEN_13517 & _GEN_15758 | _GEN_2148; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3784 = 7'h5f == _GEN_13517 & _GEN_3588 | _GEN_2660; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3785 = 7'h60 == _GEN_13517 & _GEN_15758 | _GEN_2149; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3786 = 7'h60 == _GEN_13517 & _GEN_3588 | _GEN_2661; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3787 = 7'h61 == _GEN_13517 & _GEN_15758 | _GEN_2150; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3788 = 7'h61 == _GEN_13517 & _GEN_3588 | _GEN_2662; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3789 = 7'h62 == _GEN_13517 & _GEN_15758 | _GEN_2151; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3790 = 7'h62 == _GEN_13517 & _GEN_3588 | _GEN_2663; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3791 = 7'h63 == _GEN_13517 & _GEN_15758 | _GEN_2152; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3792 = 7'h63 == _GEN_13517 & _GEN_3588 | _GEN_2664; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3793 = 7'h64 == _GEN_13517 & _GEN_15758 | _GEN_2153; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3794 = 7'h64 == _GEN_13517 & _GEN_3588 | _GEN_2665; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3795 = 7'h65 == _GEN_13517 & _GEN_15758 | _GEN_2154; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3796 = 7'h65 == _GEN_13517 & _GEN_3588 | _GEN_2666; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3797 = 7'h66 == _GEN_13517 & _GEN_15758 | _GEN_2155; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3798 = 7'h66 == _GEN_13517 & _GEN_3588 | _GEN_2667; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3799 = 7'h67 == _GEN_13517 & _GEN_15758 | _GEN_2156; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3800 = 7'h67 == _GEN_13517 & _GEN_3588 | _GEN_2668; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3801 = 7'h68 == _GEN_13517 & _GEN_15758 | _GEN_2157; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3802 = 7'h68 == _GEN_13517 & _GEN_3588 | _GEN_2669; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3803 = 7'h69 == _GEN_13517 & _GEN_15758 | _GEN_2158; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3804 = 7'h69 == _GEN_13517 & _GEN_3588 | _GEN_2670; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3805 = 7'h6a == _GEN_13517 & _GEN_15758 | _GEN_2159; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3806 = 7'h6a == _GEN_13517 & _GEN_3588 | _GEN_2671; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3807 = 7'h6b == _GEN_13517 & _GEN_15758 | _GEN_2160; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3808 = 7'h6b == _GEN_13517 & _GEN_3588 | _GEN_2672; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3809 = 7'h6c == _GEN_13517 & _GEN_15758 | _GEN_2161; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3810 = 7'h6c == _GEN_13517 & _GEN_3588 | _GEN_2673; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3811 = 7'h6d == _GEN_13517 & _GEN_15758 | _GEN_2162; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3812 = 7'h6d == _GEN_13517 & _GEN_3588 | _GEN_2674; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3813 = 7'h6e == _GEN_13517 & _GEN_15758 | _GEN_2163; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3814 = 7'h6e == _GEN_13517 & _GEN_3588 | _GEN_2675; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3815 = 7'h6f == _GEN_13517 & _GEN_15758 | _GEN_2164; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3816 = 7'h6f == _GEN_13517 & _GEN_3588 | _GEN_2676; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3817 = 7'h70 == _GEN_13517 & _GEN_15758 | _GEN_2165; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3818 = 7'h70 == _GEN_13517 & _GEN_3588 | _GEN_2677; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3819 = 7'h71 == _GEN_13517 & _GEN_15758 | _GEN_2166; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3820 = 7'h71 == _GEN_13517 & _GEN_3588 | _GEN_2678; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3821 = 7'h72 == _GEN_13517 & _GEN_15758 | _GEN_2167; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3822 = 7'h72 == _GEN_13517 & _GEN_3588 | _GEN_2679; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3823 = 7'h73 == _GEN_13517 & _GEN_15758 | _GEN_2168; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3824 = 7'h73 == _GEN_13517 & _GEN_3588 | _GEN_2680; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3825 = 7'h74 == _GEN_13517 & _GEN_15758 | _GEN_2169; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3826 = 7'h74 == _GEN_13517 & _GEN_3588 | _GEN_2681; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3827 = 7'h75 == _GEN_13517 & _GEN_15758 | _GEN_2170; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3828 = 7'h75 == _GEN_13517 & _GEN_3588 | _GEN_2682; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3829 = 7'h76 == _GEN_13517 & _GEN_15758 | _GEN_2171; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3830 = 7'h76 == _GEN_13517 & _GEN_3588 | _GEN_2683; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3831 = 7'h77 == _GEN_13517 & _GEN_15758 | _GEN_2172; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3832 = 7'h77 == _GEN_13517 & _GEN_3588 | _GEN_2684; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3833 = 7'h78 == _GEN_13517 & _GEN_15758 | _GEN_2173; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3834 = 7'h78 == _GEN_13517 & _GEN_3588 | _GEN_2685; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3835 = 7'h79 == _GEN_13517 & _GEN_15758 | _GEN_2174; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3836 = 7'h79 == _GEN_13517 & _GEN_3588 | _GEN_2686; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3837 = 7'h7a == _GEN_13517 & _GEN_15758 | _GEN_2175; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3838 = 7'h7a == _GEN_13517 & _GEN_3588 | _GEN_2687; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3839 = 7'h7b == _GEN_13517 & _GEN_15758 | _GEN_2176; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3840 = 7'h7b == _GEN_13517 & _GEN_3588 | _GEN_2688; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3841 = 7'h7c == _GEN_13517 & _GEN_15758 | _GEN_2177; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3842 = 7'h7c == _GEN_13517 & _GEN_3588 | _GEN_2689; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3843 = 7'h7d == _GEN_13517 & _GEN_15758 | _GEN_2178; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3844 = 7'h7d == _GEN_13517 & _GEN_3588 | _GEN_2690; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3845 = 7'h7e == _GEN_13517 & _GEN_15758 | _GEN_2179; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3846 = 7'h7e == _GEN_13517 & _GEN_3588 | _GEN_2691; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3847 = 7'h7f == _GEN_13517 & _GEN_15758 | _GEN_2180; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3848 = 7'h7f == _GEN_13517 & _GEN_3588 | _GEN_2692; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3849 = 8'h80 == _GEN_13581 & _GEN_15758 | _GEN_2181; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3850 = 8'h80 == _GEN_13581 & _GEN_3588 | _GEN_2693; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3851 = 8'h81 == _GEN_13581 & _GEN_15758 | _GEN_2182; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3852 = 8'h81 == _GEN_13581 & _GEN_3588 | _GEN_2694; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3853 = 8'h82 == _GEN_13581 & _GEN_15758 | _GEN_2183; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3854 = 8'h82 == _GEN_13581 & _GEN_3588 | _GEN_2695; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3855 = 8'h83 == _GEN_13581 & _GEN_15758 | _GEN_2184; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3856 = 8'h83 == _GEN_13581 & _GEN_3588 | _GEN_2696; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3857 = 8'h84 == _GEN_13581 & _GEN_15758 | _GEN_2185; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3858 = 8'h84 == _GEN_13581 & _GEN_3588 | _GEN_2697; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3859 = 8'h85 == _GEN_13581 & _GEN_15758 | _GEN_2186; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3860 = 8'h85 == _GEN_13581 & _GEN_3588 | _GEN_2698; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3861 = 8'h86 == _GEN_13581 & _GEN_15758 | _GEN_2187; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3862 = 8'h86 == _GEN_13581 & _GEN_3588 | _GEN_2699; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3863 = 8'h87 == _GEN_13581 & _GEN_15758 | _GEN_2188; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3864 = 8'h87 == _GEN_13581 & _GEN_3588 | _GEN_2700; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3865 = 8'h88 == _GEN_13581 & _GEN_15758 | _GEN_2189; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3866 = 8'h88 == _GEN_13581 & _GEN_3588 | _GEN_2701; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3867 = 8'h89 == _GEN_13581 & _GEN_15758 | _GEN_2190; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3868 = 8'h89 == _GEN_13581 & _GEN_3588 | _GEN_2702; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3869 = 8'h8a == _GEN_13581 & _GEN_15758 | _GEN_2191; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3870 = 8'h8a == _GEN_13581 & _GEN_3588 | _GEN_2703; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3871 = 8'h8b == _GEN_13581 & _GEN_15758 | _GEN_2192; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3872 = 8'h8b == _GEN_13581 & _GEN_3588 | _GEN_2704; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3873 = 8'h8c == _GEN_13581 & _GEN_15758 | _GEN_2193; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3874 = 8'h8c == _GEN_13581 & _GEN_3588 | _GEN_2705; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3875 = 8'h8d == _GEN_13581 & _GEN_15758 | _GEN_2194; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3876 = 8'h8d == _GEN_13581 & _GEN_3588 | _GEN_2706; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3877 = 8'h8e == _GEN_13581 & _GEN_15758 | _GEN_2195; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3878 = 8'h8e == _GEN_13581 & _GEN_3588 | _GEN_2707; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3879 = 8'h8f == _GEN_13581 & _GEN_15758 | _GEN_2196; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3880 = 8'h8f == _GEN_13581 & _GEN_3588 | _GEN_2708; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3881 = 8'h90 == _GEN_13581 & _GEN_15758 | _GEN_2197; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3882 = 8'h90 == _GEN_13581 & _GEN_3588 | _GEN_2709; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3883 = 8'h91 == _GEN_13581 & _GEN_15758 | _GEN_2198; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3884 = 8'h91 == _GEN_13581 & _GEN_3588 | _GEN_2710; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3885 = 8'h92 == _GEN_13581 & _GEN_15758 | _GEN_2199; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3886 = 8'h92 == _GEN_13581 & _GEN_3588 | _GEN_2711; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3887 = 8'h93 == _GEN_13581 & _GEN_15758 | _GEN_2200; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3888 = 8'h93 == _GEN_13581 & _GEN_3588 | _GEN_2712; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3889 = 8'h94 == _GEN_13581 & _GEN_15758 | _GEN_2201; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3890 = 8'h94 == _GEN_13581 & _GEN_3588 | _GEN_2713; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3891 = 8'h95 == _GEN_13581 & _GEN_15758 | _GEN_2202; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3892 = 8'h95 == _GEN_13581 & _GEN_3588 | _GEN_2714; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3893 = 8'h96 == _GEN_13581 & _GEN_15758 | _GEN_2203; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3894 = 8'h96 == _GEN_13581 & _GEN_3588 | _GEN_2715; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3895 = 8'h97 == _GEN_13581 & _GEN_15758 | _GEN_2204; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3896 = 8'h97 == _GEN_13581 & _GEN_3588 | _GEN_2716; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3897 = 8'h98 == _GEN_13581 & _GEN_15758 | _GEN_2205; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3898 = 8'h98 == _GEN_13581 & _GEN_3588 | _GEN_2717; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3899 = 8'h99 == _GEN_13581 & _GEN_15758 | _GEN_2206; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3900 = 8'h99 == _GEN_13581 & _GEN_3588 | _GEN_2718; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3901 = 8'h9a == _GEN_13581 & _GEN_15758 | _GEN_2207; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3902 = 8'h9a == _GEN_13581 & _GEN_3588 | _GEN_2719; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3903 = 8'h9b == _GEN_13581 & _GEN_15758 | _GEN_2208; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3904 = 8'h9b == _GEN_13581 & _GEN_3588 | _GEN_2720; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3905 = 8'h9c == _GEN_13581 & _GEN_15758 | _GEN_2209; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3906 = 8'h9c == _GEN_13581 & _GEN_3588 | _GEN_2721; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3907 = 8'h9d == _GEN_13581 & _GEN_15758 | _GEN_2210; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3908 = 8'h9d == _GEN_13581 & _GEN_3588 | _GEN_2722; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3909 = 8'h9e == _GEN_13581 & _GEN_15758 | _GEN_2211; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3910 = 8'h9e == _GEN_13581 & _GEN_3588 | _GEN_2723; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3911 = 8'h9f == _GEN_13581 & _GEN_15758 | _GEN_2212; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3912 = 8'h9f == _GEN_13581 & _GEN_3588 | _GEN_2724; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3913 = 8'ha0 == _GEN_13581 & _GEN_15758 | _GEN_2213; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3914 = 8'ha0 == _GEN_13581 & _GEN_3588 | _GEN_2725; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3915 = 8'ha1 == _GEN_13581 & _GEN_15758 | _GEN_2214; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3916 = 8'ha1 == _GEN_13581 & _GEN_3588 | _GEN_2726; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3917 = 8'ha2 == _GEN_13581 & _GEN_15758 | _GEN_2215; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3918 = 8'ha2 == _GEN_13581 & _GEN_3588 | _GEN_2727; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3919 = 8'ha3 == _GEN_13581 & _GEN_15758 | _GEN_2216; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3920 = 8'ha3 == _GEN_13581 & _GEN_3588 | _GEN_2728; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3921 = 8'ha4 == _GEN_13581 & _GEN_15758 | _GEN_2217; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3922 = 8'ha4 == _GEN_13581 & _GEN_3588 | _GEN_2729; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3923 = 8'ha5 == _GEN_13581 & _GEN_15758 | _GEN_2218; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3924 = 8'ha5 == _GEN_13581 & _GEN_3588 | _GEN_2730; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3925 = 8'ha6 == _GEN_13581 & _GEN_15758 | _GEN_2219; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3926 = 8'ha6 == _GEN_13581 & _GEN_3588 | _GEN_2731; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3927 = 8'ha7 == _GEN_13581 & _GEN_15758 | _GEN_2220; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3928 = 8'ha7 == _GEN_13581 & _GEN_3588 | _GEN_2732; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3929 = 8'ha8 == _GEN_13581 & _GEN_15758 | _GEN_2221; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3930 = 8'ha8 == _GEN_13581 & _GEN_3588 | _GEN_2733; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3931 = 8'ha9 == _GEN_13581 & _GEN_15758 | _GEN_2222; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3932 = 8'ha9 == _GEN_13581 & _GEN_3588 | _GEN_2734; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3933 = 8'haa == _GEN_13581 & _GEN_15758 | _GEN_2223; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3934 = 8'haa == _GEN_13581 & _GEN_3588 | _GEN_2735; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3935 = 8'hab == _GEN_13581 & _GEN_15758 | _GEN_2224; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3936 = 8'hab == _GEN_13581 & _GEN_3588 | _GEN_2736; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3937 = 8'hac == _GEN_13581 & _GEN_15758 | _GEN_2225; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3938 = 8'hac == _GEN_13581 & _GEN_3588 | _GEN_2737; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3939 = 8'had == _GEN_13581 & _GEN_15758 | _GEN_2226; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3940 = 8'had == _GEN_13581 & _GEN_3588 | _GEN_2738; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3941 = 8'hae == _GEN_13581 & _GEN_15758 | _GEN_2227; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3942 = 8'hae == _GEN_13581 & _GEN_3588 | _GEN_2739; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3943 = 8'haf == _GEN_13581 & _GEN_15758 | _GEN_2228; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3944 = 8'haf == _GEN_13581 & _GEN_3588 | _GEN_2740; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3945 = 8'hb0 == _GEN_13581 & _GEN_15758 | _GEN_2229; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3946 = 8'hb0 == _GEN_13581 & _GEN_3588 | _GEN_2741; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3947 = 8'hb1 == _GEN_13581 & _GEN_15758 | _GEN_2230; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3948 = 8'hb1 == _GEN_13581 & _GEN_3588 | _GEN_2742; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3949 = 8'hb2 == _GEN_13581 & _GEN_15758 | _GEN_2231; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3950 = 8'hb2 == _GEN_13581 & _GEN_3588 | _GEN_2743; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3951 = 8'hb3 == _GEN_13581 & _GEN_15758 | _GEN_2232; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3952 = 8'hb3 == _GEN_13581 & _GEN_3588 | _GEN_2744; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3953 = 8'hb4 == _GEN_13581 & _GEN_15758 | _GEN_2233; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3954 = 8'hb4 == _GEN_13581 & _GEN_3588 | _GEN_2745; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3955 = 8'hb5 == _GEN_13581 & _GEN_15758 | _GEN_2234; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3956 = 8'hb5 == _GEN_13581 & _GEN_3588 | _GEN_2746; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3957 = 8'hb6 == _GEN_13581 & _GEN_15758 | _GEN_2235; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3958 = 8'hb6 == _GEN_13581 & _GEN_3588 | _GEN_2747; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3959 = 8'hb7 == _GEN_13581 & _GEN_15758 | _GEN_2236; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3960 = 8'hb7 == _GEN_13581 & _GEN_3588 | _GEN_2748; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3961 = 8'hb8 == _GEN_13581 & _GEN_15758 | _GEN_2237; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3962 = 8'hb8 == _GEN_13581 & _GEN_3588 | _GEN_2749; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3963 = 8'hb9 == _GEN_13581 & _GEN_15758 | _GEN_2238; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3964 = 8'hb9 == _GEN_13581 & _GEN_3588 | _GEN_2750; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3965 = 8'hba == _GEN_13581 & _GEN_15758 | _GEN_2239; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3966 = 8'hba == _GEN_13581 & _GEN_3588 | _GEN_2751; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3967 = 8'hbb == _GEN_13581 & _GEN_15758 | _GEN_2240; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3968 = 8'hbb == _GEN_13581 & _GEN_3588 | _GEN_2752; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3969 = 8'hbc == _GEN_13581 & _GEN_15758 | _GEN_2241; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3970 = 8'hbc == _GEN_13581 & _GEN_3588 | _GEN_2753; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3971 = 8'hbd == _GEN_13581 & _GEN_15758 | _GEN_2242; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3972 = 8'hbd == _GEN_13581 & _GEN_3588 | _GEN_2754; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3973 = 8'hbe == _GEN_13581 & _GEN_15758 | _GEN_2243; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3974 = 8'hbe == _GEN_13581 & _GEN_3588 | _GEN_2755; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3975 = 8'hbf == _GEN_13581 & _GEN_15758 | _GEN_2244; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3976 = 8'hbf == _GEN_13581 & _GEN_3588 | _GEN_2756; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3977 = 8'hc0 == _GEN_13581 & _GEN_15758 | _GEN_2245; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3978 = 8'hc0 == _GEN_13581 & _GEN_3588 | _GEN_2757; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3979 = 8'hc1 == _GEN_13581 & _GEN_15758 | _GEN_2246; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3980 = 8'hc1 == _GEN_13581 & _GEN_3588 | _GEN_2758; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3981 = 8'hc2 == _GEN_13581 & _GEN_15758 | _GEN_2247; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3982 = 8'hc2 == _GEN_13581 & _GEN_3588 | _GEN_2759; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3983 = 8'hc3 == _GEN_13581 & _GEN_15758 | _GEN_2248; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3984 = 8'hc3 == _GEN_13581 & _GEN_3588 | _GEN_2760; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3985 = 8'hc4 == _GEN_13581 & _GEN_15758 | _GEN_2249; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3986 = 8'hc4 == _GEN_13581 & _GEN_3588 | _GEN_2761; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3987 = 8'hc5 == _GEN_13581 & _GEN_15758 | _GEN_2250; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3988 = 8'hc5 == _GEN_13581 & _GEN_3588 | _GEN_2762; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3989 = 8'hc6 == _GEN_13581 & _GEN_15758 | _GEN_2251; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3990 = 8'hc6 == _GEN_13581 & _GEN_3588 | _GEN_2763; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3991 = 8'hc7 == _GEN_13581 & _GEN_15758 | _GEN_2252; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3992 = 8'hc7 == _GEN_13581 & _GEN_3588 | _GEN_2764; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3993 = 8'hc8 == _GEN_13581 & _GEN_15758 | _GEN_2253; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3994 = 8'hc8 == _GEN_13581 & _GEN_3588 | _GEN_2765; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3995 = 8'hc9 == _GEN_13581 & _GEN_15758 | _GEN_2254; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3996 = 8'hc9 == _GEN_13581 & _GEN_3588 | _GEN_2766; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3997 = 8'hca == _GEN_13581 & _GEN_15758 | _GEN_2255; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3998 = 8'hca == _GEN_13581 & _GEN_3588 | _GEN_2767; // @[ICache.scala 186:{60,60}]
  wire  _GEN_3999 = 8'hcb == _GEN_13581 & _GEN_15758 | _GEN_2256; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4000 = 8'hcb == _GEN_13581 & _GEN_3588 | _GEN_2768; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4001 = 8'hcc == _GEN_13581 & _GEN_15758 | _GEN_2257; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4002 = 8'hcc == _GEN_13581 & _GEN_3588 | _GEN_2769; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4003 = 8'hcd == _GEN_13581 & _GEN_15758 | _GEN_2258; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4004 = 8'hcd == _GEN_13581 & _GEN_3588 | _GEN_2770; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4005 = 8'hce == _GEN_13581 & _GEN_15758 | _GEN_2259; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4006 = 8'hce == _GEN_13581 & _GEN_3588 | _GEN_2771; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4007 = 8'hcf == _GEN_13581 & _GEN_15758 | _GEN_2260; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4008 = 8'hcf == _GEN_13581 & _GEN_3588 | _GEN_2772; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4009 = 8'hd0 == _GEN_13581 & _GEN_15758 | _GEN_2261; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4010 = 8'hd0 == _GEN_13581 & _GEN_3588 | _GEN_2773; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4011 = 8'hd1 == _GEN_13581 & _GEN_15758 | _GEN_2262; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4012 = 8'hd1 == _GEN_13581 & _GEN_3588 | _GEN_2774; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4013 = 8'hd2 == _GEN_13581 & _GEN_15758 | _GEN_2263; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4014 = 8'hd2 == _GEN_13581 & _GEN_3588 | _GEN_2775; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4015 = 8'hd3 == _GEN_13581 & _GEN_15758 | _GEN_2264; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4016 = 8'hd3 == _GEN_13581 & _GEN_3588 | _GEN_2776; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4017 = 8'hd4 == _GEN_13581 & _GEN_15758 | _GEN_2265; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4018 = 8'hd4 == _GEN_13581 & _GEN_3588 | _GEN_2777; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4019 = 8'hd5 == _GEN_13581 & _GEN_15758 | _GEN_2266; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4020 = 8'hd5 == _GEN_13581 & _GEN_3588 | _GEN_2778; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4021 = 8'hd6 == _GEN_13581 & _GEN_15758 | _GEN_2267; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4022 = 8'hd6 == _GEN_13581 & _GEN_3588 | _GEN_2779; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4023 = 8'hd7 == _GEN_13581 & _GEN_15758 | _GEN_2268; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4024 = 8'hd7 == _GEN_13581 & _GEN_3588 | _GEN_2780; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4025 = 8'hd8 == _GEN_13581 & _GEN_15758 | _GEN_2269; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4026 = 8'hd8 == _GEN_13581 & _GEN_3588 | _GEN_2781; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4027 = 8'hd9 == _GEN_13581 & _GEN_15758 | _GEN_2270; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4028 = 8'hd9 == _GEN_13581 & _GEN_3588 | _GEN_2782; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4029 = 8'hda == _GEN_13581 & _GEN_15758 | _GEN_2271; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4030 = 8'hda == _GEN_13581 & _GEN_3588 | _GEN_2783; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4031 = 8'hdb == _GEN_13581 & _GEN_15758 | _GEN_2272; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4032 = 8'hdb == _GEN_13581 & _GEN_3588 | _GEN_2784; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4033 = 8'hdc == _GEN_13581 & _GEN_15758 | _GEN_2273; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4034 = 8'hdc == _GEN_13581 & _GEN_3588 | _GEN_2785; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4035 = 8'hdd == _GEN_13581 & _GEN_15758 | _GEN_2274; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4036 = 8'hdd == _GEN_13581 & _GEN_3588 | _GEN_2786; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4037 = 8'hde == _GEN_13581 & _GEN_15758 | _GEN_2275; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4038 = 8'hde == _GEN_13581 & _GEN_3588 | _GEN_2787; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4039 = 8'hdf == _GEN_13581 & _GEN_15758 | _GEN_2276; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4040 = 8'hdf == _GEN_13581 & _GEN_3588 | _GEN_2788; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4041 = 8'he0 == _GEN_13581 & _GEN_15758 | _GEN_2277; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4042 = 8'he0 == _GEN_13581 & _GEN_3588 | _GEN_2789; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4043 = 8'he1 == _GEN_13581 & _GEN_15758 | _GEN_2278; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4044 = 8'he1 == _GEN_13581 & _GEN_3588 | _GEN_2790; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4045 = 8'he2 == _GEN_13581 & _GEN_15758 | _GEN_2279; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4046 = 8'he2 == _GEN_13581 & _GEN_3588 | _GEN_2791; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4047 = 8'he3 == _GEN_13581 & _GEN_15758 | _GEN_2280; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4048 = 8'he3 == _GEN_13581 & _GEN_3588 | _GEN_2792; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4049 = 8'he4 == _GEN_13581 & _GEN_15758 | _GEN_2281; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4050 = 8'he4 == _GEN_13581 & _GEN_3588 | _GEN_2793; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4051 = 8'he5 == _GEN_13581 & _GEN_15758 | _GEN_2282; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4052 = 8'he5 == _GEN_13581 & _GEN_3588 | _GEN_2794; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4053 = 8'he6 == _GEN_13581 & _GEN_15758 | _GEN_2283; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4054 = 8'he6 == _GEN_13581 & _GEN_3588 | _GEN_2795; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4055 = 8'he7 == _GEN_13581 & _GEN_15758 | _GEN_2284; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4056 = 8'he7 == _GEN_13581 & _GEN_3588 | _GEN_2796; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4057 = 8'he8 == _GEN_13581 & _GEN_15758 | _GEN_2285; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4058 = 8'he8 == _GEN_13581 & _GEN_3588 | _GEN_2797; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4059 = 8'he9 == _GEN_13581 & _GEN_15758 | _GEN_2286; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4060 = 8'he9 == _GEN_13581 & _GEN_3588 | _GEN_2798; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4061 = 8'hea == _GEN_13581 & _GEN_15758 | _GEN_2287; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4062 = 8'hea == _GEN_13581 & _GEN_3588 | _GEN_2799; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4063 = 8'heb == _GEN_13581 & _GEN_15758 | _GEN_2288; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4064 = 8'heb == _GEN_13581 & _GEN_3588 | _GEN_2800; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4065 = 8'hec == _GEN_13581 & _GEN_15758 | _GEN_2289; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4066 = 8'hec == _GEN_13581 & _GEN_3588 | _GEN_2801; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4067 = 8'hed == _GEN_13581 & _GEN_15758 | _GEN_2290; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4068 = 8'hed == _GEN_13581 & _GEN_3588 | _GEN_2802; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4069 = 8'hee == _GEN_13581 & _GEN_15758 | _GEN_2291; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4070 = 8'hee == _GEN_13581 & _GEN_3588 | _GEN_2803; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4071 = 8'hef == _GEN_13581 & _GEN_15758 | _GEN_2292; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4072 = 8'hef == _GEN_13581 & _GEN_3588 | _GEN_2804; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4073 = 8'hf0 == _GEN_13581 & _GEN_15758 | _GEN_2293; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4074 = 8'hf0 == _GEN_13581 & _GEN_3588 | _GEN_2805; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4075 = 8'hf1 == _GEN_13581 & _GEN_15758 | _GEN_2294; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4076 = 8'hf1 == _GEN_13581 & _GEN_3588 | _GEN_2806; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4077 = 8'hf2 == _GEN_13581 & _GEN_15758 | _GEN_2295; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4078 = 8'hf2 == _GEN_13581 & _GEN_3588 | _GEN_2807; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4079 = 8'hf3 == _GEN_13581 & _GEN_15758 | _GEN_2296; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4080 = 8'hf3 == _GEN_13581 & _GEN_3588 | _GEN_2808; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4081 = 8'hf4 == _GEN_13581 & _GEN_15758 | _GEN_2297; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4082 = 8'hf4 == _GEN_13581 & _GEN_3588 | _GEN_2809; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4083 = 8'hf5 == _GEN_13581 & _GEN_15758 | _GEN_2298; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4084 = 8'hf5 == _GEN_13581 & _GEN_3588 | _GEN_2810; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4085 = 8'hf6 == _GEN_13581 & _GEN_15758 | _GEN_2299; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4086 = 8'hf6 == _GEN_13581 & _GEN_3588 | _GEN_2811; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4087 = 8'hf7 == _GEN_13581 & _GEN_15758 | _GEN_2300; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4088 = 8'hf7 == _GEN_13581 & _GEN_3588 | _GEN_2812; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4089 = 8'hf8 == _GEN_13581 & _GEN_15758 | _GEN_2301; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4090 = 8'hf8 == _GEN_13581 & _GEN_3588 | _GEN_2813; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4091 = 8'hf9 == _GEN_13581 & _GEN_15758 | _GEN_2302; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4092 = 8'hf9 == _GEN_13581 & _GEN_3588 | _GEN_2814; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4093 = 8'hfa == _GEN_13581 & _GEN_15758 | _GEN_2303; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4094 = 8'hfa == _GEN_13581 & _GEN_3588 | _GEN_2815; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4095 = 8'hfb == _GEN_13581 & _GEN_15758 | _GEN_2304; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4096 = 8'hfb == _GEN_13581 & _GEN_3588 | _GEN_2816; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4097 = 8'hfc == _GEN_13581 & _GEN_15758 | _GEN_2305; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4098 = 8'hfc == _GEN_13581 & _GEN_3588 | _GEN_2817; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4099 = 8'hfd == _GEN_13581 & _GEN_15758 | _GEN_2306; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4100 = 8'hfd == _GEN_13581 & _GEN_3588 | _GEN_2818; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4101 = 8'hfe == _GEN_13581 & _GEN_15758 | _GEN_2307; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4102 = 8'hfe == _GEN_13581 & _GEN_3588 | _GEN_2819; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4103 = 8'hff == _GEN_13581 & _GEN_15758 | _GEN_2308; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4104 = 8'hff == _GEN_13581 & _GEN_3588 | _GEN_2820; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4105 = 9'h100 == _GEN_13709 & _GEN_15758 | _GEN_2309; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4106 = 9'h100 == _GEN_13709 & _GEN_3588 | _GEN_2821; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4107 = 9'h101 == _GEN_13709 & _GEN_15758 | _GEN_2310; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4108 = 9'h101 == _GEN_13709 & _GEN_3588 | _GEN_2822; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4109 = 9'h102 == _GEN_13709 & _GEN_15758 | _GEN_2311; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4110 = 9'h102 == _GEN_13709 & _GEN_3588 | _GEN_2823; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4111 = 9'h103 == _GEN_13709 & _GEN_15758 | _GEN_2312; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4112 = 9'h103 == _GEN_13709 & _GEN_3588 | _GEN_2824; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4113 = 9'h104 == _GEN_13709 & _GEN_15758 | _GEN_2313; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4114 = 9'h104 == _GEN_13709 & _GEN_3588 | _GEN_2825; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4115 = 9'h105 == _GEN_13709 & _GEN_15758 | _GEN_2314; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4116 = 9'h105 == _GEN_13709 & _GEN_3588 | _GEN_2826; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4117 = 9'h106 == _GEN_13709 & _GEN_15758 | _GEN_2315; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4118 = 9'h106 == _GEN_13709 & _GEN_3588 | _GEN_2827; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4119 = 9'h107 == _GEN_13709 & _GEN_15758 | _GEN_2316; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4120 = 9'h107 == _GEN_13709 & _GEN_3588 | _GEN_2828; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4121 = 9'h108 == _GEN_13709 & _GEN_15758 | _GEN_2317; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4122 = 9'h108 == _GEN_13709 & _GEN_3588 | _GEN_2829; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4123 = 9'h109 == _GEN_13709 & _GEN_15758 | _GEN_2318; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4124 = 9'h109 == _GEN_13709 & _GEN_3588 | _GEN_2830; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4125 = 9'h10a == _GEN_13709 & _GEN_15758 | _GEN_2319; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4126 = 9'h10a == _GEN_13709 & _GEN_3588 | _GEN_2831; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4127 = 9'h10b == _GEN_13709 & _GEN_15758 | _GEN_2320; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4128 = 9'h10b == _GEN_13709 & _GEN_3588 | _GEN_2832; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4129 = 9'h10c == _GEN_13709 & _GEN_15758 | _GEN_2321; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4130 = 9'h10c == _GEN_13709 & _GEN_3588 | _GEN_2833; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4131 = 9'h10d == _GEN_13709 & _GEN_15758 | _GEN_2322; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4132 = 9'h10d == _GEN_13709 & _GEN_3588 | _GEN_2834; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4133 = 9'h10e == _GEN_13709 & _GEN_15758 | _GEN_2323; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4134 = 9'h10e == _GEN_13709 & _GEN_3588 | _GEN_2835; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4135 = 9'h10f == _GEN_13709 & _GEN_15758 | _GEN_2324; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4136 = 9'h10f == _GEN_13709 & _GEN_3588 | _GEN_2836; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4137 = 9'h110 == _GEN_13709 & _GEN_15758 | _GEN_2325; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4138 = 9'h110 == _GEN_13709 & _GEN_3588 | _GEN_2837; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4139 = 9'h111 == _GEN_13709 & _GEN_15758 | _GEN_2326; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4140 = 9'h111 == _GEN_13709 & _GEN_3588 | _GEN_2838; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4141 = 9'h112 == _GEN_13709 & _GEN_15758 | _GEN_2327; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4142 = 9'h112 == _GEN_13709 & _GEN_3588 | _GEN_2839; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4143 = 9'h113 == _GEN_13709 & _GEN_15758 | _GEN_2328; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4144 = 9'h113 == _GEN_13709 & _GEN_3588 | _GEN_2840; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4145 = 9'h114 == _GEN_13709 & _GEN_15758 | _GEN_2329; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4146 = 9'h114 == _GEN_13709 & _GEN_3588 | _GEN_2841; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4147 = 9'h115 == _GEN_13709 & _GEN_15758 | _GEN_2330; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4148 = 9'h115 == _GEN_13709 & _GEN_3588 | _GEN_2842; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4149 = 9'h116 == _GEN_13709 & _GEN_15758 | _GEN_2331; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4150 = 9'h116 == _GEN_13709 & _GEN_3588 | _GEN_2843; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4151 = 9'h117 == _GEN_13709 & _GEN_15758 | _GEN_2332; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4152 = 9'h117 == _GEN_13709 & _GEN_3588 | _GEN_2844; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4153 = 9'h118 == _GEN_13709 & _GEN_15758 | _GEN_2333; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4154 = 9'h118 == _GEN_13709 & _GEN_3588 | _GEN_2845; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4155 = 9'h119 == _GEN_13709 & _GEN_15758 | _GEN_2334; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4156 = 9'h119 == _GEN_13709 & _GEN_3588 | _GEN_2846; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4157 = 9'h11a == _GEN_13709 & _GEN_15758 | _GEN_2335; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4158 = 9'h11a == _GEN_13709 & _GEN_3588 | _GEN_2847; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4159 = 9'h11b == _GEN_13709 & _GEN_15758 | _GEN_2336; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4160 = 9'h11b == _GEN_13709 & _GEN_3588 | _GEN_2848; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4161 = 9'h11c == _GEN_13709 & _GEN_15758 | _GEN_2337; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4162 = 9'h11c == _GEN_13709 & _GEN_3588 | _GEN_2849; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4163 = 9'h11d == _GEN_13709 & _GEN_15758 | _GEN_2338; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4164 = 9'h11d == _GEN_13709 & _GEN_3588 | _GEN_2850; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4165 = 9'h11e == _GEN_13709 & _GEN_15758 | _GEN_2339; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4166 = 9'h11e == _GEN_13709 & _GEN_3588 | _GEN_2851; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4167 = 9'h11f == _GEN_13709 & _GEN_15758 | _GEN_2340; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4168 = 9'h11f == _GEN_13709 & _GEN_3588 | _GEN_2852; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4169 = 9'h120 == _GEN_13709 & _GEN_15758 | _GEN_2341; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4170 = 9'h120 == _GEN_13709 & _GEN_3588 | _GEN_2853; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4171 = 9'h121 == _GEN_13709 & _GEN_15758 | _GEN_2342; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4172 = 9'h121 == _GEN_13709 & _GEN_3588 | _GEN_2854; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4173 = 9'h122 == _GEN_13709 & _GEN_15758 | _GEN_2343; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4174 = 9'h122 == _GEN_13709 & _GEN_3588 | _GEN_2855; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4175 = 9'h123 == _GEN_13709 & _GEN_15758 | _GEN_2344; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4176 = 9'h123 == _GEN_13709 & _GEN_3588 | _GEN_2856; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4177 = 9'h124 == _GEN_13709 & _GEN_15758 | _GEN_2345; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4178 = 9'h124 == _GEN_13709 & _GEN_3588 | _GEN_2857; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4179 = 9'h125 == _GEN_13709 & _GEN_15758 | _GEN_2346; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4180 = 9'h125 == _GEN_13709 & _GEN_3588 | _GEN_2858; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4181 = 9'h126 == _GEN_13709 & _GEN_15758 | _GEN_2347; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4182 = 9'h126 == _GEN_13709 & _GEN_3588 | _GEN_2859; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4183 = 9'h127 == _GEN_13709 & _GEN_15758 | _GEN_2348; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4184 = 9'h127 == _GEN_13709 & _GEN_3588 | _GEN_2860; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4185 = 9'h128 == _GEN_13709 & _GEN_15758 | _GEN_2349; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4186 = 9'h128 == _GEN_13709 & _GEN_3588 | _GEN_2861; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4187 = 9'h129 == _GEN_13709 & _GEN_15758 | _GEN_2350; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4188 = 9'h129 == _GEN_13709 & _GEN_3588 | _GEN_2862; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4189 = 9'h12a == _GEN_13709 & _GEN_15758 | _GEN_2351; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4190 = 9'h12a == _GEN_13709 & _GEN_3588 | _GEN_2863; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4191 = 9'h12b == _GEN_13709 & _GEN_15758 | _GEN_2352; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4192 = 9'h12b == _GEN_13709 & _GEN_3588 | _GEN_2864; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4193 = 9'h12c == _GEN_13709 & _GEN_15758 | _GEN_2353; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4194 = 9'h12c == _GEN_13709 & _GEN_3588 | _GEN_2865; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4195 = 9'h12d == _GEN_13709 & _GEN_15758 | _GEN_2354; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4196 = 9'h12d == _GEN_13709 & _GEN_3588 | _GEN_2866; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4197 = 9'h12e == _GEN_13709 & _GEN_15758 | _GEN_2355; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4198 = 9'h12e == _GEN_13709 & _GEN_3588 | _GEN_2867; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4199 = 9'h12f == _GEN_13709 & _GEN_15758 | _GEN_2356; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4200 = 9'h12f == _GEN_13709 & _GEN_3588 | _GEN_2868; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4201 = 9'h130 == _GEN_13709 & _GEN_15758 | _GEN_2357; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4202 = 9'h130 == _GEN_13709 & _GEN_3588 | _GEN_2869; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4203 = 9'h131 == _GEN_13709 & _GEN_15758 | _GEN_2358; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4204 = 9'h131 == _GEN_13709 & _GEN_3588 | _GEN_2870; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4205 = 9'h132 == _GEN_13709 & _GEN_15758 | _GEN_2359; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4206 = 9'h132 == _GEN_13709 & _GEN_3588 | _GEN_2871; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4207 = 9'h133 == _GEN_13709 & _GEN_15758 | _GEN_2360; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4208 = 9'h133 == _GEN_13709 & _GEN_3588 | _GEN_2872; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4209 = 9'h134 == _GEN_13709 & _GEN_15758 | _GEN_2361; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4210 = 9'h134 == _GEN_13709 & _GEN_3588 | _GEN_2873; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4211 = 9'h135 == _GEN_13709 & _GEN_15758 | _GEN_2362; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4212 = 9'h135 == _GEN_13709 & _GEN_3588 | _GEN_2874; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4213 = 9'h136 == _GEN_13709 & _GEN_15758 | _GEN_2363; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4214 = 9'h136 == _GEN_13709 & _GEN_3588 | _GEN_2875; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4215 = 9'h137 == _GEN_13709 & _GEN_15758 | _GEN_2364; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4216 = 9'h137 == _GEN_13709 & _GEN_3588 | _GEN_2876; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4217 = 9'h138 == _GEN_13709 & _GEN_15758 | _GEN_2365; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4218 = 9'h138 == _GEN_13709 & _GEN_3588 | _GEN_2877; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4219 = 9'h139 == _GEN_13709 & _GEN_15758 | _GEN_2366; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4220 = 9'h139 == _GEN_13709 & _GEN_3588 | _GEN_2878; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4221 = 9'h13a == _GEN_13709 & _GEN_15758 | _GEN_2367; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4222 = 9'h13a == _GEN_13709 & _GEN_3588 | _GEN_2879; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4223 = 9'h13b == _GEN_13709 & _GEN_15758 | _GEN_2368; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4224 = 9'h13b == _GEN_13709 & _GEN_3588 | _GEN_2880; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4225 = 9'h13c == _GEN_13709 & _GEN_15758 | _GEN_2369; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4226 = 9'h13c == _GEN_13709 & _GEN_3588 | _GEN_2881; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4227 = 9'h13d == _GEN_13709 & _GEN_15758 | _GEN_2370; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4228 = 9'h13d == _GEN_13709 & _GEN_3588 | _GEN_2882; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4229 = 9'h13e == _GEN_13709 & _GEN_15758 | _GEN_2371; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4230 = 9'h13e == _GEN_13709 & _GEN_3588 | _GEN_2883; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4231 = 9'h13f == _GEN_13709 & _GEN_15758 | _GEN_2372; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4232 = 9'h13f == _GEN_13709 & _GEN_3588 | _GEN_2884; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4233 = 9'h140 == _GEN_13709 & _GEN_15758 | _GEN_2373; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4234 = 9'h140 == _GEN_13709 & _GEN_3588 | _GEN_2885; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4235 = 9'h141 == _GEN_13709 & _GEN_15758 | _GEN_2374; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4236 = 9'h141 == _GEN_13709 & _GEN_3588 | _GEN_2886; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4237 = 9'h142 == _GEN_13709 & _GEN_15758 | _GEN_2375; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4238 = 9'h142 == _GEN_13709 & _GEN_3588 | _GEN_2887; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4239 = 9'h143 == _GEN_13709 & _GEN_15758 | _GEN_2376; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4240 = 9'h143 == _GEN_13709 & _GEN_3588 | _GEN_2888; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4241 = 9'h144 == _GEN_13709 & _GEN_15758 | _GEN_2377; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4242 = 9'h144 == _GEN_13709 & _GEN_3588 | _GEN_2889; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4243 = 9'h145 == _GEN_13709 & _GEN_15758 | _GEN_2378; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4244 = 9'h145 == _GEN_13709 & _GEN_3588 | _GEN_2890; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4245 = 9'h146 == _GEN_13709 & _GEN_15758 | _GEN_2379; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4246 = 9'h146 == _GEN_13709 & _GEN_3588 | _GEN_2891; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4247 = 9'h147 == _GEN_13709 & _GEN_15758 | _GEN_2380; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4248 = 9'h147 == _GEN_13709 & _GEN_3588 | _GEN_2892; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4249 = 9'h148 == _GEN_13709 & _GEN_15758 | _GEN_2381; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4250 = 9'h148 == _GEN_13709 & _GEN_3588 | _GEN_2893; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4251 = 9'h149 == _GEN_13709 & _GEN_15758 | _GEN_2382; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4252 = 9'h149 == _GEN_13709 & _GEN_3588 | _GEN_2894; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4253 = 9'h14a == _GEN_13709 & _GEN_15758 | _GEN_2383; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4254 = 9'h14a == _GEN_13709 & _GEN_3588 | _GEN_2895; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4255 = 9'h14b == _GEN_13709 & _GEN_15758 | _GEN_2384; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4256 = 9'h14b == _GEN_13709 & _GEN_3588 | _GEN_2896; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4257 = 9'h14c == _GEN_13709 & _GEN_15758 | _GEN_2385; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4258 = 9'h14c == _GEN_13709 & _GEN_3588 | _GEN_2897; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4259 = 9'h14d == _GEN_13709 & _GEN_15758 | _GEN_2386; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4260 = 9'h14d == _GEN_13709 & _GEN_3588 | _GEN_2898; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4261 = 9'h14e == _GEN_13709 & _GEN_15758 | _GEN_2387; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4262 = 9'h14e == _GEN_13709 & _GEN_3588 | _GEN_2899; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4263 = 9'h14f == _GEN_13709 & _GEN_15758 | _GEN_2388; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4264 = 9'h14f == _GEN_13709 & _GEN_3588 | _GEN_2900; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4265 = 9'h150 == _GEN_13709 & _GEN_15758 | _GEN_2389; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4266 = 9'h150 == _GEN_13709 & _GEN_3588 | _GEN_2901; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4267 = 9'h151 == _GEN_13709 & _GEN_15758 | _GEN_2390; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4268 = 9'h151 == _GEN_13709 & _GEN_3588 | _GEN_2902; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4269 = 9'h152 == _GEN_13709 & _GEN_15758 | _GEN_2391; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4270 = 9'h152 == _GEN_13709 & _GEN_3588 | _GEN_2903; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4271 = 9'h153 == _GEN_13709 & _GEN_15758 | _GEN_2392; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4272 = 9'h153 == _GEN_13709 & _GEN_3588 | _GEN_2904; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4273 = 9'h154 == _GEN_13709 & _GEN_15758 | _GEN_2393; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4274 = 9'h154 == _GEN_13709 & _GEN_3588 | _GEN_2905; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4275 = 9'h155 == _GEN_13709 & _GEN_15758 | _GEN_2394; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4276 = 9'h155 == _GEN_13709 & _GEN_3588 | _GEN_2906; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4277 = 9'h156 == _GEN_13709 & _GEN_15758 | _GEN_2395; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4278 = 9'h156 == _GEN_13709 & _GEN_3588 | _GEN_2907; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4279 = 9'h157 == _GEN_13709 & _GEN_15758 | _GEN_2396; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4280 = 9'h157 == _GEN_13709 & _GEN_3588 | _GEN_2908; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4281 = 9'h158 == _GEN_13709 & _GEN_15758 | _GEN_2397; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4282 = 9'h158 == _GEN_13709 & _GEN_3588 | _GEN_2909; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4283 = 9'h159 == _GEN_13709 & _GEN_15758 | _GEN_2398; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4284 = 9'h159 == _GEN_13709 & _GEN_3588 | _GEN_2910; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4285 = 9'h15a == _GEN_13709 & _GEN_15758 | _GEN_2399; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4286 = 9'h15a == _GEN_13709 & _GEN_3588 | _GEN_2911; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4287 = 9'h15b == _GEN_13709 & _GEN_15758 | _GEN_2400; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4288 = 9'h15b == _GEN_13709 & _GEN_3588 | _GEN_2912; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4289 = 9'h15c == _GEN_13709 & _GEN_15758 | _GEN_2401; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4290 = 9'h15c == _GEN_13709 & _GEN_3588 | _GEN_2913; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4291 = 9'h15d == _GEN_13709 & _GEN_15758 | _GEN_2402; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4292 = 9'h15d == _GEN_13709 & _GEN_3588 | _GEN_2914; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4293 = 9'h15e == _GEN_13709 & _GEN_15758 | _GEN_2403; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4294 = 9'h15e == _GEN_13709 & _GEN_3588 | _GEN_2915; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4295 = 9'h15f == _GEN_13709 & _GEN_15758 | _GEN_2404; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4296 = 9'h15f == _GEN_13709 & _GEN_3588 | _GEN_2916; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4297 = 9'h160 == _GEN_13709 & _GEN_15758 | _GEN_2405; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4298 = 9'h160 == _GEN_13709 & _GEN_3588 | _GEN_2917; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4299 = 9'h161 == _GEN_13709 & _GEN_15758 | _GEN_2406; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4300 = 9'h161 == _GEN_13709 & _GEN_3588 | _GEN_2918; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4301 = 9'h162 == _GEN_13709 & _GEN_15758 | _GEN_2407; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4302 = 9'h162 == _GEN_13709 & _GEN_3588 | _GEN_2919; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4303 = 9'h163 == _GEN_13709 & _GEN_15758 | _GEN_2408; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4304 = 9'h163 == _GEN_13709 & _GEN_3588 | _GEN_2920; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4305 = 9'h164 == _GEN_13709 & _GEN_15758 | _GEN_2409; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4306 = 9'h164 == _GEN_13709 & _GEN_3588 | _GEN_2921; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4307 = 9'h165 == _GEN_13709 & _GEN_15758 | _GEN_2410; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4308 = 9'h165 == _GEN_13709 & _GEN_3588 | _GEN_2922; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4309 = 9'h166 == _GEN_13709 & _GEN_15758 | _GEN_2411; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4310 = 9'h166 == _GEN_13709 & _GEN_3588 | _GEN_2923; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4311 = 9'h167 == _GEN_13709 & _GEN_15758 | _GEN_2412; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4312 = 9'h167 == _GEN_13709 & _GEN_3588 | _GEN_2924; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4313 = 9'h168 == _GEN_13709 & _GEN_15758 | _GEN_2413; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4314 = 9'h168 == _GEN_13709 & _GEN_3588 | _GEN_2925; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4315 = 9'h169 == _GEN_13709 & _GEN_15758 | _GEN_2414; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4316 = 9'h169 == _GEN_13709 & _GEN_3588 | _GEN_2926; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4317 = 9'h16a == _GEN_13709 & _GEN_15758 | _GEN_2415; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4318 = 9'h16a == _GEN_13709 & _GEN_3588 | _GEN_2927; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4319 = 9'h16b == _GEN_13709 & _GEN_15758 | _GEN_2416; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4320 = 9'h16b == _GEN_13709 & _GEN_3588 | _GEN_2928; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4321 = 9'h16c == _GEN_13709 & _GEN_15758 | _GEN_2417; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4322 = 9'h16c == _GEN_13709 & _GEN_3588 | _GEN_2929; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4323 = 9'h16d == _GEN_13709 & _GEN_15758 | _GEN_2418; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4324 = 9'h16d == _GEN_13709 & _GEN_3588 | _GEN_2930; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4325 = 9'h16e == _GEN_13709 & _GEN_15758 | _GEN_2419; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4326 = 9'h16e == _GEN_13709 & _GEN_3588 | _GEN_2931; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4327 = 9'h16f == _GEN_13709 & _GEN_15758 | _GEN_2420; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4328 = 9'h16f == _GEN_13709 & _GEN_3588 | _GEN_2932; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4329 = 9'h170 == _GEN_13709 & _GEN_15758 | _GEN_2421; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4330 = 9'h170 == _GEN_13709 & _GEN_3588 | _GEN_2933; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4331 = 9'h171 == _GEN_13709 & _GEN_15758 | _GEN_2422; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4332 = 9'h171 == _GEN_13709 & _GEN_3588 | _GEN_2934; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4333 = 9'h172 == _GEN_13709 & _GEN_15758 | _GEN_2423; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4334 = 9'h172 == _GEN_13709 & _GEN_3588 | _GEN_2935; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4335 = 9'h173 == _GEN_13709 & _GEN_15758 | _GEN_2424; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4336 = 9'h173 == _GEN_13709 & _GEN_3588 | _GEN_2936; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4337 = 9'h174 == _GEN_13709 & _GEN_15758 | _GEN_2425; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4338 = 9'h174 == _GEN_13709 & _GEN_3588 | _GEN_2937; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4339 = 9'h175 == _GEN_13709 & _GEN_15758 | _GEN_2426; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4340 = 9'h175 == _GEN_13709 & _GEN_3588 | _GEN_2938; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4341 = 9'h176 == _GEN_13709 & _GEN_15758 | _GEN_2427; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4342 = 9'h176 == _GEN_13709 & _GEN_3588 | _GEN_2939; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4343 = 9'h177 == _GEN_13709 & _GEN_15758 | _GEN_2428; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4344 = 9'h177 == _GEN_13709 & _GEN_3588 | _GEN_2940; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4345 = 9'h178 == _GEN_13709 & _GEN_15758 | _GEN_2429; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4346 = 9'h178 == _GEN_13709 & _GEN_3588 | _GEN_2941; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4347 = 9'h179 == _GEN_13709 & _GEN_15758 | _GEN_2430; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4348 = 9'h179 == _GEN_13709 & _GEN_3588 | _GEN_2942; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4349 = 9'h17a == _GEN_13709 & _GEN_15758 | _GEN_2431; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4350 = 9'h17a == _GEN_13709 & _GEN_3588 | _GEN_2943; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4351 = 9'h17b == _GEN_13709 & _GEN_15758 | _GEN_2432; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4352 = 9'h17b == _GEN_13709 & _GEN_3588 | _GEN_2944; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4353 = 9'h17c == _GEN_13709 & _GEN_15758 | _GEN_2433; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4354 = 9'h17c == _GEN_13709 & _GEN_3588 | _GEN_2945; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4355 = 9'h17d == _GEN_13709 & _GEN_15758 | _GEN_2434; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4356 = 9'h17d == _GEN_13709 & _GEN_3588 | _GEN_2946; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4357 = 9'h17e == _GEN_13709 & _GEN_15758 | _GEN_2435; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4358 = 9'h17e == _GEN_13709 & _GEN_3588 | _GEN_2947; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4359 = 9'h17f == _GEN_13709 & _GEN_15758 | _GEN_2436; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4360 = 9'h17f == _GEN_13709 & _GEN_3588 | _GEN_2948; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4361 = 9'h180 == _GEN_13709 & _GEN_15758 | _GEN_2437; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4362 = 9'h180 == _GEN_13709 & _GEN_3588 | _GEN_2949; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4363 = 9'h181 == _GEN_13709 & _GEN_15758 | _GEN_2438; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4364 = 9'h181 == _GEN_13709 & _GEN_3588 | _GEN_2950; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4365 = 9'h182 == _GEN_13709 & _GEN_15758 | _GEN_2439; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4366 = 9'h182 == _GEN_13709 & _GEN_3588 | _GEN_2951; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4367 = 9'h183 == _GEN_13709 & _GEN_15758 | _GEN_2440; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4368 = 9'h183 == _GEN_13709 & _GEN_3588 | _GEN_2952; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4369 = 9'h184 == _GEN_13709 & _GEN_15758 | _GEN_2441; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4370 = 9'h184 == _GEN_13709 & _GEN_3588 | _GEN_2953; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4371 = 9'h185 == _GEN_13709 & _GEN_15758 | _GEN_2442; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4372 = 9'h185 == _GEN_13709 & _GEN_3588 | _GEN_2954; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4373 = 9'h186 == _GEN_13709 & _GEN_15758 | _GEN_2443; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4374 = 9'h186 == _GEN_13709 & _GEN_3588 | _GEN_2955; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4375 = 9'h187 == _GEN_13709 & _GEN_15758 | _GEN_2444; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4376 = 9'h187 == _GEN_13709 & _GEN_3588 | _GEN_2956; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4377 = 9'h188 == _GEN_13709 & _GEN_15758 | _GEN_2445; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4378 = 9'h188 == _GEN_13709 & _GEN_3588 | _GEN_2957; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4379 = 9'h189 == _GEN_13709 & _GEN_15758 | _GEN_2446; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4380 = 9'h189 == _GEN_13709 & _GEN_3588 | _GEN_2958; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4381 = 9'h18a == _GEN_13709 & _GEN_15758 | _GEN_2447; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4382 = 9'h18a == _GEN_13709 & _GEN_3588 | _GEN_2959; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4383 = 9'h18b == _GEN_13709 & _GEN_15758 | _GEN_2448; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4384 = 9'h18b == _GEN_13709 & _GEN_3588 | _GEN_2960; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4385 = 9'h18c == _GEN_13709 & _GEN_15758 | _GEN_2449; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4386 = 9'h18c == _GEN_13709 & _GEN_3588 | _GEN_2961; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4387 = 9'h18d == _GEN_13709 & _GEN_15758 | _GEN_2450; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4388 = 9'h18d == _GEN_13709 & _GEN_3588 | _GEN_2962; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4389 = 9'h18e == _GEN_13709 & _GEN_15758 | _GEN_2451; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4390 = 9'h18e == _GEN_13709 & _GEN_3588 | _GEN_2963; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4391 = 9'h18f == _GEN_13709 & _GEN_15758 | _GEN_2452; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4392 = 9'h18f == _GEN_13709 & _GEN_3588 | _GEN_2964; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4393 = 9'h190 == _GEN_13709 & _GEN_15758 | _GEN_2453; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4394 = 9'h190 == _GEN_13709 & _GEN_3588 | _GEN_2965; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4395 = 9'h191 == _GEN_13709 & _GEN_15758 | _GEN_2454; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4396 = 9'h191 == _GEN_13709 & _GEN_3588 | _GEN_2966; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4397 = 9'h192 == _GEN_13709 & _GEN_15758 | _GEN_2455; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4398 = 9'h192 == _GEN_13709 & _GEN_3588 | _GEN_2967; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4399 = 9'h193 == _GEN_13709 & _GEN_15758 | _GEN_2456; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4400 = 9'h193 == _GEN_13709 & _GEN_3588 | _GEN_2968; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4401 = 9'h194 == _GEN_13709 & _GEN_15758 | _GEN_2457; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4402 = 9'h194 == _GEN_13709 & _GEN_3588 | _GEN_2969; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4403 = 9'h195 == _GEN_13709 & _GEN_15758 | _GEN_2458; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4404 = 9'h195 == _GEN_13709 & _GEN_3588 | _GEN_2970; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4405 = 9'h196 == _GEN_13709 & _GEN_15758 | _GEN_2459; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4406 = 9'h196 == _GEN_13709 & _GEN_3588 | _GEN_2971; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4407 = 9'h197 == _GEN_13709 & _GEN_15758 | _GEN_2460; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4408 = 9'h197 == _GEN_13709 & _GEN_3588 | _GEN_2972; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4409 = 9'h198 == _GEN_13709 & _GEN_15758 | _GEN_2461; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4410 = 9'h198 == _GEN_13709 & _GEN_3588 | _GEN_2973; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4411 = 9'h199 == _GEN_13709 & _GEN_15758 | _GEN_2462; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4412 = 9'h199 == _GEN_13709 & _GEN_3588 | _GEN_2974; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4413 = 9'h19a == _GEN_13709 & _GEN_15758 | _GEN_2463; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4414 = 9'h19a == _GEN_13709 & _GEN_3588 | _GEN_2975; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4415 = 9'h19b == _GEN_13709 & _GEN_15758 | _GEN_2464; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4416 = 9'h19b == _GEN_13709 & _GEN_3588 | _GEN_2976; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4417 = 9'h19c == _GEN_13709 & _GEN_15758 | _GEN_2465; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4418 = 9'h19c == _GEN_13709 & _GEN_3588 | _GEN_2977; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4419 = 9'h19d == _GEN_13709 & _GEN_15758 | _GEN_2466; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4420 = 9'h19d == _GEN_13709 & _GEN_3588 | _GEN_2978; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4421 = 9'h19e == _GEN_13709 & _GEN_15758 | _GEN_2467; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4422 = 9'h19e == _GEN_13709 & _GEN_3588 | _GEN_2979; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4423 = 9'h19f == _GEN_13709 & _GEN_15758 | _GEN_2468; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4424 = 9'h19f == _GEN_13709 & _GEN_3588 | _GEN_2980; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4425 = 9'h1a0 == _GEN_13709 & _GEN_15758 | _GEN_2469; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4426 = 9'h1a0 == _GEN_13709 & _GEN_3588 | _GEN_2981; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4427 = 9'h1a1 == _GEN_13709 & _GEN_15758 | _GEN_2470; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4428 = 9'h1a1 == _GEN_13709 & _GEN_3588 | _GEN_2982; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4429 = 9'h1a2 == _GEN_13709 & _GEN_15758 | _GEN_2471; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4430 = 9'h1a2 == _GEN_13709 & _GEN_3588 | _GEN_2983; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4431 = 9'h1a3 == _GEN_13709 & _GEN_15758 | _GEN_2472; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4432 = 9'h1a3 == _GEN_13709 & _GEN_3588 | _GEN_2984; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4433 = 9'h1a4 == _GEN_13709 & _GEN_15758 | _GEN_2473; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4434 = 9'h1a4 == _GEN_13709 & _GEN_3588 | _GEN_2985; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4435 = 9'h1a5 == _GEN_13709 & _GEN_15758 | _GEN_2474; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4436 = 9'h1a5 == _GEN_13709 & _GEN_3588 | _GEN_2986; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4437 = 9'h1a6 == _GEN_13709 & _GEN_15758 | _GEN_2475; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4438 = 9'h1a6 == _GEN_13709 & _GEN_3588 | _GEN_2987; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4439 = 9'h1a7 == _GEN_13709 & _GEN_15758 | _GEN_2476; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4440 = 9'h1a7 == _GEN_13709 & _GEN_3588 | _GEN_2988; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4441 = 9'h1a8 == _GEN_13709 & _GEN_15758 | _GEN_2477; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4442 = 9'h1a8 == _GEN_13709 & _GEN_3588 | _GEN_2989; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4443 = 9'h1a9 == _GEN_13709 & _GEN_15758 | _GEN_2478; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4444 = 9'h1a9 == _GEN_13709 & _GEN_3588 | _GEN_2990; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4445 = 9'h1aa == _GEN_13709 & _GEN_15758 | _GEN_2479; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4446 = 9'h1aa == _GEN_13709 & _GEN_3588 | _GEN_2991; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4447 = 9'h1ab == _GEN_13709 & _GEN_15758 | _GEN_2480; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4448 = 9'h1ab == _GEN_13709 & _GEN_3588 | _GEN_2992; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4449 = 9'h1ac == _GEN_13709 & _GEN_15758 | _GEN_2481; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4450 = 9'h1ac == _GEN_13709 & _GEN_3588 | _GEN_2993; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4451 = 9'h1ad == _GEN_13709 & _GEN_15758 | _GEN_2482; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4452 = 9'h1ad == _GEN_13709 & _GEN_3588 | _GEN_2994; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4453 = 9'h1ae == _GEN_13709 & _GEN_15758 | _GEN_2483; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4454 = 9'h1ae == _GEN_13709 & _GEN_3588 | _GEN_2995; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4455 = 9'h1af == _GEN_13709 & _GEN_15758 | _GEN_2484; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4456 = 9'h1af == _GEN_13709 & _GEN_3588 | _GEN_2996; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4457 = 9'h1b0 == _GEN_13709 & _GEN_15758 | _GEN_2485; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4458 = 9'h1b0 == _GEN_13709 & _GEN_3588 | _GEN_2997; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4459 = 9'h1b1 == _GEN_13709 & _GEN_15758 | _GEN_2486; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4460 = 9'h1b1 == _GEN_13709 & _GEN_3588 | _GEN_2998; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4461 = 9'h1b2 == _GEN_13709 & _GEN_15758 | _GEN_2487; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4462 = 9'h1b2 == _GEN_13709 & _GEN_3588 | _GEN_2999; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4463 = 9'h1b3 == _GEN_13709 & _GEN_15758 | _GEN_2488; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4464 = 9'h1b3 == _GEN_13709 & _GEN_3588 | _GEN_3000; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4465 = 9'h1b4 == _GEN_13709 & _GEN_15758 | _GEN_2489; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4466 = 9'h1b4 == _GEN_13709 & _GEN_3588 | _GEN_3001; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4467 = 9'h1b5 == _GEN_13709 & _GEN_15758 | _GEN_2490; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4468 = 9'h1b5 == _GEN_13709 & _GEN_3588 | _GEN_3002; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4469 = 9'h1b6 == _GEN_13709 & _GEN_15758 | _GEN_2491; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4470 = 9'h1b6 == _GEN_13709 & _GEN_3588 | _GEN_3003; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4471 = 9'h1b7 == _GEN_13709 & _GEN_15758 | _GEN_2492; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4472 = 9'h1b7 == _GEN_13709 & _GEN_3588 | _GEN_3004; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4473 = 9'h1b8 == _GEN_13709 & _GEN_15758 | _GEN_2493; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4474 = 9'h1b8 == _GEN_13709 & _GEN_3588 | _GEN_3005; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4475 = 9'h1b9 == _GEN_13709 & _GEN_15758 | _GEN_2494; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4476 = 9'h1b9 == _GEN_13709 & _GEN_3588 | _GEN_3006; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4477 = 9'h1ba == _GEN_13709 & _GEN_15758 | _GEN_2495; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4478 = 9'h1ba == _GEN_13709 & _GEN_3588 | _GEN_3007; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4479 = 9'h1bb == _GEN_13709 & _GEN_15758 | _GEN_2496; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4480 = 9'h1bb == _GEN_13709 & _GEN_3588 | _GEN_3008; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4481 = 9'h1bc == _GEN_13709 & _GEN_15758 | _GEN_2497; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4482 = 9'h1bc == _GEN_13709 & _GEN_3588 | _GEN_3009; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4483 = 9'h1bd == _GEN_13709 & _GEN_15758 | _GEN_2498; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4484 = 9'h1bd == _GEN_13709 & _GEN_3588 | _GEN_3010; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4485 = 9'h1be == _GEN_13709 & _GEN_15758 | _GEN_2499; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4486 = 9'h1be == _GEN_13709 & _GEN_3588 | _GEN_3011; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4487 = 9'h1bf == _GEN_13709 & _GEN_15758 | _GEN_2500; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4488 = 9'h1bf == _GEN_13709 & _GEN_3588 | _GEN_3012; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4489 = 9'h1c0 == _GEN_13709 & _GEN_15758 | _GEN_2501; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4490 = 9'h1c0 == _GEN_13709 & _GEN_3588 | _GEN_3013; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4491 = 9'h1c1 == _GEN_13709 & _GEN_15758 | _GEN_2502; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4492 = 9'h1c1 == _GEN_13709 & _GEN_3588 | _GEN_3014; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4493 = 9'h1c2 == _GEN_13709 & _GEN_15758 | _GEN_2503; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4494 = 9'h1c2 == _GEN_13709 & _GEN_3588 | _GEN_3015; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4495 = 9'h1c3 == _GEN_13709 & _GEN_15758 | _GEN_2504; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4496 = 9'h1c3 == _GEN_13709 & _GEN_3588 | _GEN_3016; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4497 = 9'h1c4 == _GEN_13709 & _GEN_15758 | _GEN_2505; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4498 = 9'h1c4 == _GEN_13709 & _GEN_3588 | _GEN_3017; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4499 = 9'h1c5 == _GEN_13709 & _GEN_15758 | _GEN_2506; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4500 = 9'h1c5 == _GEN_13709 & _GEN_3588 | _GEN_3018; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4501 = 9'h1c6 == _GEN_13709 & _GEN_15758 | _GEN_2507; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4502 = 9'h1c6 == _GEN_13709 & _GEN_3588 | _GEN_3019; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4503 = 9'h1c7 == _GEN_13709 & _GEN_15758 | _GEN_2508; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4504 = 9'h1c7 == _GEN_13709 & _GEN_3588 | _GEN_3020; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4505 = 9'h1c8 == _GEN_13709 & _GEN_15758 | _GEN_2509; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4506 = 9'h1c8 == _GEN_13709 & _GEN_3588 | _GEN_3021; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4507 = 9'h1c9 == _GEN_13709 & _GEN_15758 | _GEN_2510; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4508 = 9'h1c9 == _GEN_13709 & _GEN_3588 | _GEN_3022; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4509 = 9'h1ca == _GEN_13709 & _GEN_15758 | _GEN_2511; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4510 = 9'h1ca == _GEN_13709 & _GEN_3588 | _GEN_3023; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4511 = 9'h1cb == _GEN_13709 & _GEN_15758 | _GEN_2512; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4512 = 9'h1cb == _GEN_13709 & _GEN_3588 | _GEN_3024; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4513 = 9'h1cc == _GEN_13709 & _GEN_15758 | _GEN_2513; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4514 = 9'h1cc == _GEN_13709 & _GEN_3588 | _GEN_3025; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4515 = 9'h1cd == _GEN_13709 & _GEN_15758 | _GEN_2514; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4516 = 9'h1cd == _GEN_13709 & _GEN_3588 | _GEN_3026; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4517 = 9'h1ce == _GEN_13709 & _GEN_15758 | _GEN_2515; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4518 = 9'h1ce == _GEN_13709 & _GEN_3588 | _GEN_3027; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4519 = 9'h1cf == _GEN_13709 & _GEN_15758 | _GEN_2516; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4520 = 9'h1cf == _GEN_13709 & _GEN_3588 | _GEN_3028; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4521 = 9'h1d0 == _GEN_13709 & _GEN_15758 | _GEN_2517; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4522 = 9'h1d0 == _GEN_13709 & _GEN_3588 | _GEN_3029; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4523 = 9'h1d1 == _GEN_13709 & _GEN_15758 | _GEN_2518; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4524 = 9'h1d1 == _GEN_13709 & _GEN_3588 | _GEN_3030; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4525 = 9'h1d2 == _GEN_13709 & _GEN_15758 | _GEN_2519; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4526 = 9'h1d2 == _GEN_13709 & _GEN_3588 | _GEN_3031; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4527 = 9'h1d3 == _GEN_13709 & _GEN_15758 | _GEN_2520; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4528 = 9'h1d3 == _GEN_13709 & _GEN_3588 | _GEN_3032; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4529 = 9'h1d4 == _GEN_13709 & _GEN_15758 | _GEN_2521; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4530 = 9'h1d4 == _GEN_13709 & _GEN_3588 | _GEN_3033; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4531 = 9'h1d5 == _GEN_13709 & _GEN_15758 | _GEN_2522; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4532 = 9'h1d5 == _GEN_13709 & _GEN_3588 | _GEN_3034; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4533 = 9'h1d6 == _GEN_13709 & _GEN_15758 | _GEN_2523; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4534 = 9'h1d6 == _GEN_13709 & _GEN_3588 | _GEN_3035; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4535 = 9'h1d7 == _GEN_13709 & _GEN_15758 | _GEN_2524; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4536 = 9'h1d7 == _GEN_13709 & _GEN_3588 | _GEN_3036; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4537 = 9'h1d8 == _GEN_13709 & _GEN_15758 | _GEN_2525; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4538 = 9'h1d8 == _GEN_13709 & _GEN_3588 | _GEN_3037; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4539 = 9'h1d9 == _GEN_13709 & _GEN_15758 | _GEN_2526; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4540 = 9'h1d9 == _GEN_13709 & _GEN_3588 | _GEN_3038; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4541 = 9'h1da == _GEN_13709 & _GEN_15758 | _GEN_2527; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4542 = 9'h1da == _GEN_13709 & _GEN_3588 | _GEN_3039; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4543 = 9'h1db == _GEN_13709 & _GEN_15758 | _GEN_2528; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4544 = 9'h1db == _GEN_13709 & _GEN_3588 | _GEN_3040; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4545 = 9'h1dc == _GEN_13709 & _GEN_15758 | _GEN_2529; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4546 = 9'h1dc == _GEN_13709 & _GEN_3588 | _GEN_3041; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4547 = 9'h1dd == _GEN_13709 & _GEN_15758 | _GEN_2530; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4548 = 9'h1dd == _GEN_13709 & _GEN_3588 | _GEN_3042; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4549 = 9'h1de == _GEN_13709 & _GEN_15758 | _GEN_2531; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4550 = 9'h1de == _GEN_13709 & _GEN_3588 | _GEN_3043; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4551 = 9'h1df == _GEN_13709 & _GEN_15758 | _GEN_2532; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4552 = 9'h1df == _GEN_13709 & _GEN_3588 | _GEN_3044; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4553 = 9'h1e0 == _GEN_13709 & _GEN_15758 | _GEN_2533; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4554 = 9'h1e0 == _GEN_13709 & _GEN_3588 | _GEN_3045; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4555 = 9'h1e1 == _GEN_13709 & _GEN_15758 | _GEN_2534; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4556 = 9'h1e1 == _GEN_13709 & _GEN_3588 | _GEN_3046; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4557 = 9'h1e2 == _GEN_13709 & _GEN_15758 | _GEN_2535; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4558 = 9'h1e2 == _GEN_13709 & _GEN_3588 | _GEN_3047; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4559 = 9'h1e3 == _GEN_13709 & _GEN_15758 | _GEN_2536; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4560 = 9'h1e3 == _GEN_13709 & _GEN_3588 | _GEN_3048; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4561 = 9'h1e4 == _GEN_13709 & _GEN_15758 | _GEN_2537; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4562 = 9'h1e4 == _GEN_13709 & _GEN_3588 | _GEN_3049; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4563 = 9'h1e5 == _GEN_13709 & _GEN_15758 | _GEN_2538; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4564 = 9'h1e5 == _GEN_13709 & _GEN_3588 | _GEN_3050; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4565 = 9'h1e6 == _GEN_13709 & _GEN_15758 | _GEN_2539; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4566 = 9'h1e6 == _GEN_13709 & _GEN_3588 | _GEN_3051; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4567 = 9'h1e7 == _GEN_13709 & _GEN_15758 | _GEN_2540; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4568 = 9'h1e7 == _GEN_13709 & _GEN_3588 | _GEN_3052; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4569 = 9'h1e8 == _GEN_13709 & _GEN_15758 | _GEN_2541; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4570 = 9'h1e8 == _GEN_13709 & _GEN_3588 | _GEN_3053; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4571 = 9'h1e9 == _GEN_13709 & _GEN_15758 | _GEN_2542; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4572 = 9'h1e9 == _GEN_13709 & _GEN_3588 | _GEN_3054; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4573 = 9'h1ea == _GEN_13709 & _GEN_15758 | _GEN_2543; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4574 = 9'h1ea == _GEN_13709 & _GEN_3588 | _GEN_3055; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4575 = 9'h1eb == _GEN_13709 & _GEN_15758 | _GEN_2544; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4576 = 9'h1eb == _GEN_13709 & _GEN_3588 | _GEN_3056; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4577 = 9'h1ec == _GEN_13709 & _GEN_15758 | _GEN_2545; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4578 = 9'h1ec == _GEN_13709 & _GEN_3588 | _GEN_3057; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4579 = 9'h1ed == _GEN_13709 & _GEN_15758 | _GEN_2546; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4580 = 9'h1ed == _GEN_13709 & _GEN_3588 | _GEN_3058; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4581 = 9'h1ee == _GEN_13709 & _GEN_15758 | _GEN_2547; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4582 = 9'h1ee == _GEN_13709 & _GEN_3588 | _GEN_3059; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4583 = 9'h1ef == _GEN_13709 & _GEN_15758 | _GEN_2548; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4584 = 9'h1ef == _GEN_13709 & _GEN_3588 | _GEN_3060; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4585 = 9'h1f0 == _GEN_13709 & _GEN_15758 | _GEN_2549; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4586 = 9'h1f0 == _GEN_13709 & _GEN_3588 | _GEN_3061; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4587 = 9'h1f1 == _GEN_13709 & _GEN_15758 | _GEN_2550; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4588 = 9'h1f1 == _GEN_13709 & _GEN_3588 | _GEN_3062; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4589 = 9'h1f2 == _GEN_13709 & _GEN_15758 | _GEN_2551; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4590 = 9'h1f2 == _GEN_13709 & _GEN_3588 | _GEN_3063; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4591 = 9'h1f3 == _GEN_13709 & _GEN_15758 | _GEN_2552; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4592 = 9'h1f3 == _GEN_13709 & _GEN_3588 | _GEN_3064; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4593 = 9'h1f4 == _GEN_13709 & _GEN_15758 | _GEN_2553; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4594 = 9'h1f4 == _GEN_13709 & _GEN_3588 | _GEN_3065; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4595 = 9'h1f5 == _GEN_13709 & _GEN_15758 | _GEN_2554; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4596 = 9'h1f5 == _GEN_13709 & _GEN_3588 | _GEN_3066; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4597 = 9'h1f6 == _GEN_13709 & _GEN_15758 | _GEN_2555; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4598 = 9'h1f6 == _GEN_13709 & _GEN_3588 | _GEN_3067; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4599 = 9'h1f7 == _GEN_13709 & _GEN_15758 | _GEN_2556; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4600 = 9'h1f7 == _GEN_13709 & _GEN_3588 | _GEN_3068; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4601 = 9'h1f8 == _GEN_13709 & _GEN_15758 | _GEN_2557; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4602 = 9'h1f8 == _GEN_13709 & _GEN_3588 | _GEN_3069; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4603 = 9'h1f9 == _GEN_13709 & _GEN_15758 | _GEN_2558; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4604 = 9'h1f9 == _GEN_13709 & _GEN_3588 | _GEN_3070; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4605 = 9'h1fa == _GEN_13709 & _GEN_15758 | _GEN_2559; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4606 = 9'h1fa == _GEN_13709 & _GEN_3588 | _GEN_3071; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4607 = 9'h1fb == _GEN_13709 & _GEN_15758 | _GEN_2560; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4608 = 9'h1fb == _GEN_13709 & _GEN_3588 | _GEN_3072; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4609 = 9'h1fc == _GEN_13709 & _GEN_15758 | _GEN_2561; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4610 = 9'h1fc == _GEN_13709 & _GEN_3588 | _GEN_3073; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4611 = 9'h1fd == _GEN_13709 & _GEN_15758 | _GEN_2562; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4612 = 9'h1fd == _GEN_13709 & _GEN_3588 | _GEN_3074; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4613 = 9'h1fe == _GEN_13709 & _GEN_15758 | _GEN_2563; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4614 = 9'h1fe == _GEN_13709 & _GEN_3588 | _GEN_3075; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4615 = 9'h1ff == _GEN_13709 & _GEN_15758 | _GEN_2564; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4616 = 9'h1ff == _GEN_13709 & _GEN_3588 | _GEN_3076; // @[ICache.scala 186:{60,60}]
  wire  _GEN_4617 = 6'h0 == va_line_addr ? ~tag_compare_valid_1 : meta_0_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4618 = 6'h1 == va_line_addr ? ~tag_compare_valid_1 : meta_1_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4619 = 6'h2 == va_line_addr ? ~tag_compare_valid_1 : meta_2_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4620 = 6'h3 == va_line_addr ? ~tag_compare_valid_1 : meta_3_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4621 = 6'h4 == va_line_addr ? ~tag_compare_valid_1 : meta_4_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4622 = 6'h5 == va_line_addr ? ~tag_compare_valid_1 : meta_5_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4623 = 6'h6 == va_line_addr ? ~tag_compare_valid_1 : meta_6_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4624 = 6'h7 == va_line_addr ? ~tag_compare_valid_1 : meta_7_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4625 = 6'h8 == va_line_addr ? ~tag_compare_valid_1 : meta_8_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4626 = 6'h9 == va_line_addr ? ~tag_compare_valid_1 : meta_9_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4627 = 6'ha == va_line_addr ? ~tag_compare_valid_1 : meta_10_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4628 = 6'hb == va_line_addr ? ~tag_compare_valid_1 : meta_11_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4629 = 6'hc == va_line_addr ? ~tag_compare_valid_1 : meta_12_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4630 = 6'hd == va_line_addr ? ~tag_compare_valid_1 : meta_13_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4631 = 6'he == va_line_addr ? ~tag_compare_valid_1 : meta_14_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4632 = 6'hf == va_line_addr ? ~tag_compare_valid_1 : meta_15_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4633 = 6'h10 == va_line_addr ? ~tag_compare_valid_1 : meta_16_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4634 = 6'h11 == va_line_addr ? ~tag_compare_valid_1 : meta_17_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4635 = 6'h12 == va_line_addr ? ~tag_compare_valid_1 : meta_18_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4636 = 6'h13 == va_line_addr ? ~tag_compare_valid_1 : meta_19_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4637 = 6'h14 == va_line_addr ? ~tag_compare_valid_1 : meta_20_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4638 = 6'h15 == va_line_addr ? ~tag_compare_valid_1 : meta_21_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4639 = 6'h16 == va_line_addr ? ~tag_compare_valid_1 : meta_22_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4640 = 6'h17 == va_line_addr ? ~tag_compare_valid_1 : meta_23_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4641 = 6'h18 == va_line_addr ? ~tag_compare_valid_1 : meta_24_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4642 = 6'h19 == va_line_addr ? ~tag_compare_valid_1 : meta_25_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4643 = 6'h1a == va_line_addr ? ~tag_compare_valid_1 : meta_26_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4644 = 6'h1b == va_line_addr ? ~tag_compare_valid_1 : meta_27_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4645 = 6'h1c == va_line_addr ? ~tag_compare_valid_1 : meta_28_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4646 = 6'h1d == va_line_addr ? ~tag_compare_valid_1 : meta_29_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4647 = 6'h1e == va_line_addr ? ~tag_compare_valid_1 : meta_30_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4648 = 6'h1f == va_line_addr ? ~tag_compare_valid_1 : meta_31_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4649 = 6'h20 == va_line_addr ? ~tag_compare_valid_1 : meta_32_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4650 = 6'h21 == va_line_addr ? ~tag_compare_valid_1 : meta_33_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4651 = 6'h22 == va_line_addr ? ~tag_compare_valid_1 : meta_34_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4652 = 6'h23 == va_line_addr ? ~tag_compare_valid_1 : meta_35_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4653 = 6'h24 == va_line_addr ? ~tag_compare_valid_1 : meta_36_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4654 = 6'h25 == va_line_addr ? ~tag_compare_valid_1 : meta_37_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4655 = 6'h26 == va_line_addr ? ~tag_compare_valid_1 : meta_38_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4656 = 6'h27 == va_line_addr ? ~tag_compare_valid_1 : meta_39_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4657 = 6'h28 == va_line_addr ? ~tag_compare_valid_1 : meta_40_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4658 = 6'h29 == va_line_addr ? ~tag_compare_valid_1 : meta_41_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4659 = 6'h2a == va_line_addr ? ~tag_compare_valid_1 : meta_42_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4660 = 6'h2b == va_line_addr ? ~tag_compare_valid_1 : meta_43_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4661 = 6'h2c == va_line_addr ? ~tag_compare_valid_1 : meta_44_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4662 = 6'h2d == va_line_addr ? ~tag_compare_valid_1 : meta_45_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4663 = 6'h2e == va_line_addr ? ~tag_compare_valid_1 : meta_46_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4664 = 6'h2f == va_line_addr ? ~tag_compare_valid_1 : meta_47_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4665 = 6'h30 == va_line_addr ? ~tag_compare_valid_1 : meta_48_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4666 = 6'h31 == va_line_addr ? ~tag_compare_valid_1 : meta_49_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4667 = 6'h32 == va_line_addr ? ~tag_compare_valid_1 : meta_50_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4668 = 6'h33 == va_line_addr ? ~tag_compare_valid_1 : meta_51_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4669 = 6'h34 == va_line_addr ? ~tag_compare_valid_1 : meta_52_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4670 = 6'h35 == va_line_addr ? ~tag_compare_valid_1 : meta_53_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4671 = 6'h36 == va_line_addr ? ~tag_compare_valid_1 : meta_54_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4672 = 6'h37 == va_line_addr ? ~tag_compare_valid_1 : meta_55_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4673 = 6'h38 == va_line_addr ? ~tag_compare_valid_1 : meta_56_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4674 = 6'h39 == va_line_addr ? ~tag_compare_valid_1 : meta_57_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4675 = 6'h3a == va_line_addr ? ~tag_compare_valid_1 : meta_58_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4676 = 6'h3b == va_line_addr ? ~tag_compare_valid_1 : meta_59_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4677 = 6'h3c == va_line_addr ? ~tag_compare_valid_1 : meta_60_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4678 = 6'h3d == va_line_addr ? ~tag_compare_valid_1 : meta_61_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4679 = 6'h3e == va_line_addr ? ~tag_compare_valid_1 : meta_62_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4680 = 6'h3f == va_line_addr ? ~tag_compare_valid_1 : meta_63_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4681 = 7'h40 == _GEN_13517 ? ~tag_compare_valid_1 : meta_64_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4682 = 7'h41 == _GEN_13517 ? ~tag_compare_valid_1 : meta_65_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4683 = 7'h42 == _GEN_13517 ? ~tag_compare_valid_1 : meta_66_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4684 = 7'h43 == _GEN_13517 ? ~tag_compare_valid_1 : meta_67_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4685 = 7'h44 == _GEN_13517 ? ~tag_compare_valid_1 : meta_68_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4686 = 7'h45 == _GEN_13517 ? ~tag_compare_valid_1 : meta_69_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4687 = 7'h46 == _GEN_13517 ? ~tag_compare_valid_1 : meta_70_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4688 = 7'h47 == _GEN_13517 ? ~tag_compare_valid_1 : meta_71_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4689 = 7'h48 == _GEN_13517 ? ~tag_compare_valid_1 : meta_72_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4690 = 7'h49 == _GEN_13517 ? ~tag_compare_valid_1 : meta_73_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4691 = 7'h4a == _GEN_13517 ? ~tag_compare_valid_1 : meta_74_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4692 = 7'h4b == _GEN_13517 ? ~tag_compare_valid_1 : meta_75_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4693 = 7'h4c == _GEN_13517 ? ~tag_compare_valid_1 : meta_76_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4694 = 7'h4d == _GEN_13517 ? ~tag_compare_valid_1 : meta_77_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4695 = 7'h4e == _GEN_13517 ? ~tag_compare_valid_1 : meta_78_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4696 = 7'h4f == _GEN_13517 ? ~tag_compare_valid_1 : meta_79_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4697 = 7'h50 == _GEN_13517 ? ~tag_compare_valid_1 : meta_80_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4698 = 7'h51 == _GEN_13517 ? ~tag_compare_valid_1 : meta_81_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4699 = 7'h52 == _GEN_13517 ? ~tag_compare_valid_1 : meta_82_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4700 = 7'h53 == _GEN_13517 ? ~tag_compare_valid_1 : meta_83_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4701 = 7'h54 == _GEN_13517 ? ~tag_compare_valid_1 : meta_84_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4702 = 7'h55 == _GEN_13517 ? ~tag_compare_valid_1 : meta_85_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4703 = 7'h56 == _GEN_13517 ? ~tag_compare_valid_1 : meta_86_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4704 = 7'h57 == _GEN_13517 ? ~tag_compare_valid_1 : meta_87_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4705 = 7'h58 == _GEN_13517 ? ~tag_compare_valid_1 : meta_88_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4706 = 7'h59 == _GEN_13517 ? ~tag_compare_valid_1 : meta_89_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4707 = 7'h5a == _GEN_13517 ? ~tag_compare_valid_1 : meta_90_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4708 = 7'h5b == _GEN_13517 ? ~tag_compare_valid_1 : meta_91_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4709 = 7'h5c == _GEN_13517 ? ~tag_compare_valid_1 : meta_92_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4710 = 7'h5d == _GEN_13517 ? ~tag_compare_valid_1 : meta_93_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4711 = 7'h5e == _GEN_13517 ? ~tag_compare_valid_1 : meta_94_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4712 = 7'h5f == _GEN_13517 ? ~tag_compare_valid_1 : meta_95_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4713 = 7'h60 == _GEN_13517 ? ~tag_compare_valid_1 : meta_96_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4714 = 7'h61 == _GEN_13517 ? ~tag_compare_valid_1 : meta_97_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4715 = 7'h62 == _GEN_13517 ? ~tag_compare_valid_1 : meta_98_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4716 = 7'h63 == _GEN_13517 ? ~tag_compare_valid_1 : meta_99_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4717 = 7'h64 == _GEN_13517 ? ~tag_compare_valid_1 : meta_100_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4718 = 7'h65 == _GEN_13517 ? ~tag_compare_valid_1 : meta_101_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4719 = 7'h66 == _GEN_13517 ? ~tag_compare_valid_1 : meta_102_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4720 = 7'h67 == _GEN_13517 ? ~tag_compare_valid_1 : meta_103_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4721 = 7'h68 == _GEN_13517 ? ~tag_compare_valid_1 : meta_104_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4722 = 7'h69 == _GEN_13517 ? ~tag_compare_valid_1 : meta_105_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4723 = 7'h6a == _GEN_13517 ? ~tag_compare_valid_1 : meta_106_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4724 = 7'h6b == _GEN_13517 ? ~tag_compare_valid_1 : meta_107_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4725 = 7'h6c == _GEN_13517 ? ~tag_compare_valid_1 : meta_108_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4726 = 7'h6d == _GEN_13517 ? ~tag_compare_valid_1 : meta_109_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4727 = 7'h6e == _GEN_13517 ? ~tag_compare_valid_1 : meta_110_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4728 = 7'h6f == _GEN_13517 ? ~tag_compare_valid_1 : meta_111_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4729 = 7'h70 == _GEN_13517 ? ~tag_compare_valid_1 : meta_112_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4730 = 7'h71 == _GEN_13517 ? ~tag_compare_valid_1 : meta_113_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4731 = 7'h72 == _GEN_13517 ? ~tag_compare_valid_1 : meta_114_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4732 = 7'h73 == _GEN_13517 ? ~tag_compare_valid_1 : meta_115_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4733 = 7'h74 == _GEN_13517 ? ~tag_compare_valid_1 : meta_116_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4734 = 7'h75 == _GEN_13517 ? ~tag_compare_valid_1 : meta_117_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4735 = 7'h76 == _GEN_13517 ? ~tag_compare_valid_1 : meta_118_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4736 = 7'h77 == _GEN_13517 ? ~tag_compare_valid_1 : meta_119_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4737 = 7'h78 == _GEN_13517 ? ~tag_compare_valid_1 : meta_120_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4738 = 7'h79 == _GEN_13517 ? ~tag_compare_valid_1 : meta_121_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4739 = 7'h7a == _GEN_13517 ? ~tag_compare_valid_1 : meta_122_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4740 = 7'h7b == _GEN_13517 ? ~tag_compare_valid_1 : meta_123_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4741 = 7'h7c == _GEN_13517 ? ~tag_compare_valid_1 : meta_124_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4742 = 7'h7d == _GEN_13517 ? ~tag_compare_valid_1 : meta_125_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4743 = 7'h7e == _GEN_13517 ? ~tag_compare_valid_1 : meta_126_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4744 = 7'h7f == _GEN_13517 ? ~tag_compare_valid_1 : meta_127_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4745 = 8'h80 == _GEN_13581 ? ~tag_compare_valid_1 : meta_128_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4746 = 8'h81 == _GEN_13581 ? ~tag_compare_valid_1 : meta_129_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4747 = 8'h82 == _GEN_13581 ? ~tag_compare_valid_1 : meta_130_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4748 = 8'h83 == _GEN_13581 ? ~tag_compare_valid_1 : meta_131_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4749 = 8'h84 == _GEN_13581 ? ~tag_compare_valid_1 : meta_132_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4750 = 8'h85 == _GEN_13581 ? ~tag_compare_valid_1 : meta_133_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4751 = 8'h86 == _GEN_13581 ? ~tag_compare_valid_1 : meta_134_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4752 = 8'h87 == _GEN_13581 ? ~tag_compare_valid_1 : meta_135_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4753 = 8'h88 == _GEN_13581 ? ~tag_compare_valid_1 : meta_136_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4754 = 8'h89 == _GEN_13581 ? ~tag_compare_valid_1 : meta_137_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4755 = 8'h8a == _GEN_13581 ? ~tag_compare_valid_1 : meta_138_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4756 = 8'h8b == _GEN_13581 ? ~tag_compare_valid_1 : meta_139_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4757 = 8'h8c == _GEN_13581 ? ~tag_compare_valid_1 : meta_140_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4758 = 8'h8d == _GEN_13581 ? ~tag_compare_valid_1 : meta_141_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4759 = 8'h8e == _GEN_13581 ? ~tag_compare_valid_1 : meta_142_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4760 = 8'h8f == _GEN_13581 ? ~tag_compare_valid_1 : meta_143_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4761 = 8'h90 == _GEN_13581 ? ~tag_compare_valid_1 : meta_144_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4762 = 8'h91 == _GEN_13581 ? ~tag_compare_valid_1 : meta_145_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4763 = 8'h92 == _GEN_13581 ? ~tag_compare_valid_1 : meta_146_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4764 = 8'h93 == _GEN_13581 ? ~tag_compare_valid_1 : meta_147_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4765 = 8'h94 == _GEN_13581 ? ~tag_compare_valid_1 : meta_148_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4766 = 8'h95 == _GEN_13581 ? ~tag_compare_valid_1 : meta_149_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4767 = 8'h96 == _GEN_13581 ? ~tag_compare_valid_1 : meta_150_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4768 = 8'h97 == _GEN_13581 ? ~tag_compare_valid_1 : meta_151_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4769 = 8'h98 == _GEN_13581 ? ~tag_compare_valid_1 : meta_152_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4770 = 8'h99 == _GEN_13581 ? ~tag_compare_valid_1 : meta_153_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4771 = 8'h9a == _GEN_13581 ? ~tag_compare_valid_1 : meta_154_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4772 = 8'h9b == _GEN_13581 ? ~tag_compare_valid_1 : meta_155_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4773 = 8'h9c == _GEN_13581 ? ~tag_compare_valid_1 : meta_156_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4774 = 8'h9d == _GEN_13581 ? ~tag_compare_valid_1 : meta_157_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4775 = 8'h9e == _GEN_13581 ? ~tag_compare_valid_1 : meta_158_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4776 = 8'h9f == _GEN_13581 ? ~tag_compare_valid_1 : meta_159_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4777 = 8'ha0 == _GEN_13581 ? ~tag_compare_valid_1 : meta_160_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4778 = 8'ha1 == _GEN_13581 ? ~tag_compare_valid_1 : meta_161_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4779 = 8'ha2 == _GEN_13581 ? ~tag_compare_valid_1 : meta_162_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4780 = 8'ha3 == _GEN_13581 ? ~tag_compare_valid_1 : meta_163_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4781 = 8'ha4 == _GEN_13581 ? ~tag_compare_valid_1 : meta_164_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4782 = 8'ha5 == _GEN_13581 ? ~tag_compare_valid_1 : meta_165_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4783 = 8'ha6 == _GEN_13581 ? ~tag_compare_valid_1 : meta_166_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4784 = 8'ha7 == _GEN_13581 ? ~tag_compare_valid_1 : meta_167_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4785 = 8'ha8 == _GEN_13581 ? ~tag_compare_valid_1 : meta_168_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4786 = 8'ha9 == _GEN_13581 ? ~tag_compare_valid_1 : meta_169_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4787 = 8'haa == _GEN_13581 ? ~tag_compare_valid_1 : meta_170_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4788 = 8'hab == _GEN_13581 ? ~tag_compare_valid_1 : meta_171_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4789 = 8'hac == _GEN_13581 ? ~tag_compare_valid_1 : meta_172_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4790 = 8'had == _GEN_13581 ? ~tag_compare_valid_1 : meta_173_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4791 = 8'hae == _GEN_13581 ? ~tag_compare_valid_1 : meta_174_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4792 = 8'haf == _GEN_13581 ? ~tag_compare_valid_1 : meta_175_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4793 = 8'hb0 == _GEN_13581 ? ~tag_compare_valid_1 : meta_176_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4794 = 8'hb1 == _GEN_13581 ? ~tag_compare_valid_1 : meta_177_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4795 = 8'hb2 == _GEN_13581 ? ~tag_compare_valid_1 : meta_178_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4796 = 8'hb3 == _GEN_13581 ? ~tag_compare_valid_1 : meta_179_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4797 = 8'hb4 == _GEN_13581 ? ~tag_compare_valid_1 : meta_180_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4798 = 8'hb5 == _GEN_13581 ? ~tag_compare_valid_1 : meta_181_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4799 = 8'hb6 == _GEN_13581 ? ~tag_compare_valid_1 : meta_182_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4800 = 8'hb7 == _GEN_13581 ? ~tag_compare_valid_1 : meta_183_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4801 = 8'hb8 == _GEN_13581 ? ~tag_compare_valid_1 : meta_184_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4802 = 8'hb9 == _GEN_13581 ? ~tag_compare_valid_1 : meta_185_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4803 = 8'hba == _GEN_13581 ? ~tag_compare_valid_1 : meta_186_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4804 = 8'hbb == _GEN_13581 ? ~tag_compare_valid_1 : meta_187_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4805 = 8'hbc == _GEN_13581 ? ~tag_compare_valid_1 : meta_188_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4806 = 8'hbd == _GEN_13581 ? ~tag_compare_valid_1 : meta_189_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4807 = 8'hbe == _GEN_13581 ? ~tag_compare_valid_1 : meta_190_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4808 = 8'hbf == _GEN_13581 ? ~tag_compare_valid_1 : meta_191_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4809 = 8'hc0 == _GEN_13581 ? ~tag_compare_valid_1 : meta_192_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4810 = 8'hc1 == _GEN_13581 ? ~tag_compare_valid_1 : meta_193_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4811 = 8'hc2 == _GEN_13581 ? ~tag_compare_valid_1 : meta_194_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4812 = 8'hc3 == _GEN_13581 ? ~tag_compare_valid_1 : meta_195_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4813 = 8'hc4 == _GEN_13581 ? ~tag_compare_valid_1 : meta_196_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4814 = 8'hc5 == _GEN_13581 ? ~tag_compare_valid_1 : meta_197_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4815 = 8'hc6 == _GEN_13581 ? ~tag_compare_valid_1 : meta_198_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4816 = 8'hc7 == _GEN_13581 ? ~tag_compare_valid_1 : meta_199_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4817 = 8'hc8 == _GEN_13581 ? ~tag_compare_valid_1 : meta_200_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4818 = 8'hc9 == _GEN_13581 ? ~tag_compare_valid_1 : meta_201_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4819 = 8'hca == _GEN_13581 ? ~tag_compare_valid_1 : meta_202_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4820 = 8'hcb == _GEN_13581 ? ~tag_compare_valid_1 : meta_203_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4821 = 8'hcc == _GEN_13581 ? ~tag_compare_valid_1 : meta_204_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4822 = 8'hcd == _GEN_13581 ? ~tag_compare_valid_1 : meta_205_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4823 = 8'hce == _GEN_13581 ? ~tag_compare_valid_1 : meta_206_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4824 = 8'hcf == _GEN_13581 ? ~tag_compare_valid_1 : meta_207_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4825 = 8'hd0 == _GEN_13581 ? ~tag_compare_valid_1 : meta_208_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4826 = 8'hd1 == _GEN_13581 ? ~tag_compare_valid_1 : meta_209_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4827 = 8'hd2 == _GEN_13581 ? ~tag_compare_valid_1 : meta_210_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4828 = 8'hd3 == _GEN_13581 ? ~tag_compare_valid_1 : meta_211_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4829 = 8'hd4 == _GEN_13581 ? ~tag_compare_valid_1 : meta_212_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4830 = 8'hd5 == _GEN_13581 ? ~tag_compare_valid_1 : meta_213_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4831 = 8'hd6 == _GEN_13581 ? ~tag_compare_valid_1 : meta_214_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4832 = 8'hd7 == _GEN_13581 ? ~tag_compare_valid_1 : meta_215_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4833 = 8'hd8 == _GEN_13581 ? ~tag_compare_valid_1 : meta_216_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4834 = 8'hd9 == _GEN_13581 ? ~tag_compare_valid_1 : meta_217_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4835 = 8'hda == _GEN_13581 ? ~tag_compare_valid_1 : meta_218_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4836 = 8'hdb == _GEN_13581 ? ~tag_compare_valid_1 : meta_219_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4837 = 8'hdc == _GEN_13581 ? ~tag_compare_valid_1 : meta_220_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4838 = 8'hdd == _GEN_13581 ? ~tag_compare_valid_1 : meta_221_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4839 = 8'hde == _GEN_13581 ? ~tag_compare_valid_1 : meta_222_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4840 = 8'hdf == _GEN_13581 ? ~tag_compare_valid_1 : meta_223_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4841 = 8'he0 == _GEN_13581 ? ~tag_compare_valid_1 : meta_224_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4842 = 8'he1 == _GEN_13581 ? ~tag_compare_valid_1 : meta_225_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4843 = 8'he2 == _GEN_13581 ? ~tag_compare_valid_1 : meta_226_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4844 = 8'he3 == _GEN_13581 ? ~tag_compare_valid_1 : meta_227_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4845 = 8'he4 == _GEN_13581 ? ~tag_compare_valid_1 : meta_228_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4846 = 8'he5 == _GEN_13581 ? ~tag_compare_valid_1 : meta_229_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4847 = 8'he6 == _GEN_13581 ? ~tag_compare_valid_1 : meta_230_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4848 = 8'he7 == _GEN_13581 ? ~tag_compare_valid_1 : meta_231_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4849 = 8'he8 == _GEN_13581 ? ~tag_compare_valid_1 : meta_232_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4850 = 8'he9 == _GEN_13581 ? ~tag_compare_valid_1 : meta_233_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4851 = 8'hea == _GEN_13581 ? ~tag_compare_valid_1 : meta_234_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4852 = 8'heb == _GEN_13581 ? ~tag_compare_valid_1 : meta_235_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4853 = 8'hec == _GEN_13581 ? ~tag_compare_valid_1 : meta_236_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4854 = 8'hed == _GEN_13581 ? ~tag_compare_valid_1 : meta_237_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4855 = 8'hee == _GEN_13581 ? ~tag_compare_valid_1 : meta_238_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4856 = 8'hef == _GEN_13581 ? ~tag_compare_valid_1 : meta_239_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4857 = 8'hf0 == _GEN_13581 ? ~tag_compare_valid_1 : meta_240_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4858 = 8'hf1 == _GEN_13581 ? ~tag_compare_valid_1 : meta_241_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4859 = 8'hf2 == _GEN_13581 ? ~tag_compare_valid_1 : meta_242_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4860 = 8'hf3 == _GEN_13581 ? ~tag_compare_valid_1 : meta_243_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4861 = 8'hf4 == _GEN_13581 ? ~tag_compare_valid_1 : meta_244_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4862 = 8'hf5 == _GEN_13581 ? ~tag_compare_valid_1 : meta_245_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4863 = 8'hf6 == _GEN_13581 ? ~tag_compare_valid_1 : meta_246_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4864 = 8'hf7 == _GEN_13581 ? ~tag_compare_valid_1 : meta_247_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4865 = 8'hf8 == _GEN_13581 ? ~tag_compare_valid_1 : meta_248_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4866 = 8'hf9 == _GEN_13581 ? ~tag_compare_valid_1 : meta_249_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4867 = 8'hfa == _GEN_13581 ? ~tag_compare_valid_1 : meta_250_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4868 = 8'hfb == _GEN_13581 ? ~tag_compare_valid_1 : meta_251_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4869 = 8'hfc == _GEN_13581 ? ~tag_compare_valid_1 : meta_252_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4870 = 8'hfd == _GEN_13581 ? ~tag_compare_valid_1 : meta_253_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4871 = 8'hfe == _GEN_13581 ? ~tag_compare_valid_1 : meta_254_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4872 = 8'hff == _GEN_13581 ? ~tag_compare_valid_1 : meta_255_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4873 = 9'h100 == _GEN_13709 ? ~tag_compare_valid_1 : meta_256_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4874 = 9'h101 == _GEN_13709 ? ~tag_compare_valid_1 : meta_257_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4875 = 9'h102 == _GEN_13709 ? ~tag_compare_valid_1 : meta_258_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4876 = 9'h103 == _GEN_13709 ? ~tag_compare_valid_1 : meta_259_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4877 = 9'h104 == _GEN_13709 ? ~tag_compare_valid_1 : meta_260_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4878 = 9'h105 == _GEN_13709 ? ~tag_compare_valid_1 : meta_261_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4879 = 9'h106 == _GEN_13709 ? ~tag_compare_valid_1 : meta_262_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4880 = 9'h107 == _GEN_13709 ? ~tag_compare_valid_1 : meta_263_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4881 = 9'h108 == _GEN_13709 ? ~tag_compare_valid_1 : meta_264_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4882 = 9'h109 == _GEN_13709 ? ~tag_compare_valid_1 : meta_265_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4883 = 9'h10a == _GEN_13709 ? ~tag_compare_valid_1 : meta_266_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4884 = 9'h10b == _GEN_13709 ? ~tag_compare_valid_1 : meta_267_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4885 = 9'h10c == _GEN_13709 ? ~tag_compare_valid_1 : meta_268_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4886 = 9'h10d == _GEN_13709 ? ~tag_compare_valid_1 : meta_269_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4887 = 9'h10e == _GEN_13709 ? ~tag_compare_valid_1 : meta_270_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4888 = 9'h10f == _GEN_13709 ? ~tag_compare_valid_1 : meta_271_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4889 = 9'h110 == _GEN_13709 ? ~tag_compare_valid_1 : meta_272_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4890 = 9'h111 == _GEN_13709 ? ~tag_compare_valid_1 : meta_273_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4891 = 9'h112 == _GEN_13709 ? ~tag_compare_valid_1 : meta_274_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4892 = 9'h113 == _GEN_13709 ? ~tag_compare_valid_1 : meta_275_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4893 = 9'h114 == _GEN_13709 ? ~tag_compare_valid_1 : meta_276_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4894 = 9'h115 == _GEN_13709 ? ~tag_compare_valid_1 : meta_277_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4895 = 9'h116 == _GEN_13709 ? ~tag_compare_valid_1 : meta_278_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4896 = 9'h117 == _GEN_13709 ? ~tag_compare_valid_1 : meta_279_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4897 = 9'h118 == _GEN_13709 ? ~tag_compare_valid_1 : meta_280_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4898 = 9'h119 == _GEN_13709 ? ~tag_compare_valid_1 : meta_281_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4899 = 9'h11a == _GEN_13709 ? ~tag_compare_valid_1 : meta_282_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4900 = 9'h11b == _GEN_13709 ? ~tag_compare_valid_1 : meta_283_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4901 = 9'h11c == _GEN_13709 ? ~tag_compare_valid_1 : meta_284_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4902 = 9'h11d == _GEN_13709 ? ~tag_compare_valid_1 : meta_285_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4903 = 9'h11e == _GEN_13709 ? ~tag_compare_valid_1 : meta_286_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4904 = 9'h11f == _GEN_13709 ? ~tag_compare_valid_1 : meta_287_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4905 = 9'h120 == _GEN_13709 ? ~tag_compare_valid_1 : meta_288_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4906 = 9'h121 == _GEN_13709 ? ~tag_compare_valid_1 : meta_289_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4907 = 9'h122 == _GEN_13709 ? ~tag_compare_valid_1 : meta_290_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4908 = 9'h123 == _GEN_13709 ? ~tag_compare_valid_1 : meta_291_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4909 = 9'h124 == _GEN_13709 ? ~tag_compare_valid_1 : meta_292_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4910 = 9'h125 == _GEN_13709 ? ~tag_compare_valid_1 : meta_293_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4911 = 9'h126 == _GEN_13709 ? ~tag_compare_valid_1 : meta_294_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4912 = 9'h127 == _GEN_13709 ? ~tag_compare_valid_1 : meta_295_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4913 = 9'h128 == _GEN_13709 ? ~tag_compare_valid_1 : meta_296_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4914 = 9'h129 == _GEN_13709 ? ~tag_compare_valid_1 : meta_297_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4915 = 9'h12a == _GEN_13709 ? ~tag_compare_valid_1 : meta_298_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4916 = 9'h12b == _GEN_13709 ? ~tag_compare_valid_1 : meta_299_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4917 = 9'h12c == _GEN_13709 ? ~tag_compare_valid_1 : meta_300_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4918 = 9'h12d == _GEN_13709 ? ~tag_compare_valid_1 : meta_301_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4919 = 9'h12e == _GEN_13709 ? ~tag_compare_valid_1 : meta_302_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4920 = 9'h12f == _GEN_13709 ? ~tag_compare_valid_1 : meta_303_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4921 = 9'h130 == _GEN_13709 ? ~tag_compare_valid_1 : meta_304_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4922 = 9'h131 == _GEN_13709 ? ~tag_compare_valid_1 : meta_305_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4923 = 9'h132 == _GEN_13709 ? ~tag_compare_valid_1 : meta_306_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4924 = 9'h133 == _GEN_13709 ? ~tag_compare_valid_1 : meta_307_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4925 = 9'h134 == _GEN_13709 ? ~tag_compare_valid_1 : meta_308_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4926 = 9'h135 == _GEN_13709 ? ~tag_compare_valid_1 : meta_309_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4927 = 9'h136 == _GEN_13709 ? ~tag_compare_valid_1 : meta_310_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4928 = 9'h137 == _GEN_13709 ? ~tag_compare_valid_1 : meta_311_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4929 = 9'h138 == _GEN_13709 ? ~tag_compare_valid_1 : meta_312_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4930 = 9'h139 == _GEN_13709 ? ~tag_compare_valid_1 : meta_313_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4931 = 9'h13a == _GEN_13709 ? ~tag_compare_valid_1 : meta_314_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4932 = 9'h13b == _GEN_13709 ? ~tag_compare_valid_1 : meta_315_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4933 = 9'h13c == _GEN_13709 ? ~tag_compare_valid_1 : meta_316_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4934 = 9'h13d == _GEN_13709 ? ~tag_compare_valid_1 : meta_317_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4935 = 9'h13e == _GEN_13709 ? ~tag_compare_valid_1 : meta_318_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4936 = 9'h13f == _GEN_13709 ? ~tag_compare_valid_1 : meta_319_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4937 = 9'h140 == _GEN_13709 ? ~tag_compare_valid_1 : meta_320_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4938 = 9'h141 == _GEN_13709 ? ~tag_compare_valid_1 : meta_321_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4939 = 9'h142 == _GEN_13709 ? ~tag_compare_valid_1 : meta_322_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4940 = 9'h143 == _GEN_13709 ? ~tag_compare_valid_1 : meta_323_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4941 = 9'h144 == _GEN_13709 ? ~tag_compare_valid_1 : meta_324_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4942 = 9'h145 == _GEN_13709 ? ~tag_compare_valid_1 : meta_325_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4943 = 9'h146 == _GEN_13709 ? ~tag_compare_valid_1 : meta_326_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4944 = 9'h147 == _GEN_13709 ? ~tag_compare_valid_1 : meta_327_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4945 = 9'h148 == _GEN_13709 ? ~tag_compare_valid_1 : meta_328_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4946 = 9'h149 == _GEN_13709 ? ~tag_compare_valid_1 : meta_329_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4947 = 9'h14a == _GEN_13709 ? ~tag_compare_valid_1 : meta_330_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4948 = 9'h14b == _GEN_13709 ? ~tag_compare_valid_1 : meta_331_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4949 = 9'h14c == _GEN_13709 ? ~tag_compare_valid_1 : meta_332_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4950 = 9'h14d == _GEN_13709 ? ~tag_compare_valid_1 : meta_333_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4951 = 9'h14e == _GEN_13709 ? ~tag_compare_valid_1 : meta_334_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4952 = 9'h14f == _GEN_13709 ? ~tag_compare_valid_1 : meta_335_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4953 = 9'h150 == _GEN_13709 ? ~tag_compare_valid_1 : meta_336_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4954 = 9'h151 == _GEN_13709 ? ~tag_compare_valid_1 : meta_337_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4955 = 9'h152 == _GEN_13709 ? ~tag_compare_valid_1 : meta_338_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4956 = 9'h153 == _GEN_13709 ? ~tag_compare_valid_1 : meta_339_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4957 = 9'h154 == _GEN_13709 ? ~tag_compare_valid_1 : meta_340_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4958 = 9'h155 == _GEN_13709 ? ~tag_compare_valid_1 : meta_341_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4959 = 9'h156 == _GEN_13709 ? ~tag_compare_valid_1 : meta_342_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4960 = 9'h157 == _GEN_13709 ? ~tag_compare_valid_1 : meta_343_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4961 = 9'h158 == _GEN_13709 ? ~tag_compare_valid_1 : meta_344_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4962 = 9'h159 == _GEN_13709 ? ~tag_compare_valid_1 : meta_345_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4963 = 9'h15a == _GEN_13709 ? ~tag_compare_valid_1 : meta_346_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4964 = 9'h15b == _GEN_13709 ? ~tag_compare_valid_1 : meta_347_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4965 = 9'h15c == _GEN_13709 ? ~tag_compare_valid_1 : meta_348_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4966 = 9'h15d == _GEN_13709 ? ~tag_compare_valid_1 : meta_349_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4967 = 9'h15e == _GEN_13709 ? ~tag_compare_valid_1 : meta_350_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4968 = 9'h15f == _GEN_13709 ? ~tag_compare_valid_1 : meta_351_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4969 = 9'h160 == _GEN_13709 ? ~tag_compare_valid_1 : meta_352_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4970 = 9'h161 == _GEN_13709 ? ~tag_compare_valid_1 : meta_353_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4971 = 9'h162 == _GEN_13709 ? ~tag_compare_valid_1 : meta_354_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4972 = 9'h163 == _GEN_13709 ? ~tag_compare_valid_1 : meta_355_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4973 = 9'h164 == _GEN_13709 ? ~tag_compare_valid_1 : meta_356_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4974 = 9'h165 == _GEN_13709 ? ~tag_compare_valid_1 : meta_357_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4975 = 9'h166 == _GEN_13709 ? ~tag_compare_valid_1 : meta_358_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4976 = 9'h167 == _GEN_13709 ? ~tag_compare_valid_1 : meta_359_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4977 = 9'h168 == _GEN_13709 ? ~tag_compare_valid_1 : meta_360_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4978 = 9'h169 == _GEN_13709 ? ~tag_compare_valid_1 : meta_361_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4979 = 9'h16a == _GEN_13709 ? ~tag_compare_valid_1 : meta_362_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4980 = 9'h16b == _GEN_13709 ? ~tag_compare_valid_1 : meta_363_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4981 = 9'h16c == _GEN_13709 ? ~tag_compare_valid_1 : meta_364_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4982 = 9'h16d == _GEN_13709 ? ~tag_compare_valid_1 : meta_365_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4983 = 9'h16e == _GEN_13709 ? ~tag_compare_valid_1 : meta_366_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4984 = 9'h16f == _GEN_13709 ? ~tag_compare_valid_1 : meta_367_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4985 = 9'h170 == _GEN_13709 ? ~tag_compare_valid_1 : meta_368_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4986 = 9'h171 == _GEN_13709 ? ~tag_compare_valid_1 : meta_369_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4987 = 9'h172 == _GEN_13709 ? ~tag_compare_valid_1 : meta_370_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4988 = 9'h173 == _GEN_13709 ? ~tag_compare_valid_1 : meta_371_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4989 = 9'h174 == _GEN_13709 ? ~tag_compare_valid_1 : meta_372_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4990 = 9'h175 == _GEN_13709 ? ~tag_compare_valid_1 : meta_373_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4991 = 9'h176 == _GEN_13709 ? ~tag_compare_valid_1 : meta_374_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4992 = 9'h177 == _GEN_13709 ? ~tag_compare_valid_1 : meta_375_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4993 = 9'h178 == _GEN_13709 ? ~tag_compare_valid_1 : meta_376_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4994 = 9'h179 == _GEN_13709 ? ~tag_compare_valid_1 : meta_377_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4995 = 9'h17a == _GEN_13709 ? ~tag_compare_valid_1 : meta_378_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4996 = 9'h17b == _GEN_13709 ? ~tag_compare_valid_1 : meta_379_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4997 = 9'h17c == _GEN_13709 ? ~tag_compare_valid_1 : meta_380_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4998 = 9'h17d == _GEN_13709 ? ~tag_compare_valid_1 : meta_381_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_4999 = 9'h17e == _GEN_13709 ? ~tag_compare_valid_1 : meta_382_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5000 = 9'h17f == _GEN_13709 ? ~tag_compare_valid_1 : meta_383_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5001 = 9'h180 == _GEN_13709 ? ~tag_compare_valid_1 : meta_384_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5002 = 9'h181 == _GEN_13709 ? ~tag_compare_valid_1 : meta_385_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5003 = 9'h182 == _GEN_13709 ? ~tag_compare_valid_1 : meta_386_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5004 = 9'h183 == _GEN_13709 ? ~tag_compare_valid_1 : meta_387_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5005 = 9'h184 == _GEN_13709 ? ~tag_compare_valid_1 : meta_388_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5006 = 9'h185 == _GEN_13709 ? ~tag_compare_valid_1 : meta_389_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5007 = 9'h186 == _GEN_13709 ? ~tag_compare_valid_1 : meta_390_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5008 = 9'h187 == _GEN_13709 ? ~tag_compare_valid_1 : meta_391_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5009 = 9'h188 == _GEN_13709 ? ~tag_compare_valid_1 : meta_392_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5010 = 9'h189 == _GEN_13709 ? ~tag_compare_valid_1 : meta_393_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5011 = 9'h18a == _GEN_13709 ? ~tag_compare_valid_1 : meta_394_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5012 = 9'h18b == _GEN_13709 ? ~tag_compare_valid_1 : meta_395_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5013 = 9'h18c == _GEN_13709 ? ~tag_compare_valid_1 : meta_396_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5014 = 9'h18d == _GEN_13709 ? ~tag_compare_valid_1 : meta_397_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5015 = 9'h18e == _GEN_13709 ? ~tag_compare_valid_1 : meta_398_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5016 = 9'h18f == _GEN_13709 ? ~tag_compare_valid_1 : meta_399_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5017 = 9'h190 == _GEN_13709 ? ~tag_compare_valid_1 : meta_400_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5018 = 9'h191 == _GEN_13709 ? ~tag_compare_valid_1 : meta_401_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5019 = 9'h192 == _GEN_13709 ? ~tag_compare_valid_1 : meta_402_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5020 = 9'h193 == _GEN_13709 ? ~tag_compare_valid_1 : meta_403_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5021 = 9'h194 == _GEN_13709 ? ~tag_compare_valid_1 : meta_404_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5022 = 9'h195 == _GEN_13709 ? ~tag_compare_valid_1 : meta_405_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5023 = 9'h196 == _GEN_13709 ? ~tag_compare_valid_1 : meta_406_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5024 = 9'h197 == _GEN_13709 ? ~tag_compare_valid_1 : meta_407_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5025 = 9'h198 == _GEN_13709 ? ~tag_compare_valid_1 : meta_408_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5026 = 9'h199 == _GEN_13709 ? ~tag_compare_valid_1 : meta_409_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5027 = 9'h19a == _GEN_13709 ? ~tag_compare_valid_1 : meta_410_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5028 = 9'h19b == _GEN_13709 ? ~tag_compare_valid_1 : meta_411_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5029 = 9'h19c == _GEN_13709 ? ~tag_compare_valid_1 : meta_412_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5030 = 9'h19d == _GEN_13709 ? ~tag_compare_valid_1 : meta_413_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5031 = 9'h19e == _GEN_13709 ? ~tag_compare_valid_1 : meta_414_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5032 = 9'h19f == _GEN_13709 ? ~tag_compare_valid_1 : meta_415_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5033 = 9'h1a0 == _GEN_13709 ? ~tag_compare_valid_1 : meta_416_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5034 = 9'h1a1 == _GEN_13709 ? ~tag_compare_valid_1 : meta_417_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5035 = 9'h1a2 == _GEN_13709 ? ~tag_compare_valid_1 : meta_418_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5036 = 9'h1a3 == _GEN_13709 ? ~tag_compare_valid_1 : meta_419_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5037 = 9'h1a4 == _GEN_13709 ? ~tag_compare_valid_1 : meta_420_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5038 = 9'h1a5 == _GEN_13709 ? ~tag_compare_valid_1 : meta_421_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5039 = 9'h1a6 == _GEN_13709 ? ~tag_compare_valid_1 : meta_422_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5040 = 9'h1a7 == _GEN_13709 ? ~tag_compare_valid_1 : meta_423_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5041 = 9'h1a8 == _GEN_13709 ? ~tag_compare_valid_1 : meta_424_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5042 = 9'h1a9 == _GEN_13709 ? ~tag_compare_valid_1 : meta_425_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5043 = 9'h1aa == _GEN_13709 ? ~tag_compare_valid_1 : meta_426_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5044 = 9'h1ab == _GEN_13709 ? ~tag_compare_valid_1 : meta_427_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5045 = 9'h1ac == _GEN_13709 ? ~tag_compare_valid_1 : meta_428_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5046 = 9'h1ad == _GEN_13709 ? ~tag_compare_valid_1 : meta_429_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5047 = 9'h1ae == _GEN_13709 ? ~tag_compare_valid_1 : meta_430_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5048 = 9'h1af == _GEN_13709 ? ~tag_compare_valid_1 : meta_431_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5049 = 9'h1b0 == _GEN_13709 ? ~tag_compare_valid_1 : meta_432_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5050 = 9'h1b1 == _GEN_13709 ? ~tag_compare_valid_1 : meta_433_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5051 = 9'h1b2 == _GEN_13709 ? ~tag_compare_valid_1 : meta_434_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5052 = 9'h1b3 == _GEN_13709 ? ~tag_compare_valid_1 : meta_435_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5053 = 9'h1b4 == _GEN_13709 ? ~tag_compare_valid_1 : meta_436_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5054 = 9'h1b5 == _GEN_13709 ? ~tag_compare_valid_1 : meta_437_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5055 = 9'h1b6 == _GEN_13709 ? ~tag_compare_valid_1 : meta_438_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5056 = 9'h1b7 == _GEN_13709 ? ~tag_compare_valid_1 : meta_439_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5057 = 9'h1b8 == _GEN_13709 ? ~tag_compare_valid_1 : meta_440_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5058 = 9'h1b9 == _GEN_13709 ? ~tag_compare_valid_1 : meta_441_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5059 = 9'h1ba == _GEN_13709 ? ~tag_compare_valid_1 : meta_442_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5060 = 9'h1bb == _GEN_13709 ? ~tag_compare_valid_1 : meta_443_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5061 = 9'h1bc == _GEN_13709 ? ~tag_compare_valid_1 : meta_444_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5062 = 9'h1bd == _GEN_13709 ? ~tag_compare_valid_1 : meta_445_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5063 = 9'h1be == _GEN_13709 ? ~tag_compare_valid_1 : meta_446_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5064 = 9'h1bf == _GEN_13709 ? ~tag_compare_valid_1 : meta_447_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5065 = 9'h1c0 == _GEN_13709 ? ~tag_compare_valid_1 : meta_448_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5066 = 9'h1c1 == _GEN_13709 ? ~tag_compare_valid_1 : meta_449_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5067 = 9'h1c2 == _GEN_13709 ? ~tag_compare_valid_1 : meta_450_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5068 = 9'h1c3 == _GEN_13709 ? ~tag_compare_valid_1 : meta_451_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5069 = 9'h1c4 == _GEN_13709 ? ~tag_compare_valid_1 : meta_452_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5070 = 9'h1c5 == _GEN_13709 ? ~tag_compare_valid_1 : meta_453_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5071 = 9'h1c6 == _GEN_13709 ? ~tag_compare_valid_1 : meta_454_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5072 = 9'h1c7 == _GEN_13709 ? ~tag_compare_valid_1 : meta_455_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5073 = 9'h1c8 == _GEN_13709 ? ~tag_compare_valid_1 : meta_456_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5074 = 9'h1c9 == _GEN_13709 ? ~tag_compare_valid_1 : meta_457_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5075 = 9'h1ca == _GEN_13709 ? ~tag_compare_valid_1 : meta_458_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5076 = 9'h1cb == _GEN_13709 ? ~tag_compare_valid_1 : meta_459_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5077 = 9'h1cc == _GEN_13709 ? ~tag_compare_valid_1 : meta_460_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5078 = 9'h1cd == _GEN_13709 ? ~tag_compare_valid_1 : meta_461_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5079 = 9'h1ce == _GEN_13709 ? ~tag_compare_valid_1 : meta_462_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5080 = 9'h1cf == _GEN_13709 ? ~tag_compare_valid_1 : meta_463_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5081 = 9'h1d0 == _GEN_13709 ? ~tag_compare_valid_1 : meta_464_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5082 = 9'h1d1 == _GEN_13709 ? ~tag_compare_valid_1 : meta_465_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5083 = 9'h1d2 == _GEN_13709 ? ~tag_compare_valid_1 : meta_466_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5084 = 9'h1d3 == _GEN_13709 ? ~tag_compare_valid_1 : meta_467_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5085 = 9'h1d4 == _GEN_13709 ? ~tag_compare_valid_1 : meta_468_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5086 = 9'h1d5 == _GEN_13709 ? ~tag_compare_valid_1 : meta_469_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5087 = 9'h1d6 == _GEN_13709 ? ~tag_compare_valid_1 : meta_470_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5088 = 9'h1d7 == _GEN_13709 ? ~tag_compare_valid_1 : meta_471_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5089 = 9'h1d8 == _GEN_13709 ? ~tag_compare_valid_1 : meta_472_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5090 = 9'h1d9 == _GEN_13709 ? ~tag_compare_valid_1 : meta_473_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5091 = 9'h1da == _GEN_13709 ? ~tag_compare_valid_1 : meta_474_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5092 = 9'h1db == _GEN_13709 ? ~tag_compare_valid_1 : meta_475_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5093 = 9'h1dc == _GEN_13709 ? ~tag_compare_valid_1 : meta_476_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5094 = 9'h1dd == _GEN_13709 ? ~tag_compare_valid_1 : meta_477_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5095 = 9'h1de == _GEN_13709 ? ~tag_compare_valid_1 : meta_478_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5096 = 9'h1df == _GEN_13709 ? ~tag_compare_valid_1 : meta_479_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5097 = 9'h1e0 == _GEN_13709 ? ~tag_compare_valid_1 : meta_480_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5098 = 9'h1e1 == _GEN_13709 ? ~tag_compare_valid_1 : meta_481_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5099 = 9'h1e2 == _GEN_13709 ? ~tag_compare_valid_1 : meta_482_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5100 = 9'h1e3 == _GEN_13709 ? ~tag_compare_valid_1 : meta_483_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5101 = 9'h1e4 == _GEN_13709 ? ~tag_compare_valid_1 : meta_484_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5102 = 9'h1e5 == _GEN_13709 ? ~tag_compare_valid_1 : meta_485_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5103 = 9'h1e6 == _GEN_13709 ? ~tag_compare_valid_1 : meta_486_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5104 = 9'h1e7 == _GEN_13709 ? ~tag_compare_valid_1 : meta_487_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5105 = 9'h1e8 == _GEN_13709 ? ~tag_compare_valid_1 : meta_488_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5106 = 9'h1e9 == _GEN_13709 ? ~tag_compare_valid_1 : meta_489_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5107 = 9'h1ea == _GEN_13709 ? ~tag_compare_valid_1 : meta_490_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5108 = 9'h1eb == _GEN_13709 ? ~tag_compare_valid_1 : meta_491_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5109 = 9'h1ec == _GEN_13709 ? ~tag_compare_valid_1 : meta_492_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5110 = 9'h1ed == _GEN_13709 ? ~tag_compare_valid_1 : meta_493_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5111 = 9'h1ee == _GEN_13709 ? ~tag_compare_valid_1 : meta_494_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5112 = 9'h1ef == _GEN_13709 ? ~tag_compare_valid_1 : meta_495_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5113 = 9'h1f0 == _GEN_13709 ? ~tag_compare_valid_1 : meta_496_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5114 = 9'h1f1 == _GEN_13709 ? ~tag_compare_valid_1 : meta_497_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5115 = 9'h1f2 == _GEN_13709 ? ~tag_compare_valid_1 : meta_498_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5116 = 9'h1f3 == _GEN_13709 ? ~tag_compare_valid_1 : meta_499_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5117 = 9'h1f4 == _GEN_13709 ? ~tag_compare_valid_1 : meta_500_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5118 = 9'h1f5 == _GEN_13709 ? ~tag_compare_valid_1 : meta_501_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5119 = 9'h1f6 == _GEN_13709 ? ~tag_compare_valid_1 : meta_502_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5120 = 9'h1f7 == _GEN_13709 ? ~tag_compare_valid_1 : meta_503_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5121 = 9'h1f8 == _GEN_13709 ? ~tag_compare_valid_1 : meta_504_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5122 = 9'h1f9 == _GEN_13709 ? ~tag_compare_valid_1 : meta_505_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5123 = 9'h1fa == _GEN_13709 ? ~tag_compare_valid_1 : meta_506_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5124 = 9'h1fb == _GEN_13709 ? ~tag_compare_valid_1 : meta_507_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5125 = 9'h1fc == _GEN_13709 ? ~tag_compare_valid_1 : meta_508_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5126 = 9'h1fd == _GEN_13709 ? ~tag_compare_valid_1 : meta_509_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5127 = 9'h1fe == _GEN_13709 ? ~tag_compare_valid_1 : meta_510_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire  _GEN_5128 = 9'h1ff == _GEN_13709 ? ~tag_compare_valid_1 : meta_511_lru; // @[ICache.scala 189:{34,34} 34:21]
  wire [2:0] _GEN_5129 = io_cpu_cpu_stall ? 3'h4 : state; // @[ICache.scala 190:34 191:28 48:81]
  wire [63:0] _GEN_5130 = io_cpu_cpu_stall ? cache_data_1 : {{32'd0}, saved_1_inst}; // @[ICache.scala 190:34 192:28 91:22]
  wire  _GEN_5131 = io_cpu_cpu_stall ? cache_hit_available : saved_0_valid; // @[ICache.scala 190:34 193:28 91:22]
  wire  _GEN_5132 = io_cpu_cpu_stall ? cache_inst_ok_1 : saved_1_valid; // @[ICache.scala 190:34 194:28 91:22]
  wire  _GEN_5133 = _T ? _GEN_4617 : meta_0_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5134 = _T ? _GEN_4618 : meta_1_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5135 = _T ? _GEN_4619 : meta_2_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5136 = _T ? _GEN_4620 : meta_3_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5137 = _T ? _GEN_4621 : meta_4_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5138 = _T ? _GEN_4622 : meta_5_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5139 = _T ? _GEN_4623 : meta_6_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5140 = _T ? _GEN_4624 : meta_7_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5141 = _T ? _GEN_4625 : meta_8_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5142 = _T ? _GEN_4626 : meta_9_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5143 = _T ? _GEN_4627 : meta_10_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5144 = _T ? _GEN_4628 : meta_11_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5145 = _T ? _GEN_4629 : meta_12_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5146 = _T ? _GEN_4630 : meta_13_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5147 = _T ? _GEN_4631 : meta_14_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5148 = _T ? _GEN_4632 : meta_15_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5149 = _T ? _GEN_4633 : meta_16_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5150 = _T ? _GEN_4634 : meta_17_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5151 = _T ? _GEN_4635 : meta_18_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5152 = _T ? _GEN_4636 : meta_19_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5153 = _T ? _GEN_4637 : meta_20_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5154 = _T ? _GEN_4638 : meta_21_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5155 = _T ? _GEN_4639 : meta_22_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5156 = _T ? _GEN_4640 : meta_23_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5157 = _T ? _GEN_4641 : meta_24_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5158 = _T ? _GEN_4642 : meta_25_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5159 = _T ? _GEN_4643 : meta_26_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5160 = _T ? _GEN_4644 : meta_27_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5161 = _T ? _GEN_4645 : meta_28_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5162 = _T ? _GEN_4646 : meta_29_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5163 = _T ? _GEN_4647 : meta_30_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5164 = _T ? _GEN_4648 : meta_31_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5165 = _T ? _GEN_4649 : meta_32_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5166 = _T ? _GEN_4650 : meta_33_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5167 = _T ? _GEN_4651 : meta_34_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5168 = _T ? _GEN_4652 : meta_35_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5169 = _T ? _GEN_4653 : meta_36_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5170 = _T ? _GEN_4654 : meta_37_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5171 = _T ? _GEN_4655 : meta_38_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5172 = _T ? _GEN_4656 : meta_39_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5173 = _T ? _GEN_4657 : meta_40_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5174 = _T ? _GEN_4658 : meta_41_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5175 = _T ? _GEN_4659 : meta_42_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5176 = _T ? _GEN_4660 : meta_43_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5177 = _T ? _GEN_4661 : meta_44_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5178 = _T ? _GEN_4662 : meta_45_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5179 = _T ? _GEN_4663 : meta_46_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5180 = _T ? _GEN_4664 : meta_47_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5181 = _T ? _GEN_4665 : meta_48_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5182 = _T ? _GEN_4666 : meta_49_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5183 = _T ? _GEN_4667 : meta_50_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5184 = _T ? _GEN_4668 : meta_51_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5185 = _T ? _GEN_4669 : meta_52_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5186 = _T ? _GEN_4670 : meta_53_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5187 = _T ? _GEN_4671 : meta_54_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5188 = _T ? _GEN_4672 : meta_55_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5189 = _T ? _GEN_4673 : meta_56_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5190 = _T ? _GEN_4674 : meta_57_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5191 = _T ? _GEN_4675 : meta_58_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5192 = _T ? _GEN_4676 : meta_59_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5193 = _T ? _GEN_4677 : meta_60_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5194 = _T ? _GEN_4678 : meta_61_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5195 = _T ? _GEN_4679 : meta_62_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5196 = _T ? _GEN_4680 : meta_63_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5197 = _T ? _GEN_4681 : meta_64_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5198 = _T ? _GEN_4682 : meta_65_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5199 = _T ? _GEN_4683 : meta_66_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5200 = _T ? _GEN_4684 : meta_67_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5201 = _T ? _GEN_4685 : meta_68_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5202 = _T ? _GEN_4686 : meta_69_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5203 = _T ? _GEN_4687 : meta_70_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5204 = _T ? _GEN_4688 : meta_71_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5205 = _T ? _GEN_4689 : meta_72_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5206 = _T ? _GEN_4690 : meta_73_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5207 = _T ? _GEN_4691 : meta_74_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5208 = _T ? _GEN_4692 : meta_75_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5209 = _T ? _GEN_4693 : meta_76_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5210 = _T ? _GEN_4694 : meta_77_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5211 = _T ? _GEN_4695 : meta_78_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5212 = _T ? _GEN_4696 : meta_79_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5213 = _T ? _GEN_4697 : meta_80_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5214 = _T ? _GEN_4698 : meta_81_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5215 = _T ? _GEN_4699 : meta_82_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5216 = _T ? _GEN_4700 : meta_83_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5217 = _T ? _GEN_4701 : meta_84_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5218 = _T ? _GEN_4702 : meta_85_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5219 = _T ? _GEN_4703 : meta_86_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5220 = _T ? _GEN_4704 : meta_87_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5221 = _T ? _GEN_4705 : meta_88_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5222 = _T ? _GEN_4706 : meta_89_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5223 = _T ? _GEN_4707 : meta_90_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5224 = _T ? _GEN_4708 : meta_91_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5225 = _T ? _GEN_4709 : meta_92_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5226 = _T ? _GEN_4710 : meta_93_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5227 = _T ? _GEN_4711 : meta_94_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5228 = _T ? _GEN_4712 : meta_95_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5229 = _T ? _GEN_4713 : meta_96_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5230 = _T ? _GEN_4714 : meta_97_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5231 = _T ? _GEN_4715 : meta_98_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5232 = _T ? _GEN_4716 : meta_99_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5233 = _T ? _GEN_4717 : meta_100_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5234 = _T ? _GEN_4718 : meta_101_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5235 = _T ? _GEN_4719 : meta_102_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5236 = _T ? _GEN_4720 : meta_103_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5237 = _T ? _GEN_4721 : meta_104_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5238 = _T ? _GEN_4722 : meta_105_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5239 = _T ? _GEN_4723 : meta_106_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5240 = _T ? _GEN_4724 : meta_107_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5241 = _T ? _GEN_4725 : meta_108_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5242 = _T ? _GEN_4726 : meta_109_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5243 = _T ? _GEN_4727 : meta_110_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5244 = _T ? _GEN_4728 : meta_111_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5245 = _T ? _GEN_4729 : meta_112_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5246 = _T ? _GEN_4730 : meta_113_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5247 = _T ? _GEN_4731 : meta_114_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5248 = _T ? _GEN_4732 : meta_115_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5249 = _T ? _GEN_4733 : meta_116_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5250 = _T ? _GEN_4734 : meta_117_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5251 = _T ? _GEN_4735 : meta_118_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5252 = _T ? _GEN_4736 : meta_119_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5253 = _T ? _GEN_4737 : meta_120_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5254 = _T ? _GEN_4738 : meta_121_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5255 = _T ? _GEN_4739 : meta_122_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5256 = _T ? _GEN_4740 : meta_123_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5257 = _T ? _GEN_4741 : meta_124_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5258 = _T ? _GEN_4742 : meta_125_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5259 = _T ? _GEN_4743 : meta_126_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5260 = _T ? _GEN_4744 : meta_127_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5261 = _T ? _GEN_4745 : meta_128_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5262 = _T ? _GEN_4746 : meta_129_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5263 = _T ? _GEN_4747 : meta_130_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5264 = _T ? _GEN_4748 : meta_131_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5265 = _T ? _GEN_4749 : meta_132_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5266 = _T ? _GEN_4750 : meta_133_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5267 = _T ? _GEN_4751 : meta_134_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5268 = _T ? _GEN_4752 : meta_135_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5269 = _T ? _GEN_4753 : meta_136_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5270 = _T ? _GEN_4754 : meta_137_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5271 = _T ? _GEN_4755 : meta_138_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5272 = _T ? _GEN_4756 : meta_139_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5273 = _T ? _GEN_4757 : meta_140_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5274 = _T ? _GEN_4758 : meta_141_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5275 = _T ? _GEN_4759 : meta_142_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5276 = _T ? _GEN_4760 : meta_143_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5277 = _T ? _GEN_4761 : meta_144_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5278 = _T ? _GEN_4762 : meta_145_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5279 = _T ? _GEN_4763 : meta_146_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5280 = _T ? _GEN_4764 : meta_147_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5281 = _T ? _GEN_4765 : meta_148_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5282 = _T ? _GEN_4766 : meta_149_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5283 = _T ? _GEN_4767 : meta_150_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5284 = _T ? _GEN_4768 : meta_151_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5285 = _T ? _GEN_4769 : meta_152_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5286 = _T ? _GEN_4770 : meta_153_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5287 = _T ? _GEN_4771 : meta_154_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5288 = _T ? _GEN_4772 : meta_155_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5289 = _T ? _GEN_4773 : meta_156_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5290 = _T ? _GEN_4774 : meta_157_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5291 = _T ? _GEN_4775 : meta_158_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5292 = _T ? _GEN_4776 : meta_159_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5293 = _T ? _GEN_4777 : meta_160_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5294 = _T ? _GEN_4778 : meta_161_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5295 = _T ? _GEN_4779 : meta_162_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5296 = _T ? _GEN_4780 : meta_163_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5297 = _T ? _GEN_4781 : meta_164_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5298 = _T ? _GEN_4782 : meta_165_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5299 = _T ? _GEN_4783 : meta_166_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5300 = _T ? _GEN_4784 : meta_167_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5301 = _T ? _GEN_4785 : meta_168_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5302 = _T ? _GEN_4786 : meta_169_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5303 = _T ? _GEN_4787 : meta_170_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5304 = _T ? _GEN_4788 : meta_171_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5305 = _T ? _GEN_4789 : meta_172_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5306 = _T ? _GEN_4790 : meta_173_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5307 = _T ? _GEN_4791 : meta_174_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5308 = _T ? _GEN_4792 : meta_175_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5309 = _T ? _GEN_4793 : meta_176_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5310 = _T ? _GEN_4794 : meta_177_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5311 = _T ? _GEN_4795 : meta_178_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5312 = _T ? _GEN_4796 : meta_179_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5313 = _T ? _GEN_4797 : meta_180_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5314 = _T ? _GEN_4798 : meta_181_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5315 = _T ? _GEN_4799 : meta_182_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5316 = _T ? _GEN_4800 : meta_183_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5317 = _T ? _GEN_4801 : meta_184_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5318 = _T ? _GEN_4802 : meta_185_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5319 = _T ? _GEN_4803 : meta_186_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5320 = _T ? _GEN_4804 : meta_187_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5321 = _T ? _GEN_4805 : meta_188_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5322 = _T ? _GEN_4806 : meta_189_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5323 = _T ? _GEN_4807 : meta_190_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5324 = _T ? _GEN_4808 : meta_191_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5325 = _T ? _GEN_4809 : meta_192_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5326 = _T ? _GEN_4810 : meta_193_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5327 = _T ? _GEN_4811 : meta_194_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5328 = _T ? _GEN_4812 : meta_195_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5329 = _T ? _GEN_4813 : meta_196_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5330 = _T ? _GEN_4814 : meta_197_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5331 = _T ? _GEN_4815 : meta_198_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5332 = _T ? _GEN_4816 : meta_199_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5333 = _T ? _GEN_4817 : meta_200_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5334 = _T ? _GEN_4818 : meta_201_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5335 = _T ? _GEN_4819 : meta_202_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5336 = _T ? _GEN_4820 : meta_203_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5337 = _T ? _GEN_4821 : meta_204_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5338 = _T ? _GEN_4822 : meta_205_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5339 = _T ? _GEN_4823 : meta_206_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5340 = _T ? _GEN_4824 : meta_207_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5341 = _T ? _GEN_4825 : meta_208_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5342 = _T ? _GEN_4826 : meta_209_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5343 = _T ? _GEN_4827 : meta_210_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5344 = _T ? _GEN_4828 : meta_211_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5345 = _T ? _GEN_4829 : meta_212_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5346 = _T ? _GEN_4830 : meta_213_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5347 = _T ? _GEN_4831 : meta_214_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5348 = _T ? _GEN_4832 : meta_215_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5349 = _T ? _GEN_4833 : meta_216_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5350 = _T ? _GEN_4834 : meta_217_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5351 = _T ? _GEN_4835 : meta_218_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5352 = _T ? _GEN_4836 : meta_219_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5353 = _T ? _GEN_4837 : meta_220_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5354 = _T ? _GEN_4838 : meta_221_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5355 = _T ? _GEN_4839 : meta_222_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5356 = _T ? _GEN_4840 : meta_223_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5357 = _T ? _GEN_4841 : meta_224_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5358 = _T ? _GEN_4842 : meta_225_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5359 = _T ? _GEN_4843 : meta_226_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5360 = _T ? _GEN_4844 : meta_227_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5361 = _T ? _GEN_4845 : meta_228_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5362 = _T ? _GEN_4846 : meta_229_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5363 = _T ? _GEN_4847 : meta_230_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5364 = _T ? _GEN_4848 : meta_231_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5365 = _T ? _GEN_4849 : meta_232_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5366 = _T ? _GEN_4850 : meta_233_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5367 = _T ? _GEN_4851 : meta_234_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5368 = _T ? _GEN_4852 : meta_235_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5369 = _T ? _GEN_4853 : meta_236_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5370 = _T ? _GEN_4854 : meta_237_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5371 = _T ? _GEN_4855 : meta_238_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5372 = _T ? _GEN_4856 : meta_239_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5373 = _T ? _GEN_4857 : meta_240_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5374 = _T ? _GEN_4858 : meta_241_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5375 = _T ? _GEN_4859 : meta_242_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5376 = _T ? _GEN_4860 : meta_243_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5377 = _T ? _GEN_4861 : meta_244_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5378 = _T ? _GEN_4862 : meta_245_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5379 = _T ? _GEN_4863 : meta_246_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5380 = _T ? _GEN_4864 : meta_247_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5381 = _T ? _GEN_4865 : meta_248_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5382 = _T ? _GEN_4866 : meta_249_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5383 = _T ? _GEN_4867 : meta_250_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5384 = _T ? _GEN_4868 : meta_251_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5385 = _T ? _GEN_4869 : meta_252_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5386 = _T ? _GEN_4870 : meta_253_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5387 = _T ? _GEN_4871 : meta_254_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5388 = _T ? _GEN_4872 : meta_255_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5389 = _T ? _GEN_4873 : meta_256_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5390 = _T ? _GEN_4874 : meta_257_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5391 = _T ? _GEN_4875 : meta_258_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5392 = _T ? _GEN_4876 : meta_259_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5393 = _T ? _GEN_4877 : meta_260_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5394 = _T ? _GEN_4878 : meta_261_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5395 = _T ? _GEN_4879 : meta_262_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5396 = _T ? _GEN_4880 : meta_263_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5397 = _T ? _GEN_4881 : meta_264_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5398 = _T ? _GEN_4882 : meta_265_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5399 = _T ? _GEN_4883 : meta_266_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5400 = _T ? _GEN_4884 : meta_267_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5401 = _T ? _GEN_4885 : meta_268_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5402 = _T ? _GEN_4886 : meta_269_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5403 = _T ? _GEN_4887 : meta_270_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5404 = _T ? _GEN_4888 : meta_271_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5405 = _T ? _GEN_4889 : meta_272_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5406 = _T ? _GEN_4890 : meta_273_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5407 = _T ? _GEN_4891 : meta_274_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5408 = _T ? _GEN_4892 : meta_275_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5409 = _T ? _GEN_4893 : meta_276_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5410 = _T ? _GEN_4894 : meta_277_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5411 = _T ? _GEN_4895 : meta_278_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5412 = _T ? _GEN_4896 : meta_279_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5413 = _T ? _GEN_4897 : meta_280_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5414 = _T ? _GEN_4898 : meta_281_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5415 = _T ? _GEN_4899 : meta_282_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5416 = _T ? _GEN_4900 : meta_283_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5417 = _T ? _GEN_4901 : meta_284_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5418 = _T ? _GEN_4902 : meta_285_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5419 = _T ? _GEN_4903 : meta_286_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5420 = _T ? _GEN_4904 : meta_287_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5421 = _T ? _GEN_4905 : meta_288_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5422 = _T ? _GEN_4906 : meta_289_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5423 = _T ? _GEN_4907 : meta_290_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5424 = _T ? _GEN_4908 : meta_291_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5425 = _T ? _GEN_4909 : meta_292_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5426 = _T ? _GEN_4910 : meta_293_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5427 = _T ? _GEN_4911 : meta_294_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5428 = _T ? _GEN_4912 : meta_295_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5429 = _T ? _GEN_4913 : meta_296_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5430 = _T ? _GEN_4914 : meta_297_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5431 = _T ? _GEN_4915 : meta_298_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5432 = _T ? _GEN_4916 : meta_299_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5433 = _T ? _GEN_4917 : meta_300_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5434 = _T ? _GEN_4918 : meta_301_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5435 = _T ? _GEN_4919 : meta_302_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5436 = _T ? _GEN_4920 : meta_303_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5437 = _T ? _GEN_4921 : meta_304_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5438 = _T ? _GEN_4922 : meta_305_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5439 = _T ? _GEN_4923 : meta_306_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5440 = _T ? _GEN_4924 : meta_307_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5441 = _T ? _GEN_4925 : meta_308_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5442 = _T ? _GEN_4926 : meta_309_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5443 = _T ? _GEN_4927 : meta_310_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5444 = _T ? _GEN_4928 : meta_311_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5445 = _T ? _GEN_4929 : meta_312_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5446 = _T ? _GEN_4930 : meta_313_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5447 = _T ? _GEN_4931 : meta_314_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5448 = _T ? _GEN_4932 : meta_315_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5449 = _T ? _GEN_4933 : meta_316_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5450 = _T ? _GEN_4934 : meta_317_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5451 = _T ? _GEN_4935 : meta_318_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5452 = _T ? _GEN_4936 : meta_319_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5453 = _T ? _GEN_4937 : meta_320_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5454 = _T ? _GEN_4938 : meta_321_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5455 = _T ? _GEN_4939 : meta_322_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5456 = _T ? _GEN_4940 : meta_323_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5457 = _T ? _GEN_4941 : meta_324_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5458 = _T ? _GEN_4942 : meta_325_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5459 = _T ? _GEN_4943 : meta_326_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5460 = _T ? _GEN_4944 : meta_327_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5461 = _T ? _GEN_4945 : meta_328_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5462 = _T ? _GEN_4946 : meta_329_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5463 = _T ? _GEN_4947 : meta_330_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5464 = _T ? _GEN_4948 : meta_331_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5465 = _T ? _GEN_4949 : meta_332_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5466 = _T ? _GEN_4950 : meta_333_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5467 = _T ? _GEN_4951 : meta_334_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5468 = _T ? _GEN_4952 : meta_335_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5469 = _T ? _GEN_4953 : meta_336_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5470 = _T ? _GEN_4954 : meta_337_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5471 = _T ? _GEN_4955 : meta_338_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5472 = _T ? _GEN_4956 : meta_339_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5473 = _T ? _GEN_4957 : meta_340_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5474 = _T ? _GEN_4958 : meta_341_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5475 = _T ? _GEN_4959 : meta_342_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5476 = _T ? _GEN_4960 : meta_343_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5477 = _T ? _GEN_4961 : meta_344_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5478 = _T ? _GEN_4962 : meta_345_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5479 = _T ? _GEN_4963 : meta_346_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5480 = _T ? _GEN_4964 : meta_347_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5481 = _T ? _GEN_4965 : meta_348_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5482 = _T ? _GEN_4966 : meta_349_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5483 = _T ? _GEN_4967 : meta_350_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5484 = _T ? _GEN_4968 : meta_351_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5485 = _T ? _GEN_4969 : meta_352_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5486 = _T ? _GEN_4970 : meta_353_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5487 = _T ? _GEN_4971 : meta_354_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5488 = _T ? _GEN_4972 : meta_355_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5489 = _T ? _GEN_4973 : meta_356_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5490 = _T ? _GEN_4974 : meta_357_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5491 = _T ? _GEN_4975 : meta_358_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5492 = _T ? _GEN_4976 : meta_359_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5493 = _T ? _GEN_4977 : meta_360_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5494 = _T ? _GEN_4978 : meta_361_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5495 = _T ? _GEN_4979 : meta_362_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5496 = _T ? _GEN_4980 : meta_363_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5497 = _T ? _GEN_4981 : meta_364_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5498 = _T ? _GEN_4982 : meta_365_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5499 = _T ? _GEN_4983 : meta_366_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5500 = _T ? _GEN_4984 : meta_367_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5501 = _T ? _GEN_4985 : meta_368_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5502 = _T ? _GEN_4986 : meta_369_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5503 = _T ? _GEN_4987 : meta_370_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5504 = _T ? _GEN_4988 : meta_371_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5505 = _T ? _GEN_4989 : meta_372_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5506 = _T ? _GEN_4990 : meta_373_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5507 = _T ? _GEN_4991 : meta_374_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5508 = _T ? _GEN_4992 : meta_375_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5509 = _T ? _GEN_4993 : meta_376_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5510 = _T ? _GEN_4994 : meta_377_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5511 = _T ? _GEN_4995 : meta_378_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5512 = _T ? _GEN_4996 : meta_379_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5513 = _T ? _GEN_4997 : meta_380_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5514 = _T ? _GEN_4998 : meta_381_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5515 = _T ? _GEN_4999 : meta_382_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5516 = _T ? _GEN_5000 : meta_383_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5517 = _T ? _GEN_5001 : meta_384_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5518 = _T ? _GEN_5002 : meta_385_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5519 = _T ? _GEN_5003 : meta_386_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5520 = _T ? _GEN_5004 : meta_387_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5521 = _T ? _GEN_5005 : meta_388_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5522 = _T ? _GEN_5006 : meta_389_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5523 = _T ? _GEN_5007 : meta_390_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5524 = _T ? _GEN_5008 : meta_391_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5525 = _T ? _GEN_5009 : meta_392_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5526 = _T ? _GEN_5010 : meta_393_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5527 = _T ? _GEN_5011 : meta_394_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5528 = _T ? _GEN_5012 : meta_395_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5529 = _T ? _GEN_5013 : meta_396_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5530 = _T ? _GEN_5014 : meta_397_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5531 = _T ? _GEN_5015 : meta_398_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5532 = _T ? _GEN_5016 : meta_399_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5533 = _T ? _GEN_5017 : meta_400_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5534 = _T ? _GEN_5018 : meta_401_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5535 = _T ? _GEN_5019 : meta_402_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5536 = _T ? _GEN_5020 : meta_403_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5537 = _T ? _GEN_5021 : meta_404_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5538 = _T ? _GEN_5022 : meta_405_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5539 = _T ? _GEN_5023 : meta_406_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5540 = _T ? _GEN_5024 : meta_407_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5541 = _T ? _GEN_5025 : meta_408_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5542 = _T ? _GEN_5026 : meta_409_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5543 = _T ? _GEN_5027 : meta_410_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5544 = _T ? _GEN_5028 : meta_411_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5545 = _T ? _GEN_5029 : meta_412_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5546 = _T ? _GEN_5030 : meta_413_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5547 = _T ? _GEN_5031 : meta_414_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5548 = _T ? _GEN_5032 : meta_415_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5549 = _T ? _GEN_5033 : meta_416_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5550 = _T ? _GEN_5034 : meta_417_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5551 = _T ? _GEN_5035 : meta_418_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5552 = _T ? _GEN_5036 : meta_419_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5553 = _T ? _GEN_5037 : meta_420_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5554 = _T ? _GEN_5038 : meta_421_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5555 = _T ? _GEN_5039 : meta_422_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5556 = _T ? _GEN_5040 : meta_423_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5557 = _T ? _GEN_5041 : meta_424_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5558 = _T ? _GEN_5042 : meta_425_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5559 = _T ? _GEN_5043 : meta_426_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5560 = _T ? _GEN_5044 : meta_427_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5561 = _T ? _GEN_5045 : meta_428_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5562 = _T ? _GEN_5046 : meta_429_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5563 = _T ? _GEN_5047 : meta_430_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5564 = _T ? _GEN_5048 : meta_431_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5565 = _T ? _GEN_5049 : meta_432_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5566 = _T ? _GEN_5050 : meta_433_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5567 = _T ? _GEN_5051 : meta_434_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5568 = _T ? _GEN_5052 : meta_435_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5569 = _T ? _GEN_5053 : meta_436_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5570 = _T ? _GEN_5054 : meta_437_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5571 = _T ? _GEN_5055 : meta_438_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5572 = _T ? _GEN_5056 : meta_439_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5573 = _T ? _GEN_5057 : meta_440_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5574 = _T ? _GEN_5058 : meta_441_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5575 = _T ? _GEN_5059 : meta_442_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5576 = _T ? _GEN_5060 : meta_443_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5577 = _T ? _GEN_5061 : meta_444_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5578 = _T ? _GEN_5062 : meta_445_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5579 = _T ? _GEN_5063 : meta_446_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5580 = _T ? _GEN_5064 : meta_447_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5581 = _T ? _GEN_5065 : meta_448_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5582 = _T ? _GEN_5066 : meta_449_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5583 = _T ? _GEN_5067 : meta_450_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5584 = _T ? _GEN_5068 : meta_451_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5585 = _T ? _GEN_5069 : meta_452_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5586 = _T ? _GEN_5070 : meta_453_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5587 = _T ? _GEN_5071 : meta_454_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5588 = _T ? _GEN_5072 : meta_455_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5589 = _T ? _GEN_5073 : meta_456_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5590 = _T ? _GEN_5074 : meta_457_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5591 = _T ? _GEN_5075 : meta_458_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5592 = _T ? _GEN_5076 : meta_459_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5593 = _T ? _GEN_5077 : meta_460_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5594 = _T ? _GEN_5078 : meta_461_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5595 = _T ? _GEN_5079 : meta_462_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5596 = _T ? _GEN_5080 : meta_463_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5597 = _T ? _GEN_5081 : meta_464_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5598 = _T ? _GEN_5082 : meta_465_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5599 = _T ? _GEN_5083 : meta_466_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5600 = _T ? _GEN_5084 : meta_467_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5601 = _T ? _GEN_5085 : meta_468_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5602 = _T ? _GEN_5086 : meta_469_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5603 = _T ? _GEN_5087 : meta_470_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5604 = _T ? _GEN_5088 : meta_471_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5605 = _T ? _GEN_5089 : meta_472_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5606 = _T ? _GEN_5090 : meta_473_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5607 = _T ? _GEN_5091 : meta_474_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5608 = _T ? _GEN_5092 : meta_475_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5609 = _T ? _GEN_5093 : meta_476_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5610 = _T ? _GEN_5094 : meta_477_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5611 = _T ? _GEN_5095 : meta_478_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5612 = _T ? _GEN_5096 : meta_479_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5613 = _T ? _GEN_5097 : meta_480_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5614 = _T ? _GEN_5098 : meta_481_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5615 = _T ? _GEN_5099 : meta_482_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5616 = _T ? _GEN_5100 : meta_483_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5617 = _T ? _GEN_5101 : meta_484_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5618 = _T ? _GEN_5102 : meta_485_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5619 = _T ? _GEN_5103 : meta_486_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5620 = _T ? _GEN_5104 : meta_487_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5621 = _T ? _GEN_5105 : meta_488_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5622 = _T ? _GEN_5106 : meta_489_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5623 = _T ? _GEN_5107 : meta_490_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5624 = _T ? _GEN_5108 : meta_491_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5625 = _T ? _GEN_5109 : meta_492_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5626 = _T ? _GEN_5110 : meta_493_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5627 = _T ? _GEN_5111 : meta_494_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5628 = _T ? _GEN_5112 : meta_495_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5629 = _T ? _GEN_5113 : meta_496_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5630 = _T ? _GEN_5114 : meta_497_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5631 = _T ? _GEN_5115 : meta_498_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5632 = _T ? _GEN_5116 : meta_499_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5633 = _T ? _GEN_5117 : meta_500_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5634 = _T ? _GEN_5118 : meta_501_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5635 = _T ? _GEN_5119 : meta_502_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5636 = _T ? _GEN_5120 : meta_503_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5637 = _T ? _GEN_5121 : meta_504_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5638 = _T ? _GEN_5122 : meta_505_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5639 = _T ? _GEN_5123 : meta_506_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5640 = _T ? _GEN_5124 : meta_507_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5641 = _T ? _GEN_5125 : meta_508_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5642 = _T ? _GEN_5126 : meta_509_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5643 = _T ? _GEN_5127 : meta_510_lru; // @[ICache.scala 188:42 34:21]
  wire  _GEN_5644 = _T ? _GEN_5128 : meta_511_lru; // @[ICache.scala 188:42 34:21]
  wire [2:0] _GEN_5645 = _T ? _GEN_5129 : state; // @[ICache.scala 188:42 48:81]
  wire [63:0] _GEN_5646 = _T ? _GEN_5130 : {{32'd0}, saved_1_inst}; // @[ICache.scala 188:42 91:22]
  wire  _GEN_5647 = _T ? _GEN_5131 : saved_0_valid; // @[ICache.scala 188:42 91:22]
  wire  _GEN_5648 = _T ? _GEN_5132 : saved_1_valid; // @[ICache.scala 188:42 91:22]
  wire [2:0] _GEN_5649 = ~cache_hit ? 3'h3 : _GEN_5645; // @[ICache.scala 175:32 176:19]
  wire [31:0] _GEN_5650 = ~cache_hit ? _ar_addr_T_1 : ar_addr; // @[ICache.scala 175:32 177:19 141:24]
  wire [7:0] _GEN_5651 = ~cache_hit ? 8'hf : ar_len; // @[ICache.scala 175:32 178:19 141:24]
  wire [2:0] _GEN_5652 = ~cache_hit ? 3'h2 : ar_size; // @[ICache.scala 175:32 179:19 141:24]
  wire  _GEN_5653 = ~cache_hit | arvalid; // @[ICache.scala 175:32 180:19 142:24]
  wire [5:0] _GEN_5654 = ~cache_hit ? va_line_addr : replace_line_addr; // @[ICache.scala 175:32 182:60 58:38]
  wire [7:0] _GEN_5655 = ~cache_hit ? _GEN_3589 : data_wen_0; // @[ICache.scala 175:32 66:30]
  wire [7:0] _GEN_5656 = ~cache_hit ? _GEN_3590 : data_wen_1; // @[ICache.scala 175:32 66:30]
  wire  _GEN_5657 = ~cache_hit ? _GEN_3591 : tag_wen_0; // @[ICache.scala 175:32 67:30]
  wire  _GEN_5658 = ~cache_hit ? _GEN_3592 : tag_wen_1; // @[ICache.scala 175:32 67:30]
  wire [19:0] _GEN_5659 = ~cache_hit ? inst_tag : {{3'd0}, tag_ram_wdata}; // @[ICache.scala 175:32 185:60 68:30]
  wire  _GEN_5660 = ~cache_hit ? _GEN_3593 : _GEN_2053; // @[ICache.scala 175:32]
  wire  _GEN_5661 = ~cache_hit ? _GEN_3594 : _GEN_2565; // @[ICache.scala 175:32]
  wire  _GEN_5662 = ~cache_hit ? _GEN_3595 : _GEN_2054; // @[ICache.scala 175:32]
  wire  _GEN_5663 = ~cache_hit ? _GEN_3596 : _GEN_2566; // @[ICache.scala 175:32]
  wire  _GEN_5664 = ~cache_hit ? _GEN_3597 : _GEN_2055; // @[ICache.scala 175:32]
  wire  _GEN_5665 = ~cache_hit ? _GEN_3598 : _GEN_2567; // @[ICache.scala 175:32]
  wire  _GEN_5666 = ~cache_hit ? _GEN_3599 : _GEN_2056; // @[ICache.scala 175:32]
  wire  _GEN_5667 = ~cache_hit ? _GEN_3600 : _GEN_2568; // @[ICache.scala 175:32]
  wire  _GEN_5668 = ~cache_hit ? _GEN_3601 : _GEN_2057; // @[ICache.scala 175:32]
  wire  _GEN_5669 = ~cache_hit ? _GEN_3602 : _GEN_2569; // @[ICache.scala 175:32]
  wire  _GEN_5670 = ~cache_hit ? _GEN_3603 : _GEN_2058; // @[ICache.scala 175:32]
  wire  _GEN_5671 = ~cache_hit ? _GEN_3604 : _GEN_2570; // @[ICache.scala 175:32]
  wire  _GEN_5672 = ~cache_hit ? _GEN_3605 : _GEN_2059; // @[ICache.scala 175:32]
  wire  _GEN_5673 = ~cache_hit ? _GEN_3606 : _GEN_2571; // @[ICache.scala 175:32]
  wire  _GEN_5674 = ~cache_hit ? _GEN_3607 : _GEN_2060; // @[ICache.scala 175:32]
  wire  _GEN_5675 = ~cache_hit ? _GEN_3608 : _GEN_2572; // @[ICache.scala 175:32]
  wire  _GEN_5676 = ~cache_hit ? _GEN_3609 : _GEN_2061; // @[ICache.scala 175:32]
  wire  _GEN_5677 = ~cache_hit ? _GEN_3610 : _GEN_2573; // @[ICache.scala 175:32]
  wire  _GEN_5678 = ~cache_hit ? _GEN_3611 : _GEN_2062; // @[ICache.scala 175:32]
  wire  _GEN_5679 = ~cache_hit ? _GEN_3612 : _GEN_2574; // @[ICache.scala 175:32]
  wire  _GEN_5680 = ~cache_hit ? _GEN_3613 : _GEN_2063; // @[ICache.scala 175:32]
  wire  _GEN_5681 = ~cache_hit ? _GEN_3614 : _GEN_2575; // @[ICache.scala 175:32]
  wire  _GEN_5682 = ~cache_hit ? _GEN_3615 : _GEN_2064; // @[ICache.scala 175:32]
  wire  _GEN_5683 = ~cache_hit ? _GEN_3616 : _GEN_2576; // @[ICache.scala 175:32]
  wire  _GEN_5684 = ~cache_hit ? _GEN_3617 : _GEN_2065; // @[ICache.scala 175:32]
  wire  _GEN_5685 = ~cache_hit ? _GEN_3618 : _GEN_2577; // @[ICache.scala 175:32]
  wire  _GEN_5686 = ~cache_hit ? _GEN_3619 : _GEN_2066; // @[ICache.scala 175:32]
  wire  _GEN_5687 = ~cache_hit ? _GEN_3620 : _GEN_2578; // @[ICache.scala 175:32]
  wire  _GEN_5688 = ~cache_hit ? _GEN_3621 : _GEN_2067; // @[ICache.scala 175:32]
  wire  _GEN_5689 = ~cache_hit ? _GEN_3622 : _GEN_2579; // @[ICache.scala 175:32]
  wire  _GEN_5690 = ~cache_hit ? _GEN_3623 : _GEN_2068; // @[ICache.scala 175:32]
  wire  _GEN_5691 = ~cache_hit ? _GEN_3624 : _GEN_2580; // @[ICache.scala 175:32]
  wire  _GEN_5692 = ~cache_hit ? _GEN_3625 : _GEN_2069; // @[ICache.scala 175:32]
  wire  _GEN_5693 = ~cache_hit ? _GEN_3626 : _GEN_2581; // @[ICache.scala 175:32]
  wire  _GEN_5694 = ~cache_hit ? _GEN_3627 : _GEN_2070; // @[ICache.scala 175:32]
  wire  _GEN_5695 = ~cache_hit ? _GEN_3628 : _GEN_2582; // @[ICache.scala 175:32]
  wire  _GEN_5696 = ~cache_hit ? _GEN_3629 : _GEN_2071; // @[ICache.scala 175:32]
  wire  _GEN_5697 = ~cache_hit ? _GEN_3630 : _GEN_2583; // @[ICache.scala 175:32]
  wire  _GEN_5698 = ~cache_hit ? _GEN_3631 : _GEN_2072; // @[ICache.scala 175:32]
  wire  _GEN_5699 = ~cache_hit ? _GEN_3632 : _GEN_2584; // @[ICache.scala 175:32]
  wire  _GEN_5700 = ~cache_hit ? _GEN_3633 : _GEN_2073; // @[ICache.scala 175:32]
  wire  _GEN_5701 = ~cache_hit ? _GEN_3634 : _GEN_2585; // @[ICache.scala 175:32]
  wire  _GEN_5702 = ~cache_hit ? _GEN_3635 : _GEN_2074; // @[ICache.scala 175:32]
  wire  _GEN_5703 = ~cache_hit ? _GEN_3636 : _GEN_2586; // @[ICache.scala 175:32]
  wire  _GEN_5704 = ~cache_hit ? _GEN_3637 : _GEN_2075; // @[ICache.scala 175:32]
  wire  _GEN_5705 = ~cache_hit ? _GEN_3638 : _GEN_2587; // @[ICache.scala 175:32]
  wire  _GEN_5706 = ~cache_hit ? _GEN_3639 : _GEN_2076; // @[ICache.scala 175:32]
  wire  _GEN_5707 = ~cache_hit ? _GEN_3640 : _GEN_2588; // @[ICache.scala 175:32]
  wire  _GEN_5708 = ~cache_hit ? _GEN_3641 : _GEN_2077; // @[ICache.scala 175:32]
  wire  _GEN_5709 = ~cache_hit ? _GEN_3642 : _GEN_2589; // @[ICache.scala 175:32]
  wire  _GEN_5710 = ~cache_hit ? _GEN_3643 : _GEN_2078; // @[ICache.scala 175:32]
  wire  _GEN_5711 = ~cache_hit ? _GEN_3644 : _GEN_2590; // @[ICache.scala 175:32]
  wire  _GEN_5712 = ~cache_hit ? _GEN_3645 : _GEN_2079; // @[ICache.scala 175:32]
  wire  _GEN_5713 = ~cache_hit ? _GEN_3646 : _GEN_2591; // @[ICache.scala 175:32]
  wire  _GEN_5714 = ~cache_hit ? _GEN_3647 : _GEN_2080; // @[ICache.scala 175:32]
  wire  _GEN_5715 = ~cache_hit ? _GEN_3648 : _GEN_2592; // @[ICache.scala 175:32]
  wire  _GEN_5716 = ~cache_hit ? _GEN_3649 : _GEN_2081; // @[ICache.scala 175:32]
  wire  _GEN_5717 = ~cache_hit ? _GEN_3650 : _GEN_2593; // @[ICache.scala 175:32]
  wire  _GEN_5718 = ~cache_hit ? _GEN_3651 : _GEN_2082; // @[ICache.scala 175:32]
  wire  _GEN_5719 = ~cache_hit ? _GEN_3652 : _GEN_2594; // @[ICache.scala 175:32]
  wire  _GEN_5720 = ~cache_hit ? _GEN_3653 : _GEN_2083; // @[ICache.scala 175:32]
  wire  _GEN_5721 = ~cache_hit ? _GEN_3654 : _GEN_2595; // @[ICache.scala 175:32]
  wire  _GEN_5722 = ~cache_hit ? _GEN_3655 : _GEN_2084; // @[ICache.scala 175:32]
  wire  _GEN_5723 = ~cache_hit ? _GEN_3656 : _GEN_2596; // @[ICache.scala 175:32]
  wire  _GEN_5724 = ~cache_hit ? _GEN_3657 : _GEN_2085; // @[ICache.scala 175:32]
  wire  _GEN_5725 = ~cache_hit ? _GEN_3658 : _GEN_2597; // @[ICache.scala 175:32]
  wire  _GEN_5726 = ~cache_hit ? _GEN_3659 : _GEN_2086; // @[ICache.scala 175:32]
  wire  _GEN_5727 = ~cache_hit ? _GEN_3660 : _GEN_2598; // @[ICache.scala 175:32]
  wire  _GEN_5728 = ~cache_hit ? _GEN_3661 : _GEN_2087; // @[ICache.scala 175:32]
  wire  _GEN_5729 = ~cache_hit ? _GEN_3662 : _GEN_2599; // @[ICache.scala 175:32]
  wire  _GEN_5730 = ~cache_hit ? _GEN_3663 : _GEN_2088; // @[ICache.scala 175:32]
  wire  _GEN_5731 = ~cache_hit ? _GEN_3664 : _GEN_2600; // @[ICache.scala 175:32]
  wire  _GEN_5732 = ~cache_hit ? _GEN_3665 : _GEN_2089; // @[ICache.scala 175:32]
  wire  _GEN_5733 = ~cache_hit ? _GEN_3666 : _GEN_2601; // @[ICache.scala 175:32]
  wire  _GEN_5734 = ~cache_hit ? _GEN_3667 : _GEN_2090; // @[ICache.scala 175:32]
  wire  _GEN_5735 = ~cache_hit ? _GEN_3668 : _GEN_2602; // @[ICache.scala 175:32]
  wire  _GEN_5736 = ~cache_hit ? _GEN_3669 : _GEN_2091; // @[ICache.scala 175:32]
  wire  _GEN_5737 = ~cache_hit ? _GEN_3670 : _GEN_2603; // @[ICache.scala 175:32]
  wire  _GEN_5738 = ~cache_hit ? _GEN_3671 : _GEN_2092; // @[ICache.scala 175:32]
  wire  _GEN_5739 = ~cache_hit ? _GEN_3672 : _GEN_2604; // @[ICache.scala 175:32]
  wire  _GEN_5740 = ~cache_hit ? _GEN_3673 : _GEN_2093; // @[ICache.scala 175:32]
  wire  _GEN_5741 = ~cache_hit ? _GEN_3674 : _GEN_2605; // @[ICache.scala 175:32]
  wire  _GEN_5742 = ~cache_hit ? _GEN_3675 : _GEN_2094; // @[ICache.scala 175:32]
  wire  _GEN_5743 = ~cache_hit ? _GEN_3676 : _GEN_2606; // @[ICache.scala 175:32]
  wire  _GEN_5744 = ~cache_hit ? _GEN_3677 : _GEN_2095; // @[ICache.scala 175:32]
  wire  _GEN_5745 = ~cache_hit ? _GEN_3678 : _GEN_2607; // @[ICache.scala 175:32]
  wire  _GEN_5746 = ~cache_hit ? _GEN_3679 : _GEN_2096; // @[ICache.scala 175:32]
  wire  _GEN_5747 = ~cache_hit ? _GEN_3680 : _GEN_2608; // @[ICache.scala 175:32]
  wire  _GEN_5748 = ~cache_hit ? _GEN_3681 : _GEN_2097; // @[ICache.scala 175:32]
  wire  _GEN_5749 = ~cache_hit ? _GEN_3682 : _GEN_2609; // @[ICache.scala 175:32]
  wire  _GEN_5750 = ~cache_hit ? _GEN_3683 : _GEN_2098; // @[ICache.scala 175:32]
  wire  _GEN_5751 = ~cache_hit ? _GEN_3684 : _GEN_2610; // @[ICache.scala 175:32]
  wire  _GEN_5752 = ~cache_hit ? _GEN_3685 : _GEN_2099; // @[ICache.scala 175:32]
  wire  _GEN_5753 = ~cache_hit ? _GEN_3686 : _GEN_2611; // @[ICache.scala 175:32]
  wire  _GEN_5754 = ~cache_hit ? _GEN_3687 : _GEN_2100; // @[ICache.scala 175:32]
  wire  _GEN_5755 = ~cache_hit ? _GEN_3688 : _GEN_2612; // @[ICache.scala 175:32]
  wire  _GEN_5756 = ~cache_hit ? _GEN_3689 : _GEN_2101; // @[ICache.scala 175:32]
  wire  _GEN_5757 = ~cache_hit ? _GEN_3690 : _GEN_2613; // @[ICache.scala 175:32]
  wire  _GEN_5758 = ~cache_hit ? _GEN_3691 : _GEN_2102; // @[ICache.scala 175:32]
  wire  _GEN_5759 = ~cache_hit ? _GEN_3692 : _GEN_2614; // @[ICache.scala 175:32]
  wire  _GEN_5760 = ~cache_hit ? _GEN_3693 : _GEN_2103; // @[ICache.scala 175:32]
  wire  _GEN_5761 = ~cache_hit ? _GEN_3694 : _GEN_2615; // @[ICache.scala 175:32]
  wire  _GEN_5762 = ~cache_hit ? _GEN_3695 : _GEN_2104; // @[ICache.scala 175:32]
  wire  _GEN_5763 = ~cache_hit ? _GEN_3696 : _GEN_2616; // @[ICache.scala 175:32]
  wire  _GEN_5764 = ~cache_hit ? _GEN_3697 : _GEN_2105; // @[ICache.scala 175:32]
  wire  _GEN_5765 = ~cache_hit ? _GEN_3698 : _GEN_2617; // @[ICache.scala 175:32]
  wire  _GEN_5766 = ~cache_hit ? _GEN_3699 : _GEN_2106; // @[ICache.scala 175:32]
  wire  _GEN_5767 = ~cache_hit ? _GEN_3700 : _GEN_2618; // @[ICache.scala 175:32]
  wire  _GEN_5768 = ~cache_hit ? _GEN_3701 : _GEN_2107; // @[ICache.scala 175:32]
  wire  _GEN_5769 = ~cache_hit ? _GEN_3702 : _GEN_2619; // @[ICache.scala 175:32]
  wire  _GEN_5770 = ~cache_hit ? _GEN_3703 : _GEN_2108; // @[ICache.scala 175:32]
  wire  _GEN_5771 = ~cache_hit ? _GEN_3704 : _GEN_2620; // @[ICache.scala 175:32]
  wire  _GEN_5772 = ~cache_hit ? _GEN_3705 : _GEN_2109; // @[ICache.scala 175:32]
  wire  _GEN_5773 = ~cache_hit ? _GEN_3706 : _GEN_2621; // @[ICache.scala 175:32]
  wire  _GEN_5774 = ~cache_hit ? _GEN_3707 : _GEN_2110; // @[ICache.scala 175:32]
  wire  _GEN_5775 = ~cache_hit ? _GEN_3708 : _GEN_2622; // @[ICache.scala 175:32]
  wire  _GEN_5776 = ~cache_hit ? _GEN_3709 : _GEN_2111; // @[ICache.scala 175:32]
  wire  _GEN_5777 = ~cache_hit ? _GEN_3710 : _GEN_2623; // @[ICache.scala 175:32]
  wire  _GEN_5778 = ~cache_hit ? _GEN_3711 : _GEN_2112; // @[ICache.scala 175:32]
  wire  _GEN_5779 = ~cache_hit ? _GEN_3712 : _GEN_2624; // @[ICache.scala 175:32]
  wire  _GEN_5780 = ~cache_hit ? _GEN_3713 : _GEN_2113; // @[ICache.scala 175:32]
  wire  _GEN_5781 = ~cache_hit ? _GEN_3714 : _GEN_2625; // @[ICache.scala 175:32]
  wire  _GEN_5782 = ~cache_hit ? _GEN_3715 : _GEN_2114; // @[ICache.scala 175:32]
  wire  _GEN_5783 = ~cache_hit ? _GEN_3716 : _GEN_2626; // @[ICache.scala 175:32]
  wire  _GEN_5784 = ~cache_hit ? _GEN_3717 : _GEN_2115; // @[ICache.scala 175:32]
  wire  _GEN_5785 = ~cache_hit ? _GEN_3718 : _GEN_2627; // @[ICache.scala 175:32]
  wire  _GEN_5786 = ~cache_hit ? _GEN_3719 : _GEN_2116; // @[ICache.scala 175:32]
  wire  _GEN_5787 = ~cache_hit ? _GEN_3720 : _GEN_2628; // @[ICache.scala 175:32]
  wire  _GEN_5788 = ~cache_hit ? _GEN_3721 : _GEN_2117; // @[ICache.scala 175:32]
  wire  _GEN_5789 = ~cache_hit ? _GEN_3722 : _GEN_2629; // @[ICache.scala 175:32]
  wire  _GEN_5790 = ~cache_hit ? _GEN_3723 : _GEN_2118; // @[ICache.scala 175:32]
  wire  _GEN_5791 = ~cache_hit ? _GEN_3724 : _GEN_2630; // @[ICache.scala 175:32]
  wire  _GEN_5792 = ~cache_hit ? _GEN_3725 : _GEN_2119; // @[ICache.scala 175:32]
  wire  _GEN_5793 = ~cache_hit ? _GEN_3726 : _GEN_2631; // @[ICache.scala 175:32]
  wire  _GEN_5794 = ~cache_hit ? _GEN_3727 : _GEN_2120; // @[ICache.scala 175:32]
  wire  _GEN_5795 = ~cache_hit ? _GEN_3728 : _GEN_2632; // @[ICache.scala 175:32]
  wire  _GEN_5796 = ~cache_hit ? _GEN_3729 : _GEN_2121; // @[ICache.scala 175:32]
  wire  _GEN_5797 = ~cache_hit ? _GEN_3730 : _GEN_2633; // @[ICache.scala 175:32]
  wire  _GEN_5798 = ~cache_hit ? _GEN_3731 : _GEN_2122; // @[ICache.scala 175:32]
  wire  _GEN_5799 = ~cache_hit ? _GEN_3732 : _GEN_2634; // @[ICache.scala 175:32]
  wire  _GEN_5800 = ~cache_hit ? _GEN_3733 : _GEN_2123; // @[ICache.scala 175:32]
  wire  _GEN_5801 = ~cache_hit ? _GEN_3734 : _GEN_2635; // @[ICache.scala 175:32]
  wire  _GEN_5802 = ~cache_hit ? _GEN_3735 : _GEN_2124; // @[ICache.scala 175:32]
  wire  _GEN_5803 = ~cache_hit ? _GEN_3736 : _GEN_2636; // @[ICache.scala 175:32]
  wire  _GEN_5804 = ~cache_hit ? _GEN_3737 : _GEN_2125; // @[ICache.scala 175:32]
  wire  _GEN_5805 = ~cache_hit ? _GEN_3738 : _GEN_2637; // @[ICache.scala 175:32]
  wire  _GEN_5806 = ~cache_hit ? _GEN_3739 : _GEN_2126; // @[ICache.scala 175:32]
  wire  _GEN_5807 = ~cache_hit ? _GEN_3740 : _GEN_2638; // @[ICache.scala 175:32]
  wire  _GEN_5808 = ~cache_hit ? _GEN_3741 : _GEN_2127; // @[ICache.scala 175:32]
  wire  _GEN_5809 = ~cache_hit ? _GEN_3742 : _GEN_2639; // @[ICache.scala 175:32]
  wire  _GEN_5810 = ~cache_hit ? _GEN_3743 : _GEN_2128; // @[ICache.scala 175:32]
  wire  _GEN_5811 = ~cache_hit ? _GEN_3744 : _GEN_2640; // @[ICache.scala 175:32]
  wire  _GEN_5812 = ~cache_hit ? _GEN_3745 : _GEN_2129; // @[ICache.scala 175:32]
  wire  _GEN_5813 = ~cache_hit ? _GEN_3746 : _GEN_2641; // @[ICache.scala 175:32]
  wire  _GEN_5814 = ~cache_hit ? _GEN_3747 : _GEN_2130; // @[ICache.scala 175:32]
  wire  _GEN_5815 = ~cache_hit ? _GEN_3748 : _GEN_2642; // @[ICache.scala 175:32]
  wire  _GEN_5816 = ~cache_hit ? _GEN_3749 : _GEN_2131; // @[ICache.scala 175:32]
  wire  _GEN_5817 = ~cache_hit ? _GEN_3750 : _GEN_2643; // @[ICache.scala 175:32]
  wire  _GEN_5818 = ~cache_hit ? _GEN_3751 : _GEN_2132; // @[ICache.scala 175:32]
  wire  _GEN_5819 = ~cache_hit ? _GEN_3752 : _GEN_2644; // @[ICache.scala 175:32]
  wire  _GEN_5820 = ~cache_hit ? _GEN_3753 : _GEN_2133; // @[ICache.scala 175:32]
  wire  _GEN_5821 = ~cache_hit ? _GEN_3754 : _GEN_2645; // @[ICache.scala 175:32]
  wire  _GEN_5822 = ~cache_hit ? _GEN_3755 : _GEN_2134; // @[ICache.scala 175:32]
  wire  _GEN_5823 = ~cache_hit ? _GEN_3756 : _GEN_2646; // @[ICache.scala 175:32]
  wire  _GEN_5824 = ~cache_hit ? _GEN_3757 : _GEN_2135; // @[ICache.scala 175:32]
  wire  _GEN_5825 = ~cache_hit ? _GEN_3758 : _GEN_2647; // @[ICache.scala 175:32]
  wire  _GEN_5826 = ~cache_hit ? _GEN_3759 : _GEN_2136; // @[ICache.scala 175:32]
  wire  _GEN_5827 = ~cache_hit ? _GEN_3760 : _GEN_2648; // @[ICache.scala 175:32]
  wire  _GEN_5828 = ~cache_hit ? _GEN_3761 : _GEN_2137; // @[ICache.scala 175:32]
  wire  _GEN_5829 = ~cache_hit ? _GEN_3762 : _GEN_2649; // @[ICache.scala 175:32]
  wire  _GEN_5830 = ~cache_hit ? _GEN_3763 : _GEN_2138; // @[ICache.scala 175:32]
  wire  _GEN_5831 = ~cache_hit ? _GEN_3764 : _GEN_2650; // @[ICache.scala 175:32]
  wire  _GEN_5832 = ~cache_hit ? _GEN_3765 : _GEN_2139; // @[ICache.scala 175:32]
  wire  _GEN_5833 = ~cache_hit ? _GEN_3766 : _GEN_2651; // @[ICache.scala 175:32]
  wire  _GEN_5834 = ~cache_hit ? _GEN_3767 : _GEN_2140; // @[ICache.scala 175:32]
  wire  _GEN_5835 = ~cache_hit ? _GEN_3768 : _GEN_2652; // @[ICache.scala 175:32]
  wire  _GEN_5836 = ~cache_hit ? _GEN_3769 : _GEN_2141; // @[ICache.scala 175:32]
  wire  _GEN_5837 = ~cache_hit ? _GEN_3770 : _GEN_2653; // @[ICache.scala 175:32]
  wire  _GEN_5838 = ~cache_hit ? _GEN_3771 : _GEN_2142; // @[ICache.scala 175:32]
  wire  _GEN_5839 = ~cache_hit ? _GEN_3772 : _GEN_2654; // @[ICache.scala 175:32]
  wire  _GEN_5840 = ~cache_hit ? _GEN_3773 : _GEN_2143; // @[ICache.scala 175:32]
  wire  _GEN_5841 = ~cache_hit ? _GEN_3774 : _GEN_2655; // @[ICache.scala 175:32]
  wire  _GEN_5842 = ~cache_hit ? _GEN_3775 : _GEN_2144; // @[ICache.scala 175:32]
  wire  _GEN_5843 = ~cache_hit ? _GEN_3776 : _GEN_2656; // @[ICache.scala 175:32]
  wire  _GEN_5844 = ~cache_hit ? _GEN_3777 : _GEN_2145; // @[ICache.scala 175:32]
  wire  _GEN_5845 = ~cache_hit ? _GEN_3778 : _GEN_2657; // @[ICache.scala 175:32]
  wire  _GEN_5846 = ~cache_hit ? _GEN_3779 : _GEN_2146; // @[ICache.scala 175:32]
  wire  _GEN_5847 = ~cache_hit ? _GEN_3780 : _GEN_2658; // @[ICache.scala 175:32]
  wire  _GEN_5848 = ~cache_hit ? _GEN_3781 : _GEN_2147; // @[ICache.scala 175:32]
  wire  _GEN_5849 = ~cache_hit ? _GEN_3782 : _GEN_2659; // @[ICache.scala 175:32]
  wire  _GEN_5850 = ~cache_hit ? _GEN_3783 : _GEN_2148; // @[ICache.scala 175:32]
  wire  _GEN_5851 = ~cache_hit ? _GEN_3784 : _GEN_2660; // @[ICache.scala 175:32]
  wire  _GEN_5852 = ~cache_hit ? _GEN_3785 : _GEN_2149; // @[ICache.scala 175:32]
  wire  _GEN_5853 = ~cache_hit ? _GEN_3786 : _GEN_2661; // @[ICache.scala 175:32]
  wire  _GEN_5854 = ~cache_hit ? _GEN_3787 : _GEN_2150; // @[ICache.scala 175:32]
  wire  _GEN_5855 = ~cache_hit ? _GEN_3788 : _GEN_2662; // @[ICache.scala 175:32]
  wire  _GEN_5856 = ~cache_hit ? _GEN_3789 : _GEN_2151; // @[ICache.scala 175:32]
  wire  _GEN_5857 = ~cache_hit ? _GEN_3790 : _GEN_2663; // @[ICache.scala 175:32]
  wire  _GEN_5858 = ~cache_hit ? _GEN_3791 : _GEN_2152; // @[ICache.scala 175:32]
  wire  _GEN_5859 = ~cache_hit ? _GEN_3792 : _GEN_2664; // @[ICache.scala 175:32]
  wire  _GEN_5860 = ~cache_hit ? _GEN_3793 : _GEN_2153; // @[ICache.scala 175:32]
  wire  _GEN_5861 = ~cache_hit ? _GEN_3794 : _GEN_2665; // @[ICache.scala 175:32]
  wire  _GEN_5862 = ~cache_hit ? _GEN_3795 : _GEN_2154; // @[ICache.scala 175:32]
  wire  _GEN_5863 = ~cache_hit ? _GEN_3796 : _GEN_2666; // @[ICache.scala 175:32]
  wire  _GEN_5864 = ~cache_hit ? _GEN_3797 : _GEN_2155; // @[ICache.scala 175:32]
  wire  _GEN_5865 = ~cache_hit ? _GEN_3798 : _GEN_2667; // @[ICache.scala 175:32]
  wire  _GEN_5866 = ~cache_hit ? _GEN_3799 : _GEN_2156; // @[ICache.scala 175:32]
  wire  _GEN_5867 = ~cache_hit ? _GEN_3800 : _GEN_2668; // @[ICache.scala 175:32]
  wire  _GEN_5868 = ~cache_hit ? _GEN_3801 : _GEN_2157; // @[ICache.scala 175:32]
  wire  _GEN_5869 = ~cache_hit ? _GEN_3802 : _GEN_2669; // @[ICache.scala 175:32]
  wire  _GEN_5870 = ~cache_hit ? _GEN_3803 : _GEN_2158; // @[ICache.scala 175:32]
  wire  _GEN_5871 = ~cache_hit ? _GEN_3804 : _GEN_2670; // @[ICache.scala 175:32]
  wire  _GEN_5872 = ~cache_hit ? _GEN_3805 : _GEN_2159; // @[ICache.scala 175:32]
  wire  _GEN_5873 = ~cache_hit ? _GEN_3806 : _GEN_2671; // @[ICache.scala 175:32]
  wire  _GEN_5874 = ~cache_hit ? _GEN_3807 : _GEN_2160; // @[ICache.scala 175:32]
  wire  _GEN_5875 = ~cache_hit ? _GEN_3808 : _GEN_2672; // @[ICache.scala 175:32]
  wire  _GEN_5876 = ~cache_hit ? _GEN_3809 : _GEN_2161; // @[ICache.scala 175:32]
  wire  _GEN_5877 = ~cache_hit ? _GEN_3810 : _GEN_2673; // @[ICache.scala 175:32]
  wire  _GEN_5878 = ~cache_hit ? _GEN_3811 : _GEN_2162; // @[ICache.scala 175:32]
  wire  _GEN_5879 = ~cache_hit ? _GEN_3812 : _GEN_2674; // @[ICache.scala 175:32]
  wire  _GEN_5880 = ~cache_hit ? _GEN_3813 : _GEN_2163; // @[ICache.scala 175:32]
  wire  _GEN_5881 = ~cache_hit ? _GEN_3814 : _GEN_2675; // @[ICache.scala 175:32]
  wire  _GEN_5882 = ~cache_hit ? _GEN_3815 : _GEN_2164; // @[ICache.scala 175:32]
  wire  _GEN_5883 = ~cache_hit ? _GEN_3816 : _GEN_2676; // @[ICache.scala 175:32]
  wire  _GEN_5884 = ~cache_hit ? _GEN_3817 : _GEN_2165; // @[ICache.scala 175:32]
  wire  _GEN_5885 = ~cache_hit ? _GEN_3818 : _GEN_2677; // @[ICache.scala 175:32]
  wire  _GEN_5886 = ~cache_hit ? _GEN_3819 : _GEN_2166; // @[ICache.scala 175:32]
  wire  _GEN_5887 = ~cache_hit ? _GEN_3820 : _GEN_2678; // @[ICache.scala 175:32]
  wire  _GEN_5888 = ~cache_hit ? _GEN_3821 : _GEN_2167; // @[ICache.scala 175:32]
  wire  _GEN_5889 = ~cache_hit ? _GEN_3822 : _GEN_2679; // @[ICache.scala 175:32]
  wire  _GEN_5890 = ~cache_hit ? _GEN_3823 : _GEN_2168; // @[ICache.scala 175:32]
  wire  _GEN_5891 = ~cache_hit ? _GEN_3824 : _GEN_2680; // @[ICache.scala 175:32]
  wire  _GEN_5892 = ~cache_hit ? _GEN_3825 : _GEN_2169; // @[ICache.scala 175:32]
  wire  _GEN_5893 = ~cache_hit ? _GEN_3826 : _GEN_2681; // @[ICache.scala 175:32]
  wire  _GEN_5894 = ~cache_hit ? _GEN_3827 : _GEN_2170; // @[ICache.scala 175:32]
  wire  _GEN_5895 = ~cache_hit ? _GEN_3828 : _GEN_2682; // @[ICache.scala 175:32]
  wire  _GEN_5896 = ~cache_hit ? _GEN_3829 : _GEN_2171; // @[ICache.scala 175:32]
  wire  _GEN_5897 = ~cache_hit ? _GEN_3830 : _GEN_2683; // @[ICache.scala 175:32]
  wire  _GEN_5898 = ~cache_hit ? _GEN_3831 : _GEN_2172; // @[ICache.scala 175:32]
  wire  _GEN_5899 = ~cache_hit ? _GEN_3832 : _GEN_2684; // @[ICache.scala 175:32]
  wire  _GEN_5900 = ~cache_hit ? _GEN_3833 : _GEN_2173; // @[ICache.scala 175:32]
  wire  _GEN_5901 = ~cache_hit ? _GEN_3834 : _GEN_2685; // @[ICache.scala 175:32]
  wire  _GEN_5902 = ~cache_hit ? _GEN_3835 : _GEN_2174; // @[ICache.scala 175:32]
  wire  _GEN_5903 = ~cache_hit ? _GEN_3836 : _GEN_2686; // @[ICache.scala 175:32]
  wire  _GEN_5904 = ~cache_hit ? _GEN_3837 : _GEN_2175; // @[ICache.scala 175:32]
  wire  _GEN_5905 = ~cache_hit ? _GEN_3838 : _GEN_2687; // @[ICache.scala 175:32]
  wire  _GEN_5906 = ~cache_hit ? _GEN_3839 : _GEN_2176; // @[ICache.scala 175:32]
  wire  _GEN_5907 = ~cache_hit ? _GEN_3840 : _GEN_2688; // @[ICache.scala 175:32]
  wire  _GEN_5908 = ~cache_hit ? _GEN_3841 : _GEN_2177; // @[ICache.scala 175:32]
  wire  _GEN_5909 = ~cache_hit ? _GEN_3842 : _GEN_2689; // @[ICache.scala 175:32]
  wire  _GEN_5910 = ~cache_hit ? _GEN_3843 : _GEN_2178; // @[ICache.scala 175:32]
  wire  _GEN_5911 = ~cache_hit ? _GEN_3844 : _GEN_2690; // @[ICache.scala 175:32]
  wire  _GEN_5912 = ~cache_hit ? _GEN_3845 : _GEN_2179; // @[ICache.scala 175:32]
  wire  _GEN_5913 = ~cache_hit ? _GEN_3846 : _GEN_2691; // @[ICache.scala 175:32]
  wire  _GEN_5914 = ~cache_hit ? _GEN_3847 : _GEN_2180; // @[ICache.scala 175:32]
  wire  _GEN_5915 = ~cache_hit ? _GEN_3848 : _GEN_2692; // @[ICache.scala 175:32]
  wire  _GEN_5916 = ~cache_hit ? _GEN_3849 : _GEN_2181; // @[ICache.scala 175:32]
  wire  _GEN_5917 = ~cache_hit ? _GEN_3850 : _GEN_2693; // @[ICache.scala 175:32]
  wire  _GEN_5918 = ~cache_hit ? _GEN_3851 : _GEN_2182; // @[ICache.scala 175:32]
  wire  _GEN_5919 = ~cache_hit ? _GEN_3852 : _GEN_2694; // @[ICache.scala 175:32]
  wire  _GEN_5920 = ~cache_hit ? _GEN_3853 : _GEN_2183; // @[ICache.scala 175:32]
  wire  _GEN_5921 = ~cache_hit ? _GEN_3854 : _GEN_2695; // @[ICache.scala 175:32]
  wire  _GEN_5922 = ~cache_hit ? _GEN_3855 : _GEN_2184; // @[ICache.scala 175:32]
  wire  _GEN_5923 = ~cache_hit ? _GEN_3856 : _GEN_2696; // @[ICache.scala 175:32]
  wire  _GEN_5924 = ~cache_hit ? _GEN_3857 : _GEN_2185; // @[ICache.scala 175:32]
  wire  _GEN_5925 = ~cache_hit ? _GEN_3858 : _GEN_2697; // @[ICache.scala 175:32]
  wire  _GEN_5926 = ~cache_hit ? _GEN_3859 : _GEN_2186; // @[ICache.scala 175:32]
  wire  _GEN_5927 = ~cache_hit ? _GEN_3860 : _GEN_2698; // @[ICache.scala 175:32]
  wire  _GEN_5928 = ~cache_hit ? _GEN_3861 : _GEN_2187; // @[ICache.scala 175:32]
  wire  _GEN_5929 = ~cache_hit ? _GEN_3862 : _GEN_2699; // @[ICache.scala 175:32]
  wire  _GEN_5930 = ~cache_hit ? _GEN_3863 : _GEN_2188; // @[ICache.scala 175:32]
  wire  _GEN_5931 = ~cache_hit ? _GEN_3864 : _GEN_2700; // @[ICache.scala 175:32]
  wire  _GEN_5932 = ~cache_hit ? _GEN_3865 : _GEN_2189; // @[ICache.scala 175:32]
  wire  _GEN_5933 = ~cache_hit ? _GEN_3866 : _GEN_2701; // @[ICache.scala 175:32]
  wire  _GEN_5934 = ~cache_hit ? _GEN_3867 : _GEN_2190; // @[ICache.scala 175:32]
  wire  _GEN_5935 = ~cache_hit ? _GEN_3868 : _GEN_2702; // @[ICache.scala 175:32]
  wire  _GEN_5936 = ~cache_hit ? _GEN_3869 : _GEN_2191; // @[ICache.scala 175:32]
  wire  _GEN_5937 = ~cache_hit ? _GEN_3870 : _GEN_2703; // @[ICache.scala 175:32]
  wire  _GEN_5938 = ~cache_hit ? _GEN_3871 : _GEN_2192; // @[ICache.scala 175:32]
  wire  _GEN_5939 = ~cache_hit ? _GEN_3872 : _GEN_2704; // @[ICache.scala 175:32]
  wire  _GEN_5940 = ~cache_hit ? _GEN_3873 : _GEN_2193; // @[ICache.scala 175:32]
  wire  _GEN_5941 = ~cache_hit ? _GEN_3874 : _GEN_2705; // @[ICache.scala 175:32]
  wire  _GEN_5942 = ~cache_hit ? _GEN_3875 : _GEN_2194; // @[ICache.scala 175:32]
  wire  _GEN_5943 = ~cache_hit ? _GEN_3876 : _GEN_2706; // @[ICache.scala 175:32]
  wire  _GEN_5944 = ~cache_hit ? _GEN_3877 : _GEN_2195; // @[ICache.scala 175:32]
  wire  _GEN_5945 = ~cache_hit ? _GEN_3878 : _GEN_2707; // @[ICache.scala 175:32]
  wire  _GEN_5946 = ~cache_hit ? _GEN_3879 : _GEN_2196; // @[ICache.scala 175:32]
  wire  _GEN_5947 = ~cache_hit ? _GEN_3880 : _GEN_2708; // @[ICache.scala 175:32]
  wire  _GEN_5948 = ~cache_hit ? _GEN_3881 : _GEN_2197; // @[ICache.scala 175:32]
  wire  _GEN_5949 = ~cache_hit ? _GEN_3882 : _GEN_2709; // @[ICache.scala 175:32]
  wire  _GEN_5950 = ~cache_hit ? _GEN_3883 : _GEN_2198; // @[ICache.scala 175:32]
  wire  _GEN_5951 = ~cache_hit ? _GEN_3884 : _GEN_2710; // @[ICache.scala 175:32]
  wire  _GEN_5952 = ~cache_hit ? _GEN_3885 : _GEN_2199; // @[ICache.scala 175:32]
  wire  _GEN_5953 = ~cache_hit ? _GEN_3886 : _GEN_2711; // @[ICache.scala 175:32]
  wire  _GEN_5954 = ~cache_hit ? _GEN_3887 : _GEN_2200; // @[ICache.scala 175:32]
  wire  _GEN_5955 = ~cache_hit ? _GEN_3888 : _GEN_2712; // @[ICache.scala 175:32]
  wire  _GEN_5956 = ~cache_hit ? _GEN_3889 : _GEN_2201; // @[ICache.scala 175:32]
  wire  _GEN_5957 = ~cache_hit ? _GEN_3890 : _GEN_2713; // @[ICache.scala 175:32]
  wire  _GEN_5958 = ~cache_hit ? _GEN_3891 : _GEN_2202; // @[ICache.scala 175:32]
  wire  _GEN_5959 = ~cache_hit ? _GEN_3892 : _GEN_2714; // @[ICache.scala 175:32]
  wire  _GEN_5960 = ~cache_hit ? _GEN_3893 : _GEN_2203; // @[ICache.scala 175:32]
  wire  _GEN_5961 = ~cache_hit ? _GEN_3894 : _GEN_2715; // @[ICache.scala 175:32]
  wire  _GEN_5962 = ~cache_hit ? _GEN_3895 : _GEN_2204; // @[ICache.scala 175:32]
  wire  _GEN_5963 = ~cache_hit ? _GEN_3896 : _GEN_2716; // @[ICache.scala 175:32]
  wire  _GEN_5964 = ~cache_hit ? _GEN_3897 : _GEN_2205; // @[ICache.scala 175:32]
  wire  _GEN_5965 = ~cache_hit ? _GEN_3898 : _GEN_2717; // @[ICache.scala 175:32]
  wire  _GEN_5966 = ~cache_hit ? _GEN_3899 : _GEN_2206; // @[ICache.scala 175:32]
  wire  _GEN_5967 = ~cache_hit ? _GEN_3900 : _GEN_2718; // @[ICache.scala 175:32]
  wire  _GEN_5968 = ~cache_hit ? _GEN_3901 : _GEN_2207; // @[ICache.scala 175:32]
  wire  _GEN_5969 = ~cache_hit ? _GEN_3902 : _GEN_2719; // @[ICache.scala 175:32]
  wire  _GEN_5970 = ~cache_hit ? _GEN_3903 : _GEN_2208; // @[ICache.scala 175:32]
  wire  _GEN_5971 = ~cache_hit ? _GEN_3904 : _GEN_2720; // @[ICache.scala 175:32]
  wire  _GEN_5972 = ~cache_hit ? _GEN_3905 : _GEN_2209; // @[ICache.scala 175:32]
  wire  _GEN_5973 = ~cache_hit ? _GEN_3906 : _GEN_2721; // @[ICache.scala 175:32]
  wire  _GEN_5974 = ~cache_hit ? _GEN_3907 : _GEN_2210; // @[ICache.scala 175:32]
  wire  _GEN_5975 = ~cache_hit ? _GEN_3908 : _GEN_2722; // @[ICache.scala 175:32]
  wire  _GEN_5976 = ~cache_hit ? _GEN_3909 : _GEN_2211; // @[ICache.scala 175:32]
  wire  _GEN_5977 = ~cache_hit ? _GEN_3910 : _GEN_2723; // @[ICache.scala 175:32]
  wire  _GEN_5978 = ~cache_hit ? _GEN_3911 : _GEN_2212; // @[ICache.scala 175:32]
  wire  _GEN_5979 = ~cache_hit ? _GEN_3912 : _GEN_2724; // @[ICache.scala 175:32]
  wire  _GEN_5980 = ~cache_hit ? _GEN_3913 : _GEN_2213; // @[ICache.scala 175:32]
  wire  _GEN_5981 = ~cache_hit ? _GEN_3914 : _GEN_2725; // @[ICache.scala 175:32]
  wire  _GEN_5982 = ~cache_hit ? _GEN_3915 : _GEN_2214; // @[ICache.scala 175:32]
  wire  _GEN_5983 = ~cache_hit ? _GEN_3916 : _GEN_2726; // @[ICache.scala 175:32]
  wire  _GEN_5984 = ~cache_hit ? _GEN_3917 : _GEN_2215; // @[ICache.scala 175:32]
  wire  _GEN_5985 = ~cache_hit ? _GEN_3918 : _GEN_2727; // @[ICache.scala 175:32]
  wire  _GEN_5986 = ~cache_hit ? _GEN_3919 : _GEN_2216; // @[ICache.scala 175:32]
  wire  _GEN_5987 = ~cache_hit ? _GEN_3920 : _GEN_2728; // @[ICache.scala 175:32]
  wire  _GEN_5988 = ~cache_hit ? _GEN_3921 : _GEN_2217; // @[ICache.scala 175:32]
  wire  _GEN_5989 = ~cache_hit ? _GEN_3922 : _GEN_2729; // @[ICache.scala 175:32]
  wire  _GEN_5990 = ~cache_hit ? _GEN_3923 : _GEN_2218; // @[ICache.scala 175:32]
  wire  _GEN_5991 = ~cache_hit ? _GEN_3924 : _GEN_2730; // @[ICache.scala 175:32]
  wire  _GEN_5992 = ~cache_hit ? _GEN_3925 : _GEN_2219; // @[ICache.scala 175:32]
  wire  _GEN_5993 = ~cache_hit ? _GEN_3926 : _GEN_2731; // @[ICache.scala 175:32]
  wire  _GEN_5994 = ~cache_hit ? _GEN_3927 : _GEN_2220; // @[ICache.scala 175:32]
  wire  _GEN_5995 = ~cache_hit ? _GEN_3928 : _GEN_2732; // @[ICache.scala 175:32]
  wire  _GEN_5996 = ~cache_hit ? _GEN_3929 : _GEN_2221; // @[ICache.scala 175:32]
  wire  _GEN_5997 = ~cache_hit ? _GEN_3930 : _GEN_2733; // @[ICache.scala 175:32]
  wire  _GEN_5998 = ~cache_hit ? _GEN_3931 : _GEN_2222; // @[ICache.scala 175:32]
  wire  _GEN_5999 = ~cache_hit ? _GEN_3932 : _GEN_2734; // @[ICache.scala 175:32]
  wire  _GEN_6000 = ~cache_hit ? _GEN_3933 : _GEN_2223; // @[ICache.scala 175:32]
  wire  _GEN_6001 = ~cache_hit ? _GEN_3934 : _GEN_2735; // @[ICache.scala 175:32]
  wire  _GEN_6002 = ~cache_hit ? _GEN_3935 : _GEN_2224; // @[ICache.scala 175:32]
  wire  _GEN_6003 = ~cache_hit ? _GEN_3936 : _GEN_2736; // @[ICache.scala 175:32]
  wire  _GEN_6004 = ~cache_hit ? _GEN_3937 : _GEN_2225; // @[ICache.scala 175:32]
  wire  _GEN_6005 = ~cache_hit ? _GEN_3938 : _GEN_2737; // @[ICache.scala 175:32]
  wire  _GEN_6006 = ~cache_hit ? _GEN_3939 : _GEN_2226; // @[ICache.scala 175:32]
  wire  _GEN_6007 = ~cache_hit ? _GEN_3940 : _GEN_2738; // @[ICache.scala 175:32]
  wire  _GEN_6008 = ~cache_hit ? _GEN_3941 : _GEN_2227; // @[ICache.scala 175:32]
  wire  _GEN_6009 = ~cache_hit ? _GEN_3942 : _GEN_2739; // @[ICache.scala 175:32]
  wire  _GEN_6010 = ~cache_hit ? _GEN_3943 : _GEN_2228; // @[ICache.scala 175:32]
  wire  _GEN_6011 = ~cache_hit ? _GEN_3944 : _GEN_2740; // @[ICache.scala 175:32]
  wire  _GEN_6012 = ~cache_hit ? _GEN_3945 : _GEN_2229; // @[ICache.scala 175:32]
  wire  _GEN_6013 = ~cache_hit ? _GEN_3946 : _GEN_2741; // @[ICache.scala 175:32]
  wire  _GEN_6014 = ~cache_hit ? _GEN_3947 : _GEN_2230; // @[ICache.scala 175:32]
  wire  _GEN_6015 = ~cache_hit ? _GEN_3948 : _GEN_2742; // @[ICache.scala 175:32]
  wire  _GEN_6016 = ~cache_hit ? _GEN_3949 : _GEN_2231; // @[ICache.scala 175:32]
  wire  _GEN_6017 = ~cache_hit ? _GEN_3950 : _GEN_2743; // @[ICache.scala 175:32]
  wire  _GEN_6018 = ~cache_hit ? _GEN_3951 : _GEN_2232; // @[ICache.scala 175:32]
  wire  _GEN_6019 = ~cache_hit ? _GEN_3952 : _GEN_2744; // @[ICache.scala 175:32]
  wire  _GEN_6020 = ~cache_hit ? _GEN_3953 : _GEN_2233; // @[ICache.scala 175:32]
  wire  _GEN_6021 = ~cache_hit ? _GEN_3954 : _GEN_2745; // @[ICache.scala 175:32]
  wire  _GEN_6022 = ~cache_hit ? _GEN_3955 : _GEN_2234; // @[ICache.scala 175:32]
  wire  _GEN_6023 = ~cache_hit ? _GEN_3956 : _GEN_2746; // @[ICache.scala 175:32]
  wire  _GEN_6024 = ~cache_hit ? _GEN_3957 : _GEN_2235; // @[ICache.scala 175:32]
  wire  _GEN_6025 = ~cache_hit ? _GEN_3958 : _GEN_2747; // @[ICache.scala 175:32]
  wire  _GEN_6026 = ~cache_hit ? _GEN_3959 : _GEN_2236; // @[ICache.scala 175:32]
  wire  _GEN_6027 = ~cache_hit ? _GEN_3960 : _GEN_2748; // @[ICache.scala 175:32]
  wire  _GEN_6028 = ~cache_hit ? _GEN_3961 : _GEN_2237; // @[ICache.scala 175:32]
  wire  _GEN_6029 = ~cache_hit ? _GEN_3962 : _GEN_2749; // @[ICache.scala 175:32]
  wire  _GEN_6030 = ~cache_hit ? _GEN_3963 : _GEN_2238; // @[ICache.scala 175:32]
  wire  _GEN_6031 = ~cache_hit ? _GEN_3964 : _GEN_2750; // @[ICache.scala 175:32]
  wire  _GEN_6032 = ~cache_hit ? _GEN_3965 : _GEN_2239; // @[ICache.scala 175:32]
  wire  _GEN_6033 = ~cache_hit ? _GEN_3966 : _GEN_2751; // @[ICache.scala 175:32]
  wire  _GEN_6034 = ~cache_hit ? _GEN_3967 : _GEN_2240; // @[ICache.scala 175:32]
  wire  _GEN_6035 = ~cache_hit ? _GEN_3968 : _GEN_2752; // @[ICache.scala 175:32]
  wire  _GEN_6036 = ~cache_hit ? _GEN_3969 : _GEN_2241; // @[ICache.scala 175:32]
  wire  _GEN_6037 = ~cache_hit ? _GEN_3970 : _GEN_2753; // @[ICache.scala 175:32]
  wire  _GEN_6038 = ~cache_hit ? _GEN_3971 : _GEN_2242; // @[ICache.scala 175:32]
  wire  _GEN_6039 = ~cache_hit ? _GEN_3972 : _GEN_2754; // @[ICache.scala 175:32]
  wire  _GEN_6040 = ~cache_hit ? _GEN_3973 : _GEN_2243; // @[ICache.scala 175:32]
  wire  _GEN_6041 = ~cache_hit ? _GEN_3974 : _GEN_2755; // @[ICache.scala 175:32]
  wire  _GEN_6042 = ~cache_hit ? _GEN_3975 : _GEN_2244; // @[ICache.scala 175:32]
  wire  _GEN_6043 = ~cache_hit ? _GEN_3976 : _GEN_2756; // @[ICache.scala 175:32]
  wire  _GEN_6044 = ~cache_hit ? _GEN_3977 : _GEN_2245; // @[ICache.scala 175:32]
  wire  _GEN_6045 = ~cache_hit ? _GEN_3978 : _GEN_2757; // @[ICache.scala 175:32]
  wire  _GEN_6046 = ~cache_hit ? _GEN_3979 : _GEN_2246; // @[ICache.scala 175:32]
  wire  _GEN_6047 = ~cache_hit ? _GEN_3980 : _GEN_2758; // @[ICache.scala 175:32]
  wire  _GEN_6048 = ~cache_hit ? _GEN_3981 : _GEN_2247; // @[ICache.scala 175:32]
  wire  _GEN_6049 = ~cache_hit ? _GEN_3982 : _GEN_2759; // @[ICache.scala 175:32]
  wire  _GEN_6050 = ~cache_hit ? _GEN_3983 : _GEN_2248; // @[ICache.scala 175:32]
  wire  _GEN_6051 = ~cache_hit ? _GEN_3984 : _GEN_2760; // @[ICache.scala 175:32]
  wire  _GEN_6052 = ~cache_hit ? _GEN_3985 : _GEN_2249; // @[ICache.scala 175:32]
  wire  _GEN_6053 = ~cache_hit ? _GEN_3986 : _GEN_2761; // @[ICache.scala 175:32]
  wire  _GEN_6054 = ~cache_hit ? _GEN_3987 : _GEN_2250; // @[ICache.scala 175:32]
  wire  _GEN_6055 = ~cache_hit ? _GEN_3988 : _GEN_2762; // @[ICache.scala 175:32]
  wire  _GEN_6056 = ~cache_hit ? _GEN_3989 : _GEN_2251; // @[ICache.scala 175:32]
  wire  _GEN_6057 = ~cache_hit ? _GEN_3990 : _GEN_2763; // @[ICache.scala 175:32]
  wire  _GEN_6058 = ~cache_hit ? _GEN_3991 : _GEN_2252; // @[ICache.scala 175:32]
  wire  _GEN_6059 = ~cache_hit ? _GEN_3992 : _GEN_2764; // @[ICache.scala 175:32]
  wire  _GEN_6060 = ~cache_hit ? _GEN_3993 : _GEN_2253; // @[ICache.scala 175:32]
  wire  _GEN_6061 = ~cache_hit ? _GEN_3994 : _GEN_2765; // @[ICache.scala 175:32]
  wire  _GEN_6062 = ~cache_hit ? _GEN_3995 : _GEN_2254; // @[ICache.scala 175:32]
  wire  _GEN_6063 = ~cache_hit ? _GEN_3996 : _GEN_2766; // @[ICache.scala 175:32]
  wire  _GEN_6064 = ~cache_hit ? _GEN_3997 : _GEN_2255; // @[ICache.scala 175:32]
  wire  _GEN_6065 = ~cache_hit ? _GEN_3998 : _GEN_2767; // @[ICache.scala 175:32]
  wire  _GEN_6066 = ~cache_hit ? _GEN_3999 : _GEN_2256; // @[ICache.scala 175:32]
  wire  _GEN_6067 = ~cache_hit ? _GEN_4000 : _GEN_2768; // @[ICache.scala 175:32]
  wire  _GEN_6068 = ~cache_hit ? _GEN_4001 : _GEN_2257; // @[ICache.scala 175:32]
  wire  _GEN_6069 = ~cache_hit ? _GEN_4002 : _GEN_2769; // @[ICache.scala 175:32]
  wire  _GEN_6070 = ~cache_hit ? _GEN_4003 : _GEN_2258; // @[ICache.scala 175:32]
  wire  _GEN_6071 = ~cache_hit ? _GEN_4004 : _GEN_2770; // @[ICache.scala 175:32]
  wire  _GEN_6072 = ~cache_hit ? _GEN_4005 : _GEN_2259; // @[ICache.scala 175:32]
  wire  _GEN_6073 = ~cache_hit ? _GEN_4006 : _GEN_2771; // @[ICache.scala 175:32]
  wire  _GEN_6074 = ~cache_hit ? _GEN_4007 : _GEN_2260; // @[ICache.scala 175:32]
  wire  _GEN_6075 = ~cache_hit ? _GEN_4008 : _GEN_2772; // @[ICache.scala 175:32]
  wire  _GEN_6076 = ~cache_hit ? _GEN_4009 : _GEN_2261; // @[ICache.scala 175:32]
  wire  _GEN_6077 = ~cache_hit ? _GEN_4010 : _GEN_2773; // @[ICache.scala 175:32]
  wire  _GEN_6078 = ~cache_hit ? _GEN_4011 : _GEN_2262; // @[ICache.scala 175:32]
  wire  _GEN_6079 = ~cache_hit ? _GEN_4012 : _GEN_2774; // @[ICache.scala 175:32]
  wire  _GEN_6080 = ~cache_hit ? _GEN_4013 : _GEN_2263; // @[ICache.scala 175:32]
  wire  _GEN_6081 = ~cache_hit ? _GEN_4014 : _GEN_2775; // @[ICache.scala 175:32]
  wire  _GEN_6082 = ~cache_hit ? _GEN_4015 : _GEN_2264; // @[ICache.scala 175:32]
  wire  _GEN_6083 = ~cache_hit ? _GEN_4016 : _GEN_2776; // @[ICache.scala 175:32]
  wire  _GEN_6084 = ~cache_hit ? _GEN_4017 : _GEN_2265; // @[ICache.scala 175:32]
  wire  _GEN_6085 = ~cache_hit ? _GEN_4018 : _GEN_2777; // @[ICache.scala 175:32]
  wire  _GEN_6086 = ~cache_hit ? _GEN_4019 : _GEN_2266; // @[ICache.scala 175:32]
  wire  _GEN_6087 = ~cache_hit ? _GEN_4020 : _GEN_2778; // @[ICache.scala 175:32]
  wire  _GEN_6088 = ~cache_hit ? _GEN_4021 : _GEN_2267; // @[ICache.scala 175:32]
  wire  _GEN_6089 = ~cache_hit ? _GEN_4022 : _GEN_2779; // @[ICache.scala 175:32]
  wire  _GEN_6090 = ~cache_hit ? _GEN_4023 : _GEN_2268; // @[ICache.scala 175:32]
  wire  _GEN_6091 = ~cache_hit ? _GEN_4024 : _GEN_2780; // @[ICache.scala 175:32]
  wire  _GEN_6092 = ~cache_hit ? _GEN_4025 : _GEN_2269; // @[ICache.scala 175:32]
  wire  _GEN_6093 = ~cache_hit ? _GEN_4026 : _GEN_2781; // @[ICache.scala 175:32]
  wire  _GEN_6094 = ~cache_hit ? _GEN_4027 : _GEN_2270; // @[ICache.scala 175:32]
  wire  _GEN_6095 = ~cache_hit ? _GEN_4028 : _GEN_2782; // @[ICache.scala 175:32]
  wire  _GEN_6096 = ~cache_hit ? _GEN_4029 : _GEN_2271; // @[ICache.scala 175:32]
  wire  _GEN_6097 = ~cache_hit ? _GEN_4030 : _GEN_2783; // @[ICache.scala 175:32]
  wire  _GEN_6098 = ~cache_hit ? _GEN_4031 : _GEN_2272; // @[ICache.scala 175:32]
  wire  _GEN_6099 = ~cache_hit ? _GEN_4032 : _GEN_2784; // @[ICache.scala 175:32]
  wire  _GEN_6100 = ~cache_hit ? _GEN_4033 : _GEN_2273; // @[ICache.scala 175:32]
  wire  _GEN_6101 = ~cache_hit ? _GEN_4034 : _GEN_2785; // @[ICache.scala 175:32]
  wire  _GEN_6102 = ~cache_hit ? _GEN_4035 : _GEN_2274; // @[ICache.scala 175:32]
  wire  _GEN_6103 = ~cache_hit ? _GEN_4036 : _GEN_2786; // @[ICache.scala 175:32]
  wire  _GEN_6104 = ~cache_hit ? _GEN_4037 : _GEN_2275; // @[ICache.scala 175:32]
  wire  _GEN_6105 = ~cache_hit ? _GEN_4038 : _GEN_2787; // @[ICache.scala 175:32]
  wire  _GEN_6106 = ~cache_hit ? _GEN_4039 : _GEN_2276; // @[ICache.scala 175:32]
  wire  _GEN_6107 = ~cache_hit ? _GEN_4040 : _GEN_2788; // @[ICache.scala 175:32]
  wire  _GEN_6108 = ~cache_hit ? _GEN_4041 : _GEN_2277; // @[ICache.scala 175:32]
  wire  _GEN_6109 = ~cache_hit ? _GEN_4042 : _GEN_2789; // @[ICache.scala 175:32]
  wire  _GEN_6110 = ~cache_hit ? _GEN_4043 : _GEN_2278; // @[ICache.scala 175:32]
  wire  _GEN_6111 = ~cache_hit ? _GEN_4044 : _GEN_2790; // @[ICache.scala 175:32]
  wire  _GEN_6112 = ~cache_hit ? _GEN_4045 : _GEN_2279; // @[ICache.scala 175:32]
  wire  _GEN_6113 = ~cache_hit ? _GEN_4046 : _GEN_2791; // @[ICache.scala 175:32]
  wire  _GEN_6114 = ~cache_hit ? _GEN_4047 : _GEN_2280; // @[ICache.scala 175:32]
  wire  _GEN_6115 = ~cache_hit ? _GEN_4048 : _GEN_2792; // @[ICache.scala 175:32]
  wire  _GEN_6116 = ~cache_hit ? _GEN_4049 : _GEN_2281; // @[ICache.scala 175:32]
  wire  _GEN_6117 = ~cache_hit ? _GEN_4050 : _GEN_2793; // @[ICache.scala 175:32]
  wire  _GEN_6118 = ~cache_hit ? _GEN_4051 : _GEN_2282; // @[ICache.scala 175:32]
  wire  _GEN_6119 = ~cache_hit ? _GEN_4052 : _GEN_2794; // @[ICache.scala 175:32]
  wire  _GEN_6120 = ~cache_hit ? _GEN_4053 : _GEN_2283; // @[ICache.scala 175:32]
  wire  _GEN_6121 = ~cache_hit ? _GEN_4054 : _GEN_2795; // @[ICache.scala 175:32]
  wire  _GEN_6122 = ~cache_hit ? _GEN_4055 : _GEN_2284; // @[ICache.scala 175:32]
  wire  _GEN_6123 = ~cache_hit ? _GEN_4056 : _GEN_2796; // @[ICache.scala 175:32]
  wire  _GEN_6124 = ~cache_hit ? _GEN_4057 : _GEN_2285; // @[ICache.scala 175:32]
  wire  _GEN_6125 = ~cache_hit ? _GEN_4058 : _GEN_2797; // @[ICache.scala 175:32]
  wire  _GEN_6126 = ~cache_hit ? _GEN_4059 : _GEN_2286; // @[ICache.scala 175:32]
  wire  _GEN_6127 = ~cache_hit ? _GEN_4060 : _GEN_2798; // @[ICache.scala 175:32]
  wire  _GEN_6128 = ~cache_hit ? _GEN_4061 : _GEN_2287; // @[ICache.scala 175:32]
  wire  _GEN_6129 = ~cache_hit ? _GEN_4062 : _GEN_2799; // @[ICache.scala 175:32]
  wire  _GEN_6130 = ~cache_hit ? _GEN_4063 : _GEN_2288; // @[ICache.scala 175:32]
  wire  _GEN_6131 = ~cache_hit ? _GEN_4064 : _GEN_2800; // @[ICache.scala 175:32]
  wire  _GEN_6132 = ~cache_hit ? _GEN_4065 : _GEN_2289; // @[ICache.scala 175:32]
  wire  _GEN_6133 = ~cache_hit ? _GEN_4066 : _GEN_2801; // @[ICache.scala 175:32]
  wire  _GEN_6134 = ~cache_hit ? _GEN_4067 : _GEN_2290; // @[ICache.scala 175:32]
  wire  _GEN_6135 = ~cache_hit ? _GEN_4068 : _GEN_2802; // @[ICache.scala 175:32]
  wire  _GEN_6136 = ~cache_hit ? _GEN_4069 : _GEN_2291; // @[ICache.scala 175:32]
  wire  _GEN_6137 = ~cache_hit ? _GEN_4070 : _GEN_2803; // @[ICache.scala 175:32]
  wire  _GEN_6138 = ~cache_hit ? _GEN_4071 : _GEN_2292; // @[ICache.scala 175:32]
  wire  _GEN_6139 = ~cache_hit ? _GEN_4072 : _GEN_2804; // @[ICache.scala 175:32]
  wire  _GEN_6140 = ~cache_hit ? _GEN_4073 : _GEN_2293; // @[ICache.scala 175:32]
  wire  _GEN_6141 = ~cache_hit ? _GEN_4074 : _GEN_2805; // @[ICache.scala 175:32]
  wire  _GEN_6142 = ~cache_hit ? _GEN_4075 : _GEN_2294; // @[ICache.scala 175:32]
  wire  _GEN_6143 = ~cache_hit ? _GEN_4076 : _GEN_2806; // @[ICache.scala 175:32]
  wire  _GEN_6144 = ~cache_hit ? _GEN_4077 : _GEN_2295; // @[ICache.scala 175:32]
  wire  _GEN_6145 = ~cache_hit ? _GEN_4078 : _GEN_2807; // @[ICache.scala 175:32]
  wire  _GEN_6146 = ~cache_hit ? _GEN_4079 : _GEN_2296; // @[ICache.scala 175:32]
  wire  _GEN_6147 = ~cache_hit ? _GEN_4080 : _GEN_2808; // @[ICache.scala 175:32]
  wire  _GEN_6148 = ~cache_hit ? _GEN_4081 : _GEN_2297; // @[ICache.scala 175:32]
  wire  _GEN_6149 = ~cache_hit ? _GEN_4082 : _GEN_2809; // @[ICache.scala 175:32]
  wire  _GEN_6150 = ~cache_hit ? _GEN_4083 : _GEN_2298; // @[ICache.scala 175:32]
  wire  _GEN_6151 = ~cache_hit ? _GEN_4084 : _GEN_2810; // @[ICache.scala 175:32]
  wire  _GEN_6152 = ~cache_hit ? _GEN_4085 : _GEN_2299; // @[ICache.scala 175:32]
  wire  _GEN_6153 = ~cache_hit ? _GEN_4086 : _GEN_2811; // @[ICache.scala 175:32]
  wire  _GEN_6154 = ~cache_hit ? _GEN_4087 : _GEN_2300; // @[ICache.scala 175:32]
  wire  _GEN_6155 = ~cache_hit ? _GEN_4088 : _GEN_2812; // @[ICache.scala 175:32]
  wire  _GEN_6156 = ~cache_hit ? _GEN_4089 : _GEN_2301; // @[ICache.scala 175:32]
  wire  _GEN_6157 = ~cache_hit ? _GEN_4090 : _GEN_2813; // @[ICache.scala 175:32]
  wire  _GEN_6158 = ~cache_hit ? _GEN_4091 : _GEN_2302; // @[ICache.scala 175:32]
  wire  _GEN_6159 = ~cache_hit ? _GEN_4092 : _GEN_2814; // @[ICache.scala 175:32]
  wire  _GEN_6160 = ~cache_hit ? _GEN_4093 : _GEN_2303; // @[ICache.scala 175:32]
  wire  _GEN_6161 = ~cache_hit ? _GEN_4094 : _GEN_2815; // @[ICache.scala 175:32]
  wire  _GEN_6162 = ~cache_hit ? _GEN_4095 : _GEN_2304; // @[ICache.scala 175:32]
  wire  _GEN_6163 = ~cache_hit ? _GEN_4096 : _GEN_2816; // @[ICache.scala 175:32]
  wire  _GEN_6164 = ~cache_hit ? _GEN_4097 : _GEN_2305; // @[ICache.scala 175:32]
  wire  _GEN_6165 = ~cache_hit ? _GEN_4098 : _GEN_2817; // @[ICache.scala 175:32]
  wire  _GEN_6166 = ~cache_hit ? _GEN_4099 : _GEN_2306; // @[ICache.scala 175:32]
  wire  _GEN_6167 = ~cache_hit ? _GEN_4100 : _GEN_2818; // @[ICache.scala 175:32]
  wire  _GEN_6168 = ~cache_hit ? _GEN_4101 : _GEN_2307; // @[ICache.scala 175:32]
  wire  _GEN_6169 = ~cache_hit ? _GEN_4102 : _GEN_2819; // @[ICache.scala 175:32]
  wire  _GEN_6170 = ~cache_hit ? _GEN_4103 : _GEN_2308; // @[ICache.scala 175:32]
  wire  _GEN_6171 = ~cache_hit ? _GEN_4104 : _GEN_2820; // @[ICache.scala 175:32]
  wire  _GEN_6172 = ~cache_hit ? _GEN_4105 : _GEN_2309; // @[ICache.scala 175:32]
  wire  _GEN_6173 = ~cache_hit ? _GEN_4106 : _GEN_2821; // @[ICache.scala 175:32]
  wire  _GEN_6174 = ~cache_hit ? _GEN_4107 : _GEN_2310; // @[ICache.scala 175:32]
  wire  _GEN_6175 = ~cache_hit ? _GEN_4108 : _GEN_2822; // @[ICache.scala 175:32]
  wire  _GEN_6176 = ~cache_hit ? _GEN_4109 : _GEN_2311; // @[ICache.scala 175:32]
  wire  _GEN_6177 = ~cache_hit ? _GEN_4110 : _GEN_2823; // @[ICache.scala 175:32]
  wire  _GEN_6178 = ~cache_hit ? _GEN_4111 : _GEN_2312; // @[ICache.scala 175:32]
  wire  _GEN_6179 = ~cache_hit ? _GEN_4112 : _GEN_2824; // @[ICache.scala 175:32]
  wire  _GEN_6180 = ~cache_hit ? _GEN_4113 : _GEN_2313; // @[ICache.scala 175:32]
  wire  _GEN_6181 = ~cache_hit ? _GEN_4114 : _GEN_2825; // @[ICache.scala 175:32]
  wire  _GEN_6182 = ~cache_hit ? _GEN_4115 : _GEN_2314; // @[ICache.scala 175:32]
  wire  _GEN_6183 = ~cache_hit ? _GEN_4116 : _GEN_2826; // @[ICache.scala 175:32]
  wire  _GEN_6184 = ~cache_hit ? _GEN_4117 : _GEN_2315; // @[ICache.scala 175:32]
  wire  _GEN_6185 = ~cache_hit ? _GEN_4118 : _GEN_2827; // @[ICache.scala 175:32]
  wire  _GEN_6186 = ~cache_hit ? _GEN_4119 : _GEN_2316; // @[ICache.scala 175:32]
  wire  _GEN_6187 = ~cache_hit ? _GEN_4120 : _GEN_2828; // @[ICache.scala 175:32]
  wire  _GEN_6188 = ~cache_hit ? _GEN_4121 : _GEN_2317; // @[ICache.scala 175:32]
  wire  _GEN_6189 = ~cache_hit ? _GEN_4122 : _GEN_2829; // @[ICache.scala 175:32]
  wire  _GEN_6190 = ~cache_hit ? _GEN_4123 : _GEN_2318; // @[ICache.scala 175:32]
  wire  _GEN_6191 = ~cache_hit ? _GEN_4124 : _GEN_2830; // @[ICache.scala 175:32]
  wire  _GEN_6192 = ~cache_hit ? _GEN_4125 : _GEN_2319; // @[ICache.scala 175:32]
  wire  _GEN_6193 = ~cache_hit ? _GEN_4126 : _GEN_2831; // @[ICache.scala 175:32]
  wire  _GEN_6194 = ~cache_hit ? _GEN_4127 : _GEN_2320; // @[ICache.scala 175:32]
  wire  _GEN_6195 = ~cache_hit ? _GEN_4128 : _GEN_2832; // @[ICache.scala 175:32]
  wire  _GEN_6196 = ~cache_hit ? _GEN_4129 : _GEN_2321; // @[ICache.scala 175:32]
  wire  _GEN_6197 = ~cache_hit ? _GEN_4130 : _GEN_2833; // @[ICache.scala 175:32]
  wire  _GEN_6198 = ~cache_hit ? _GEN_4131 : _GEN_2322; // @[ICache.scala 175:32]
  wire  _GEN_6199 = ~cache_hit ? _GEN_4132 : _GEN_2834; // @[ICache.scala 175:32]
  wire  _GEN_6200 = ~cache_hit ? _GEN_4133 : _GEN_2323; // @[ICache.scala 175:32]
  wire  _GEN_6201 = ~cache_hit ? _GEN_4134 : _GEN_2835; // @[ICache.scala 175:32]
  wire  _GEN_6202 = ~cache_hit ? _GEN_4135 : _GEN_2324; // @[ICache.scala 175:32]
  wire  _GEN_6203 = ~cache_hit ? _GEN_4136 : _GEN_2836; // @[ICache.scala 175:32]
  wire  _GEN_6204 = ~cache_hit ? _GEN_4137 : _GEN_2325; // @[ICache.scala 175:32]
  wire  _GEN_6205 = ~cache_hit ? _GEN_4138 : _GEN_2837; // @[ICache.scala 175:32]
  wire  _GEN_6206 = ~cache_hit ? _GEN_4139 : _GEN_2326; // @[ICache.scala 175:32]
  wire  _GEN_6207 = ~cache_hit ? _GEN_4140 : _GEN_2838; // @[ICache.scala 175:32]
  wire  _GEN_6208 = ~cache_hit ? _GEN_4141 : _GEN_2327; // @[ICache.scala 175:32]
  wire  _GEN_6209 = ~cache_hit ? _GEN_4142 : _GEN_2839; // @[ICache.scala 175:32]
  wire  _GEN_6210 = ~cache_hit ? _GEN_4143 : _GEN_2328; // @[ICache.scala 175:32]
  wire  _GEN_6211 = ~cache_hit ? _GEN_4144 : _GEN_2840; // @[ICache.scala 175:32]
  wire  _GEN_6212 = ~cache_hit ? _GEN_4145 : _GEN_2329; // @[ICache.scala 175:32]
  wire  _GEN_6213 = ~cache_hit ? _GEN_4146 : _GEN_2841; // @[ICache.scala 175:32]
  wire  _GEN_6214 = ~cache_hit ? _GEN_4147 : _GEN_2330; // @[ICache.scala 175:32]
  wire  _GEN_6215 = ~cache_hit ? _GEN_4148 : _GEN_2842; // @[ICache.scala 175:32]
  wire  _GEN_6216 = ~cache_hit ? _GEN_4149 : _GEN_2331; // @[ICache.scala 175:32]
  wire  _GEN_6217 = ~cache_hit ? _GEN_4150 : _GEN_2843; // @[ICache.scala 175:32]
  wire  _GEN_6218 = ~cache_hit ? _GEN_4151 : _GEN_2332; // @[ICache.scala 175:32]
  wire  _GEN_6219 = ~cache_hit ? _GEN_4152 : _GEN_2844; // @[ICache.scala 175:32]
  wire  _GEN_6220 = ~cache_hit ? _GEN_4153 : _GEN_2333; // @[ICache.scala 175:32]
  wire  _GEN_6221 = ~cache_hit ? _GEN_4154 : _GEN_2845; // @[ICache.scala 175:32]
  wire  _GEN_6222 = ~cache_hit ? _GEN_4155 : _GEN_2334; // @[ICache.scala 175:32]
  wire  _GEN_6223 = ~cache_hit ? _GEN_4156 : _GEN_2846; // @[ICache.scala 175:32]
  wire  _GEN_6224 = ~cache_hit ? _GEN_4157 : _GEN_2335; // @[ICache.scala 175:32]
  wire  _GEN_6225 = ~cache_hit ? _GEN_4158 : _GEN_2847; // @[ICache.scala 175:32]
  wire  _GEN_6226 = ~cache_hit ? _GEN_4159 : _GEN_2336; // @[ICache.scala 175:32]
  wire  _GEN_6227 = ~cache_hit ? _GEN_4160 : _GEN_2848; // @[ICache.scala 175:32]
  wire  _GEN_6228 = ~cache_hit ? _GEN_4161 : _GEN_2337; // @[ICache.scala 175:32]
  wire  _GEN_6229 = ~cache_hit ? _GEN_4162 : _GEN_2849; // @[ICache.scala 175:32]
  wire  _GEN_6230 = ~cache_hit ? _GEN_4163 : _GEN_2338; // @[ICache.scala 175:32]
  wire  _GEN_6231 = ~cache_hit ? _GEN_4164 : _GEN_2850; // @[ICache.scala 175:32]
  wire  _GEN_6232 = ~cache_hit ? _GEN_4165 : _GEN_2339; // @[ICache.scala 175:32]
  wire  _GEN_6233 = ~cache_hit ? _GEN_4166 : _GEN_2851; // @[ICache.scala 175:32]
  wire  _GEN_6234 = ~cache_hit ? _GEN_4167 : _GEN_2340; // @[ICache.scala 175:32]
  wire  _GEN_6235 = ~cache_hit ? _GEN_4168 : _GEN_2852; // @[ICache.scala 175:32]
  wire  _GEN_6236 = ~cache_hit ? _GEN_4169 : _GEN_2341; // @[ICache.scala 175:32]
  wire  _GEN_6237 = ~cache_hit ? _GEN_4170 : _GEN_2853; // @[ICache.scala 175:32]
  wire  _GEN_6238 = ~cache_hit ? _GEN_4171 : _GEN_2342; // @[ICache.scala 175:32]
  wire  _GEN_6239 = ~cache_hit ? _GEN_4172 : _GEN_2854; // @[ICache.scala 175:32]
  wire  _GEN_6240 = ~cache_hit ? _GEN_4173 : _GEN_2343; // @[ICache.scala 175:32]
  wire  _GEN_6241 = ~cache_hit ? _GEN_4174 : _GEN_2855; // @[ICache.scala 175:32]
  wire  _GEN_6242 = ~cache_hit ? _GEN_4175 : _GEN_2344; // @[ICache.scala 175:32]
  wire  _GEN_6243 = ~cache_hit ? _GEN_4176 : _GEN_2856; // @[ICache.scala 175:32]
  wire  _GEN_6244 = ~cache_hit ? _GEN_4177 : _GEN_2345; // @[ICache.scala 175:32]
  wire  _GEN_6245 = ~cache_hit ? _GEN_4178 : _GEN_2857; // @[ICache.scala 175:32]
  wire  _GEN_6246 = ~cache_hit ? _GEN_4179 : _GEN_2346; // @[ICache.scala 175:32]
  wire  _GEN_6247 = ~cache_hit ? _GEN_4180 : _GEN_2858; // @[ICache.scala 175:32]
  wire  _GEN_6248 = ~cache_hit ? _GEN_4181 : _GEN_2347; // @[ICache.scala 175:32]
  wire  _GEN_6249 = ~cache_hit ? _GEN_4182 : _GEN_2859; // @[ICache.scala 175:32]
  wire  _GEN_6250 = ~cache_hit ? _GEN_4183 : _GEN_2348; // @[ICache.scala 175:32]
  wire  _GEN_6251 = ~cache_hit ? _GEN_4184 : _GEN_2860; // @[ICache.scala 175:32]
  wire  _GEN_6252 = ~cache_hit ? _GEN_4185 : _GEN_2349; // @[ICache.scala 175:32]
  wire  _GEN_6253 = ~cache_hit ? _GEN_4186 : _GEN_2861; // @[ICache.scala 175:32]
  wire  _GEN_6254 = ~cache_hit ? _GEN_4187 : _GEN_2350; // @[ICache.scala 175:32]
  wire  _GEN_6255 = ~cache_hit ? _GEN_4188 : _GEN_2862; // @[ICache.scala 175:32]
  wire  _GEN_6256 = ~cache_hit ? _GEN_4189 : _GEN_2351; // @[ICache.scala 175:32]
  wire  _GEN_6257 = ~cache_hit ? _GEN_4190 : _GEN_2863; // @[ICache.scala 175:32]
  wire  _GEN_6258 = ~cache_hit ? _GEN_4191 : _GEN_2352; // @[ICache.scala 175:32]
  wire  _GEN_6259 = ~cache_hit ? _GEN_4192 : _GEN_2864; // @[ICache.scala 175:32]
  wire  _GEN_6260 = ~cache_hit ? _GEN_4193 : _GEN_2353; // @[ICache.scala 175:32]
  wire  _GEN_6261 = ~cache_hit ? _GEN_4194 : _GEN_2865; // @[ICache.scala 175:32]
  wire  _GEN_6262 = ~cache_hit ? _GEN_4195 : _GEN_2354; // @[ICache.scala 175:32]
  wire  _GEN_6263 = ~cache_hit ? _GEN_4196 : _GEN_2866; // @[ICache.scala 175:32]
  wire  _GEN_6264 = ~cache_hit ? _GEN_4197 : _GEN_2355; // @[ICache.scala 175:32]
  wire  _GEN_6265 = ~cache_hit ? _GEN_4198 : _GEN_2867; // @[ICache.scala 175:32]
  wire  _GEN_6266 = ~cache_hit ? _GEN_4199 : _GEN_2356; // @[ICache.scala 175:32]
  wire  _GEN_6267 = ~cache_hit ? _GEN_4200 : _GEN_2868; // @[ICache.scala 175:32]
  wire  _GEN_6268 = ~cache_hit ? _GEN_4201 : _GEN_2357; // @[ICache.scala 175:32]
  wire  _GEN_6269 = ~cache_hit ? _GEN_4202 : _GEN_2869; // @[ICache.scala 175:32]
  wire  _GEN_6270 = ~cache_hit ? _GEN_4203 : _GEN_2358; // @[ICache.scala 175:32]
  wire  _GEN_6271 = ~cache_hit ? _GEN_4204 : _GEN_2870; // @[ICache.scala 175:32]
  wire  _GEN_6272 = ~cache_hit ? _GEN_4205 : _GEN_2359; // @[ICache.scala 175:32]
  wire  _GEN_6273 = ~cache_hit ? _GEN_4206 : _GEN_2871; // @[ICache.scala 175:32]
  wire  _GEN_6274 = ~cache_hit ? _GEN_4207 : _GEN_2360; // @[ICache.scala 175:32]
  wire  _GEN_6275 = ~cache_hit ? _GEN_4208 : _GEN_2872; // @[ICache.scala 175:32]
  wire  _GEN_6276 = ~cache_hit ? _GEN_4209 : _GEN_2361; // @[ICache.scala 175:32]
  wire  _GEN_6277 = ~cache_hit ? _GEN_4210 : _GEN_2873; // @[ICache.scala 175:32]
  wire  _GEN_6278 = ~cache_hit ? _GEN_4211 : _GEN_2362; // @[ICache.scala 175:32]
  wire  _GEN_6279 = ~cache_hit ? _GEN_4212 : _GEN_2874; // @[ICache.scala 175:32]
  wire  _GEN_6280 = ~cache_hit ? _GEN_4213 : _GEN_2363; // @[ICache.scala 175:32]
  wire  _GEN_6281 = ~cache_hit ? _GEN_4214 : _GEN_2875; // @[ICache.scala 175:32]
  wire  _GEN_6282 = ~cache_hit ? _GEN_4215 : _GEN_2364; // @[ICache.scala 175:32]
  wire  _GEN_6283 = ~cache_hit ? _GEN_4216 : _GEN_2876; // @[ICache.scala 175:32]
  wire  _GEN_6284 = ~cache_hit ? _GEN_4217 : _GEN_2365; // @[ICache.scala 175:32]
  wire  _GEN_6285 = ~cache_hit ? _GEN_4218 : _GEN_2877; // @[ICache.scala 175:32]
  wire  _GEN_6286 = ~cache_hit ? _GEN_4219 : _GEN_2366; // @[ICache.scala 175:32]
  wire  _GEN_6287 = ~cache_hit ? _GEN_4220 : _GEN_2878; // @[ICache.scala 175:32]
  wire  _GEN_6288 = ~cache_hit ? _GEN_4221 : _GEN_2367; // @[ICache.scala 175:32]
  wire  _GEN_6289 = ~cache_hit ? _GEN_4222 : _GEN_2879; // @[ICache.scala 175:32]
  wire  _GEN_6290 = ~cache_hit ? _GEN_4223 : _GEN_2368; // @[ICache.scala 175:32]
  wire  _GEN_6291 = ~cache_hit ? _GEN_4224 : _GEN_2880; // @[ICache.scala 175:32]
  wire  _GEN_6292 = ~cache_hit ? _GEN_4225 : _GEN_2369; // @[ICache.scala 175:32]
  wire  _GEN_6293 = ~cache_hit ? _GEN_4226 : _GEN_2881; // @[ICache.scala 175:32]
  wire  _GEN_6294 = ~cache_hit ? _GEN_4227 : _GEN_2370; // @[ICache.scala 175:32]
  wire  _GEN_6295 = ~cache_hit ? _GEN_4228 : _GEN_2882; // @[ICache.scala 175:32]
  wire  _GEN_6296 = ~cache_hit ? _GEN_4229 : _GEN_2371; // @[ICache.scala 175:32]
  wire  _GEN_6297 = ~cache_hit ? _GEN_4230 : _GEN_2883; // @[ICache.scala 175:32]
  wire  _GEN_6298 = ~cache_hit ? _GEN_4231 : _GEN_2372; // @[ICache.scala 175:32]
  wire  _GEN_6299 = ~cache_hit ? _GEN_4232 : _GEN_2884; // @[ICache.scala 175:32]
  wire  _GEN_6300 = ~cache_hit ? _GEN_4233 : _GEN_2373; // @[ICache.scala 175:32]
  wire  _GEN_6301 = ~cache_hit ? _GEN_4234 : _GEN_2885; // @[ICache.scala 175:32]
  wire  _GEN_6302 = ~cache_hit ? _GEN_4235 : _GEN_2374; // @[ICache.scala 175:32]
  wire  _GEN_6303 = ~cache_hit ? _GEN_4236 : _GEN_2886; // @[ICache.scala 175:32]
  wire  _GEN_6304 = ~cache_hit ? _GEN_4237 : _GEN_2375; // @[ICache.scala 175:32]
  wire  _GEN_6305 = ~cache_hit ? _GEN_4238 : _GEN_2887; // @[ICache.scala 175:32]
  wire  _GEN_6306 = ~cache_hit ? _GEN_4239 : _GEN_2376; // @[ICache.scala 175:32]
  wire  _GEN_6307 = ~cache_hit ? _GEN_4240 : _GEN_2888; // @[ICache.scala 175:32]
  wire  _GEN_6308 = ~cache_hit ? _GEN_4241 : _GEN_2377; // @[ICache.scala 175:32]
  wire  _GEN_6309 = ~cache_hit ? _GEN_4242 : _GEN_2889; // @[ICache.scala 175:32]
  wire  _GEN_6310 = ~cache_hit ? _GEN_4243 : _GEN_2378; // @[ICache.scala 175:32]
  wire  _GEN_6311 = ~cache_hit ? _GEN_4244 : _GEN_2890; // @[ICache.scala 175:32]
  wire  _GEN_6312 = ~cache_hit ? _GEN_4245 : _GEN_2379; // @[ICache.scala 175:32]
  wire  _GEN_6313 = ~cache_hit ? _GEN_4246 : _GEN_2891; // @[ICache.scala 175:32]
  wire  _GEN_6314 = ~cache_hit ? _GEN_4247 : _GEN_2380; // @[ICache.scala 175:32]
  wire  _GEN_6315 = ~cache_hit ? _GEN_4248 : _GEN_2892; // @[ICache.scala 175:32]
  wire  _GEN_6316 = ~cache_hit ? _GEN_4249 : _GEN_2381; // @[ICache.scala 175:32]
  wire  _GEN_6317 = ~cache_hit ? _GEN_4250 : _GEN_2893; // @[ICache.scala 175:32]
  wire  _GEN_6318 = ~cache_hit ? _GEN_4251 : _GEN_2382; // @[ICache.scala 175:32]
  wire  _GEN_6319 = ~cache_hit ? _GEN_4252 : _GEN_2894; // @[ICache.scala 175:32]
  wire  _GEN_6320 = ~cache_hit ? _GEN_4253 : _GEN_2383; // @[ICache.scala 175:32]
  wire  _GEN_6321 = ~cache_hit ? _GEN_4254 : _GEN_2895; // @[ICache.scala 175:32]
  wire  _GEN_6322 = ~cache_hit ? _GEN_4255 : _GEN_2384; // @[ICache.scala 175:32]
  wire  _GEN_6323 = ~cache_hit ? _GEN_4256 : _GEN_2896; // @[ICache.scala 175:32]
  wire  _GEN_6324 = ~cache_hit ? _GEN_4257 : _GEN_2385; // @[ICache.scala 175:32]
  wire  _GEN_6325 = ~cache_hit ? _GEN_4258 : _GEN_2897; // @[ICache.scala 175:32]
  wire  _GEN_6326 = ~cache_hit ? _GEN_4259 : _GEN_2386; // @[ICache.scala 175:32]
  wire  _GEN_6327 = ~cache_hit ? _GEN_4260 : _GEN_2898; // @[ICache.scala 175:32]
  wire  _GEN_6328 = ~cache_hit ? _GEN_4261 : _GEN_2387; // @[ICache.scala 175:32]
  wire  _GEN_6329 = ~cache_hit ? _GEN_4262 : _GEN_2899; // @[ICache.scala 175:32]
  wire  _GEN_6330 = ~cache_hit ? _GEN_4263 : _GEN_2388; // @[ICache.scala 175:32]
  wire  _GEN_6331 = ~cache_hit ? _GEN_4264 : _GEN_2900; // @[ICache.scala 175:32]
  wire  _GEN_6332 = ~cache_hit ? _GEN_4265 : _GEN_2389; // @[ICache.scala 175:32]
  wire  _GEN_6333 = ~cache_hit ? _GEN_4266 : _GEN_2901; // @[ICache.scala 175:32]
  wire  _GEN_6334 = ~cache_hit ? _GEN_4267 : _GEN_2390; // @[ICache.scala 175:32]
  wire  _GEN_6335 = ~cache_hit ? _GEN_4268 : _GEN_2902; // @[ICache.scala 175:32]
  wire  _GEN_6336 = ~cache_hit ? _GEN_4269 : _GEN_2391; // @[ICache.scala 175:32]
  wire  _GEN_6337 = ~cache_hit ? _GEN_4270 : _GEN_2903; // @[ICache.scala 175:32]
  wire  _GEN_6338 = ~cache_hit ? _GEN_4271 : _GEN_2392; // @[ICache.scala 175:32]
  wire  _GEN_6339 = ~cache_hit ? _GEN_4272 : _GEN_2904; // @[ICache.scala 175:32]
  wire  _GEN_6340 = ~cache_hit ? _GEN_4273 : _GEN_2393; // @[ICache.scala 175:32]
  wire  _GEN_6341 = ~cache_hit ? _GEN_4274 : _GEN_2905; // @[ICache.scala 175:32]
  wire  _GEN_6342 = ~cache_hit ? _GEN_4275 : _GEN_2394; // @[ICache.scala 175:32]
  wire  _GEN_6343 = ~cache_hit ? _GEN_4276 : _GEN_2906; // @[ICache.scala 175:32]
  wire  _GEN_6344 = ~cache_hit ? _GEN_4277 : _GEN_2395; // @[ICache.scala 175:32]
  wire  _GEN_6345 = ~cache_hit ? _GEN_4278 : _GEN_2907; // @[ICache.scala 175:32]
  wire  _GEN_6346 = ~cache_hit ? _GEN_4279 : _GEN_2396; // @[ICache.scala 175:32]
  wire  _GEN_6347 = ~cache_hit ? _GEN_4280 : _GEN_2908; // @[ICache.scala 175:32]
  wire  _GEN_6348 = ~cache_hit ? _GEN_4281 : _GEN_2397; // @[ICache.scala 175:32]
  wire  _GEN_6349 = ~cache_hit ? _GEN_4282 : _GEN_2909; // @[ICache.scala 175:32]
  wire  _GEN_6350 = ~cache_hit ? _GEN_4283 : _GEN_2398; // @[ICache.scala 175:32]
  wire  _GEN_6351 = ~cache_hit ? _GEN_4284 : _GEN_2910; // @[ICache.scala 175:32]
  wire  _GEN_6352 = ~cache_hit ? _GEN_4285 : _GEN_2399; // @[ICache.scala 175:32]
  wire  _GEN_6353 = ~cache_hit ? _GEN_4286 : _GEN_2911; // @[ICache.scala 175:32]
  wire  _GEN_6354 = ~cache_hit ? _GEN_4287 : _GEN_2400; // @[ICache.scala 175:32]
  wire  _GEN_6355 = ~cache_hit ? _GEN_4288 : _GEN_2912; // @[ICache.scala 175:32]
  wire  _GEN_6356 = ~cache_hit ? _GEN_4289 : _GEN_2401; // @[ICache.scala 175:32]
  wire  _GEN_6357 = ~cache_hit ? _GEN_4290 : _GEN_2913; // @[ICache.scala 175:32]
  wire  _GEN_6358 = ~cache_hit ? _GEN_4291 : _GEN_2402; // @[ICache.scala 175:32]
  wire  _GEN_6359 = ~cache_hit ? _GEN_4292 : _GEN_2914; // @[ICache.scala 175:32]
  wire  _GEN_6360 = ~cache_hit ? _GEN_4293 : _GEN_2403; // @[ICache.scala 175:32]
  wire  _GEN_6361 = ~cache_hit ? _GEN_4294 : _GEN_2915; // @[ICache.scala 175:32]
  wire  _GEN_6362 = ~cache_hit ? _GEN_4295 : _GEN_2404; // @[ICache.scala 175:32]
  wire  _GEN_6363 = ~cache_hit ? _GEN_4296 : _GEN_2916; // @[ICache.scala 175:32]
  wire  _GEN_6364 = ~cache_hit ? _GEN_4297 : _GEN_2405; // @[ICache.scala 175:32]
  wire  _GEN_6365 = ~cache_hit ? _GEN_4298 : _GEN_2917; // @[ICache.scala 175:32]
  wire  _GEN_6366 = ~cache_hit ? _GEN_4299 : _GEN_2406; // @[ICache.scala 175:32]
  wire  _GEN_6367 = ~cache_hit ? _GEN_4300 : _GEN_2918; // @[ICache.scala 175:32]
  wire  _GEN_6368 = ~cache_hit ? _GEN_4301 : _GEN_2407; // @[ICache.scala 175:32]
  wire  _GEN_6369 = ~cache_hit ? _GEN_4302 : _GEN_2919; // @[ICache.scala 175:32]
  wire  _GEN_6370 = ~cache_hit ? _GEN_4303 : _GEN_2408; // @[ICache.scala 175:32]
  wire  _GEN_6371 = ~cache_hit ? _GEN_4304 : _GEN_2920; // @[ICache.scala 175:32]
  wire  _GEN_6372 = ~cache_hit ? _GEN_4305 : _GEN_2409; // @[ICache.scala 175:32]
  wire  _GEN_6373 = ~cache_hit ? _GEN_4306 : _GEN_2921; // @[ICache.scala 175:32]
  wire  _GEN_6374 = ~cache_hit ? _GEN_4307 : _GEN_2410; // @[ICache.scala 175:32]
  wire  _GEN_6375 = ~cache_hit ? _GEN_4308 : _GEN_2922; // @[ICache.scala 175:32]
  wire  _GEN_6376 = ~cache_hit ? _GEN_4309 : _GEN_2411; // @[ICache.scala 175:32]
  wire  _GEN_6377 = ~cache_hit ? _GEN_4310 : _GEN_2923; // @[ICache.scala 175:32]
  wire  _GEN_6378 = ~cache_hit ? _GEN_4311 : _GEN_2412; // @[ICache.scala 175:32]
  wire  _GEN_6379 = ~cache_hit ? _GEN_4312 : _GEN_2924; // @[ICache.scala 175:32]
  wire  _GEN_6380 = ~cache_hit ? _GEN_4313 : _GEN_2413; // @[ICache.scala 175:32]
  wire  _GEN_6381 = ~cache_hit ? _GEN_4314 : _GEN_2925; // @[ICache.scala 175:32]
  wire  _GEN_6382 = ~cache_hit ? _GEN_4315 : _GEN_2414; // @[ICache.scala 175:32]
  wire  _GEN_6383 = ~cache_hit ? _GEN_4316 : _GEN_2926; // @[ICache.scala 175:32]
  wire  _GEN_6384 = ~cache_hit ? _GEN_4317 : _GEN_2415; // @[ICache.scala 175:32]
  wire  _GEN_6385 = ~cache_hit ? _GEN_4318 : _GEN_2927; // @[ICache.scala 175:32]
  wire  _GEN_6386 = ~cache_hit ? _GEN_4319 : _GEN_2416; // @[ICache.scala 175:32]
  wire  _GEN_6387 = ~cache_hit ? _GEN_4320 : _GEN_2928; // @[ICache.scala 175:32]
  wire  _GEN_6388 = ~cache_hit ? _GEN_4321 : _GEN_2417; // @[ICache.scala 175:32]
  wire  _GEN_6389 = ~cache_hit ? _GEN_4322 : _GEN_2929; // @[ICache.scala 175:32]
  wire  _GEN_6390 = ~cache_hit ? _GEN_4323 : _GEN_2418; // @[ICache.scala 175:32]
  wire  _GEN_6391 = ~cache_hit ? _GEN_4324 : _GEN_2930; // @[ICache.scala 175:32]
  wire  _GEN_6392 = ~cache_hit ? _GEN_4325 : _GEN_2419; // @[ICache.scala 175:32]
  wire  _GEN_6393 = ~cache_hit ? _GEN_4326 : _GEN_2931; // @[ICache.scala 175:32]
  wire  _GEN_6394 = ~cache_hit ? _GEN_4327 : _GEN_2420; // @[ICache.scala 175:32]
  wire  _GEN_6395 = ~cache_hit ? _GEN_4328 : _GEN_2932; // @[ICache.scala 175:32]
  wire  _GEN_6396 = ~cache_hit ? _GEN_4329 : _GEN_2421; // @[ICache.scala 175:32]
  wire  _GEN_6397 = ~cache_hit ? _GEN_4330 : _GEN_2933; // @[ICache.scala 175:32]
  wire  _GEN_6398 = ~cache_hit ? _GEN_4331 : _GEN_2422; // @[ICache.scala 175:32]
  wire  _GEN_6399 = ~cache_hit ? _GEN_4332 : _GEN_2934; // @[ICache.scala 175:32]
  wire  _GEN_6400 = ~cache_hit ? _GEN_4333 : _GEN_2423; // @[ICache.scala 175:32]
  wire  _GEN_6401 = ~cache_hit ? _GEN_4334 : _GEN_2935; // @[ICache.scala 175:32]
  wire  _GEN_6402 = ~cache_hit ? _GEN_4335 : _GEN_2424; // @[ICache.scala 175:32]
  wire  _GEN_6403 = ~cache_hit ? _GEN_4336 : _GEN_2936; // @[ICache.scala 175:32]
  wire  _GEN_6404 = ~cache_hit ? _GEN_4337 : _GEN_2425; // @[ICache.scala 175:32]
  wire  _GEN_6405 = ~cache_hit ? _GEN_4338 : _GEN_2937; // @[ICache.scala 175:32]
  wire  _GEN_6406 = ~cache_hit ? _GEN_4339 : _GEN_2426; // @[ICache.scala 175:32]
  wire  _GEN_6407 = ~cache_hit ? _GEN_4340 : _GEN_2938; // @[ICache.scala 175:32]
  wire  _GEN_6408 = ~cache_hit ? _GEN_4341 : _GEN_2427; // @[ICache.scala 175:32]
  wire  _GEN_6409 = ~cache_hit ? _GEN_4342 : _GEN_2939; // @[ICache.scala 175:32]
  wire  _GEN_6410 = ~cache_hit ? _GEN_4343 : _GEN_2428; // @[ICache.scala 175:32]
  wire  _GEN_6411 = ~cache_hit ? _GEN_4344 : _GEN_2940; // @[ICache.scala 175:32]
  wire  _GEN_6412 = ~cache_hit ? _GEN_4345 : _GEN_2429; // @[ICache.scala 175:32]
  wire  _GEN_6413 = ~cache_hit ? _GEN_4346 : _GEN_2941; // @[ICache.scala 175:32]
  wire  _GEN_6414 = ~cache_hit ? _GEN_4347 : _GEN_2430; // @[ICache.scala 175:32]
  wire  _GEN_6415 = ~cache_hit ? _GEN_4348 : _GEN_2942; // @[ICache.scala 175:32]
  wire  _GEN_6416 = ~cache_hit ? _GEN_4349 : _GEN_2431; // @[ICache.scala 175:32]
  wire  _GEN_6417 = ~cache_hit ? _GEN_4350 : _GEN_2943; // @[ICache.scala 175:32]
  wire  _GEN_6418 = ~cache_hit ? _GEN_4351 : _GEN_2432; // @[ICache.scala 175:32]
  wire  _GEN_6419 = ~cache_hit ? _GEN_4352 : _GEN_2944; // @[ICache.scala 175:32]
  wire  _GEN_6420 = ~cache_hit ? _GEN_4353 : _GEN_2433; // @[ICache.scala 175:32]
  wire  _GEN_6421 = ~cache_hit ? _GEN_4354 : _GEN_2945; // @[ICache.scala 175:32]
  wire  _GEN_6422 = ~cache_hit ? _GEN_4355 : _GEN_2434; // @[ICache.scala 175:32]
  wire  _GEN_6423 = ~cache_hit ? _GEN_4356 : _GEN_2946; // @[ICache.scala 175:32]
  wire  _GEN_6424 = ~cache_hit ? _GEN_4357 : _GEN_2435; // @[ICache.scala 175:32]
  wire  _GEN_6425 = ~cache_hit ? _GEN_4358 : _GEN_2947; // @[ICache.scala 175:32]
  wire  _GEN_6426 = ~cache_hit ? _GEN_4359 : _GEN_2436; // @[ICache.scala 175:32]
  wire  _GEN_6427 = ~cache_hit ? _GEN_4360 : _GEN_2948; // @[ICache.scala 175:32]
  wire  _GEN_6428 = ~cache_hit ? _GEN_4361 : _GEN_2437; // @[ICache.scala 175:32]
  wire  _GEN_6429 = ~cache_hit ? _GEN_4362 : _GEN_2949; // @[ICache.scala 175:32]
  wire  _GEN_6430 = ~cache_hit ? _GEN_4363 : _GEN_2438; // @[ICache.scala 175:32]
  wire  _GEN_6431 = ~cache_hit ? _GEN_4364 : _GEN_2950; // @[ICache.scala 175:32]
  wire  _GEN_6432 = ~cache_hit ? _GEN_4365 : _GEN_2439; // @[ICache.scala 175:32]
  wire  _GEN_6433 = ~cache_hit ? _GEN_4366 : _GEN_2951; // @[ICache.scala 175:32]
  wire  _GEN_6434 = ~cache_hit ? _GEN_4367 : _GEN_2440; // @[ICache.scala 175:32]
  wire  _GEN_6435 = ~cache_hit ? _GEN_4368 : _GEN_2952; // @[ICache.scala 175:32]
  wire  _GEN_6436 = ~cache_hit ? _GEN_4369 : _GEN_2441; // @[ICache.scala 175:32]
  wire  _GEN_6437 = ~cache_hit ? _GEN_4370 : _GEN_2953; // @[ICache.scala 175:32]
  wire  _GEN_6438 = ~cache_hit ? _GEN_4371 : _GEN_2442; // @[ICache.scala 175:32]
  wire  _GEN_6439 = ~cache_hit ? _GEN_4372 : _GEN_2954; // @[ICache.scala 175:32]
  wire  _GEN_6440 = ~cache_hit ? _GEN_4373 : _GEN_2443; // @[ICache.scala 175:32]
  wire  _GEN_6441 = ~cache_hit ? _GEN_4374 : _GEN_2955; // @[ICache.scala 175:32]
  wire  _GEN_6442 = ~cache_hit ? _GEN_4375 : _GEN_2444; // @[ICache.scala 175:32]
  wire  _GEN_6443 = ~cache_hit ? _GEN_4376 : _GEN_2956; // @[ICache.scala 175:32]
  wire  _GEN_6444 = ~cache_hit ? _GEN_4377 : _GEN_2445; // @[ICache.scala 175:32]
  wire  _GEN_6445 = ~cache_hit ? _GEN_4378 : _GEN_2957; // @[ICache.scala 175:32]
  wire  _GEN_6446 = ~cache_hit ? _GEN_4379 : _GEN_2446; // @[ICache.scala 175:32]
  wire  _GEN_6447 = ~cache_hit ? _GEN_4380 : _GEN_2958; // @[ICache.scala 175:32]
  wire  _GEN_6448 = ~cache_hit ? _GEN_4381 : _GEN_2447; // @[ICache.scala 175:32]
  wire  _GEN_6449 = ~cache_hit ? _GEN_4382 : _GEN_2959; // @[ICache.scala 175:32]
  wire  _GEN_6450 = ~cache_hit ? _GEN_4383 : _GEN_2448; // @[ICache.scala 175:32]
  wire  _GEN_6451 = ~cache_hit ? _GEN_4384 : _GEN_2960; // @[ICache.scala 175:32]
  wire  _GEN_6452 = ~cache_hit ? _GEN_4385 : _GEN_2449; // @[ICache.scala 175:32]
  wire  _GEN_6453 = ~cache_hit ? _GEN_4386 : _GEN_2961; // @[ICache.scala 175:32]
  wire  _GEN_6454 = ~cache_hit ? _GEN_4387 : _GEN_2450; // @[ICache.scala 175:32]
  wire  _GEN_6455 = ~cache_hit ? _GEN_4388 : _GEN_2962; // @[ICache.scala 175:32]
  wire  _GEN_6456 = ~cache_hit ? _GEN_4389 : _GEN_2451; // @[ICache.scala 175:32]
  wire  _GEN_6457 = ~cache_hit ? _GEN_4390 : _GEN_2963; // @[ICache.scala 175:32]
  wire  _GEN_6458 = ~cache_hit ? _GEN_4391 : _GEN_2452; // @[ICache.scala 175:32]
  wire  _GEN_6459 = ~cache_hit ? _GEN_4392 : _GEN_2964; // @[ICache.scala 175:32]
  wire  _GEN_6460 = ~cache_hit ? _GEN_4393 : _GEN_2453; // @[ICache.scala 175:32]
  wire  _GEN_6461 = ~cache_hit ? _GEN_4394 : _GEN_2965; // @[ICache.scala 175:32]
  wire  _GEN_6462 = ~cache_hit ? _GEN_4395 : _GEN_2454; // @[ICache.scala 175:32]
  wire  _GEN_6463 = ~cache_hit ? _GEN_4396 : _GEN_2966; // @[ICache.scala 175:32]
  wire  _GEN_6464 = ~cache_hit ? _GEN_4397 : _GEN_2455; // @[ICache.scala 175:32]
  wire  _GEN_6465 = ~cache_hit ? _GEN_4398 : _GEN_2967; // @[ICache.scala 175:32]
  wire  _GEN_6466 = ~cache_hit ? _GEN_4399 : _GEN_2456; // @[ICache.scala 175:32]
  wire  _GEN_6467 = ~cache_hit ? _GEN_4400 : _GEN_2968; // @[ICache.scala 175:32]
  wire  _GEN_6468 = ~cache_hit ? _GEN_4401 : _GEN_2457; // @[ICache.scala 175:32]
  wire  _GEN_6469 = ~cache_hit ? _GEN_4402 : _GEN_2969; // @[ICache.scala 175:32]
  wire  _GEN_6470 = ~cache_hit ? _GEN_4403 : _GEN_2458; // @[ICache.scala 175:32]
  wire  _GEN_6471 = ~cache_hit ? _GEN_4404 : _GEN_2970; // @[ICache.scala 175:32]
  wire  _GEN_6472 = ~cache_hit ? _GEN_4405 : _GEN_2459; // @[ICache.scala 175:32]
  wire  _GEN_6473 = ~cache_hit ? _GEN_4406 : _GEN_2971; // @[ICache.scala 175:32]
  wire  _GEN_6474 = ~cache_hit ? _GEN_4407 : _GEN_2460; // @[ICache.scala 175:32]
  wire  _GEN_6475 = ~cache_hit ? _GEN_4408 : _GEN_2972; // @[ICache.scala 175:32]
  wire  _GEN_6476 = ~cache_hit ? _GEN_4409 : _GEN_2461; // @[ICache.scala 175:32]
  wire  _GEN_6477 = ~cache_hit ? _GEN_4410 : _GEN_2973; // @[ICache.scala 175:32]
  wire  _GEN_6478 = ~cache_hit ? _GEN_4411 : _GEN_2462; // @[ICache.scala 175:32]
  wire  _GEN_6479 = ~cache_hit ? _GEN_4412 : _GEN_2974; // @[ICache.scala 175:32]
  wire  _GEN_6480 = ~cache_hit ? _GEN_4413 : _GEN_2463; // @[ICache.scala 175:32]
  wire  _GEN_6481 = ~cache_hit ? _GEN_4414 : _GEN_2975; // @[ICache.scala 175:32]
  wire  _GEN_6482 = ~cache_hit ? _GEN_4415 : _GEN_2464; // @[ICache.scala 175:32]
  wire  _GEN_6483 = ~cache_hit ? _GEN_4416 : _GEN_2976; // @[ICache.scala 175:32]
  wire  _GEN_6484 = ~cache_hit ? _GEN_4417 : _GEN_2465; // @[ICache.scala 175:32]
  wire  _GEN_6485 = ~cache_hit ? _GEN_4418 : _GEN_2977; // @[ICache.scala 175:32]
  wire  _GEN_6486 = ~cache_hit ? _GEN_4419 : _GEN_2466; // @[ICache.scala 175:32]
  wire  _GEN_6487 = ~cache_hit ? _GEN_4420 : _GEN_2978; // @[ICache.scala 175:32]
  wire  _GEN_6488 = ~cache_hit ? _GEN_4421 : _GEN_2467; // @[ICache.scala 175:32]
  wire  _GEN_6489 = ~cache_hit ? _GEN_4422 : _GEN_2979; // @[ICache.scala 175:32]
  wire  _GEN_6490 = ~cache_hit ? _GEN_4423 : _GEN_2468; // @[ICache.scala 175:32]
  wire  _GEN_6491 = ~cache_hit ? _GEN_4424 : _GEN_2980; // @[ICache.scala 175:32]
  wire  _GEN_6492 = ~cache_hit ? _GEN_4425 : _GEN_2469; // @[ICache.scala 175:32]
  wire  _GEN_6493 = ~cache_hit ? _GEN_4426 : _GEN_2981; // @[ICache.scala 175:32]
  wire  _GEN_6494 = ~cache_hit ? _GEN_4427 : _GEN_2470; // @[ICache.scala 175:32]
  wire  _GEN_6495 = ~cache_hit ? _GEN_4428 : _GEN_2982; // @[ICache.scala 175:32]
  wire  _GEN_6496 = ~cache_hit ? _GEN_4429 : _GEN_2471; // @[ICache.scala 175:32]
  wire  _GEN_6497 = ~cache_hit ? _GEN_4430 : _GEN_2983; // @[ICache.scala 175:32]
  wire  _GEN_6498 = ~cache_hit ? _GEN_4431 : _GEN_2472; // @[ICache.scala 175:32]
  wire  _GEN_6499 = ~cache_hit ? _GEN_4432 : _GEN_2984; // @[ICache.scala 175:32]
  wire  _GEN_6500 = ~cache_hit ? _GEN_4433 : _GEN_2473; // @[ICache.scala 175:32]
  wire  _GEN_6501 = ~cache_hit ? _GEN_4434 : _GEN_2985; // @[ICache.scala 175:32]
  wire  _GEN_6502 = ~cache_hit ? _GEN_4435 : _GEN_2474; // @[ICache.scala 175:32]
  wire  _GEN_6503 = ~cache_hit ? _GEN_4436 : _GEN_2986; // @[ICache.scala 175:32]
  wire  _GEN_6504 = ~cache_hit ? _GEN_4437 : _GEN_2475; // @[ICache.scala 175:32]
  wire  _GEN_6505 = ~cache_hit ? _GEN_4438 : _GEN_2987; // @[ICache.scala 175:32]
  wire  _GEN_6506 = ~cache_hit ? _GEN_4439 : _GEN_2476; // @[ICache.scala 175:32]
  wire  _GEN_6507 = ~cache_hit ? _GEN_4440 : _GEN_2988; // @[ICache.scala 175:32]
  wire  _GEN_6508 = ~cache_hit ? _GEN_4441 : _GEN_2477; // @[ICache.scala 175:32]
  wire  _GEN_6509 = ~cache_hit ? _GEN_4442 : _GEN_2989; // @[ICache.scala 175:32]
  wire  _GEN_6510 = ~cache_hit ? _GEN_4443 : _GEN_2478; // @[ICache.scala 175:32]
  wire  _GEN_6511 = ~cache_hit ? _GEN_4444 : _GEN_2990; // @[ICache.scala 175:32]
  wire  _GEN_6512 = ~cache_hit ? _GEN_4445 : _GEN_2479; // @[ICache.scala 175:32]
  wire  _GEN_6513 = ~cache_hit ? _GEN_4446 : _GEN_2991; // @[ICache.scala 175:32]
  wire  _GEN_6514 = ~cache_hit ? _GEN_4447 : _GEN_2480; // @[ICache.scala 175:32]
  wire  _GEN_6515 = ~cache_hit ? _GEN_4448 : _GEN_2992; // @[ICache.scala 175:32]
  wire  _GEN_6516 = ~cache_hit ? _GEN_4449 : _GEN_2481; // @[ICache.scala 175:32]
  wire  _GEN_6517 = ~cache_hit ? _GEN_4450 : _GEN_2993; // @[ICache.scala 175:32]
  wire  _GEN_6518 = ~cache_hit ? _GEN_4451 : _GEN_2482; // @[ICache.scala 175:32]
  wire  _GEN_6519 = ~cache_hit ? _GEN_4452 : _GEN_2994; // @[ICache.scala 175:32]
  wire  _GEN_6520 = ~cache_hit ? _GEN_4453 : _GEN_2483; // @[ICache.scala 175:32]
  wire  _GEN_6521 = ~cache_hit ? _GEN_4454 : _GEN_2995; // @[ICache.scala 175:32]
  wire  _GEN_6522 = ~cache_hit ? _GEN_4455 : _GEN_2484; // @[ICache.scala 175:32]
  wire  _GEN_6523 = ~cache_hit ? _GEN_4456 : _GEN_2996; // @[ICache.scala 175:32]
  wire  _GEN_6524 = ~cache_hit ? _GEN_4457 : _GEN_2485; // @[ICache.scala 175:32]
  wire  _GEN_6525 = ~cache_hit ? _GEN_4458 : _GEN_2997; // @[ICache.scala 175:32]
  wire  _GEN_6526 = ~cache_hit ? _GEN_4459 : _GEN_2486; // @[ICache.scala 175:32]
  wire  _GEN_6527 = ~cache_hit ? _GEN_4460 : _GEN_2998; // @[ICache.scala 175:32]
  wire  _GEN_6528 = ~cache_hit ? _GEN_4461 : _GEN_2487; // @[ICache.scala 175:32]
  wire  _GEN_6529 = ~cache_hit ? _GEN_4462 : _GEN_2999; // @[ICache.scala 175:32]
  wire  _GEN_6530 = ~cache_hit ? _GEN_4463 : _GEN_2488; // @[ICache.scala 175:32]
  wire  _GEN_6531 = ~cache_hit ? _GEN_4464 : _GEN_3000; // @[ICache.scala 175:32]
  wire  _GEN_6532 = ~cache_hit ? _GEN_4465 : _GEN_2489; // @[ICache.scala 175:32]
  wire  _GEN_6533 = ~cache_hit ? _GEN_4466 : _GEN_3001; // @[ICache.scala 175:32]
  wire  _GEN_6534 = ~cache_hit ? _GEN_4467 : _GEN_2490; // @[ICache.scala 175:32]
  wire  _GEN_6535 = ~cache_hit ? _GEN_4468 : _GEN_3002; // @[ICache.scala 175:32]
  wire  _GEN_6536 = ~cache_hit ? _GEN_4469 : _GEN_2491; // @[ICache.scala 175:32]
  wire  _GEN_6537 = ~cache_hit ? _GEN_4470 : _GEN_3003; // @[ICache.scala 175:32]
  wire  _GEN_6538 = ~cache_hit ? _GEN_4471 : _GEN_2492; // @[ICache.scala 175:32]
  wire  _GEN_6539 = ~cache_hit ? _GEN_4472 : _GEN_3004; // @[ICache.scala 175:32]
  wire  _GEN_6540 = ~cache_hit ? _GEN_4473 : _GEN_2493; // @[ICache.scala 175:32]
  wire  _GEN_6541 = ~cache_hit ? _GEN_4474 : _GEN_3005; // @[ICache.scala 175:32]
  wire  _GEN_6542 = ~cache_hit ? _GEN_4475 : _GEN_2494; // @[ICache.scala 175:32]
  wire  _GEN_6543 = ~cache_hit ? _GEN_4476 : _GEN_3006; // @[ICache.scala 175:32]
  wire  _GEN_6544 = ~cache_hit ? _GEN_4477 : _GEN_2495; // @[ICache.scala 175:32]
  wire  _GEN_6545 = ~cache_hit ? _GEN_4478 : _GEN_3007; // @[ICache.scala 175:32]
  wire  _GEN_6546 = ~cache_hit ? _GEN_4479 : _GEN_2496; // @[ICache.scala 175:32]
  wire  _GEN_6547 = ~cache_hit ? _GEN_4480 : _GEN_3008; // @[ICache.scala 175:32]
  wire  _GEN_6548 = ~cache_hit ? _GEN_4481 : _GEN_2497; // @[ICache.scala 175:32]
  wire  _GEN_6549 = ~cache_hit ? _GEN_4482 : _GEN_3009; // @[ICache.scala 175:32]
  wire  _GEN_6550 = ~cache_hit ? _GEN_4483 : _GEN_2498; // @[ICache.scala 175:32]
  wire  _GEN_6551 = ~cache_hit ? _GEN_4484 : _GEN_3010; // @[ICache.scala 175:32]
  wire  _GEN_6552 = ~cache_hit ? _GEN_4485 : _GEN_2499; // @[ICache.scala 175:32]
  wire  _GEN_6553 = ~cache_hit ? _GEN_4486 : _GEN_3011; // @[ICache.scala 175:32]
  wire  _GEN_6554 = ~cache_hit ? _GEN_4487 : _GEN_2500; // @[ICache.scala 175:32]
  wire  _GEN_6555 = ~cache_hit ? _GEN_4488 : _GEN_3012; // @[ICache.scala 175:32]
  wire  _GEN_6556 = ~cache_hit ? _GEN_4489 : _GEN_2501; // @[ICache.scala 175:32]
  wire  _GEN_6557 = ~cache_hit ? _GEN_4490 : _GEN_3013; // @[ICache.scala 175:32]
  wire  _GEN_6558 = ~cache_hit ? _GEN_4491 : _GEN_2502; // @[ICache.scala 175:32]
  wire  _GEN_6559 = ~cache_hit ? _GEN_4492 : _GEN_3014; // @[ICache.scala 175:32]
  wire  _GEN_6560 = ~cache_hit ? _GEN_4493 : _GEN_2503; // @[ICache.scala 175:32]
  wire  _GEN_6561 = ~cache_hit ? _GEN_4494 : _GEN_3015; // @[ICache.scala 175:32]
  wire  _GEN_6562 = ~cache_hit ? _GEN_4495 : _GEN_2504; // @[ICache.scala 175:32]
  wire  _GEN_6563 = ~cache_hit ? _GEN_4496 : _GEN_3016; // @[ICache.scala 175:32]
  wire  _GEN_6564 = ~cache_hit ? _GEN_4497 : _GEN_2505; // @[ICache.scala 175:32]
  wire  _GEN_6565 = ~cache_hit ? _GEN_4498 : _GEN_3017; // @[ICache.scala 175:32]
  wire  _GEN_6566 = ~cache_hit ? _GEN_4499 : _GEN_2506; // @[ICache.scala 175:32]
  wire  _GEN_6567 = ~cache_hit ? _GEN_4500 : _GEN_3018; // @[ICache.scala 175:32]
  wire  _GEN_6568 = ~cache_hit ? _GEN_4501 : _GEN_2507; // @[ICache.scala 175:32]
  wire  _GEN_6569 = ~cache_hit ? _GEN_4502 : _GEN_3019; // @[ICache.scala 175:32]
  wire  _GEN_6570 = ~cache_hit ? _GEN_4503 : _GEN_2508; // @[ICache.scala 175:32]
  wire  _GEN_6571 = ~cache_hit ? _GEN_4504 : _GEN_3020; // @[ICache.scala 175:32]
  wire  _GEN_6572 = ~cache_hit ? _GEN_4505 : _GEN_2509; // @[ICache.scala 175:32]
  wire  _GEN_6573 = ~cache_hit ? _GEN_4506 : _GEN_3021; // @[ICache.scala 175:32]
  wire  _GEN_6574 = ~cache_hit ? _GEN_4507 : _GEN_2510; // @[ICache.scala 175:32]
  wire  _GEN_6575 = ~cache_hit ? _GEN_4508 : _GEN_3022; // @[ICache.scala 175:32]
  wire  _GEN_6576 = ~cache_hit ? _GEN_4509 : _GEN_2511; // @[ICache.scala 175:32]
  wire  _GEN_6577 = ~cache_hit ? _GEN_4510 : _GEN_3023; // @[ICache.scala 175:32]
  wire  _GEN_6578 = ~cache_hit ? _GEN_4511 : _GEN_2512; // @[ICache.scala 175:32]
  wire  _GEN_6579 = ~cache_hit ? _GEN_4512 : _GEN_3024; // @[ICache.scala 175:32]
  wire  _GEN_6580 = ~cache_hit ? _GEN_4513 : _GEN_2513; // @[ICache.scala 175:32]
  wire  _GEN_6581 = ~cache_hit ? _GEN_4514 : _GEN_3025; // @[ICache.scala 175:32]
  wire  _GEN_6582 = ~cache_hit ? _GEN_4515 : _GEN_2514; // @[ICache.scala 175:32]
  wire  _GEN_6583 = ~cache_hit ? _GEN_4516 : _GEN_3026; // @[ICache.scala 175:32]
  wire  _GEN_6584 = ~cache_hit ? _GEN_4517 : _GEN_2515; // @[ICache.scala 175:32]
  wire  _GEN_6585 = ~cache_hit ? _GEN_4518 : _GEN_3027; // @[ICache.scala 175:32]
  wire  _GEN_6586 = ~cache_hit ? _GEN_4519 : _GEN_2516; // @[ICache.scala 175:32]
  wire  _GEN_6587 = ~cache_hit ? _GEN_4520 : _GEN_3028; // @[ICache.scala 175:32]
  wire  _GEN_6588 = ~cache_hit ? _GEN_4521 : _GEN_2517; // @[ICache.scala 175:32]
  wire  _GEN_6589 = ~cache_hit ? _GEN_4522 : _GEN_3029; // @[ICache.scala 175:32]
  wire  _GEN_6590 = ~cache_hit ? _GEN_4523 : _GEN_2518; // @[ICache.scala 175:32]
  wire  _GEN_6591 = ~cache_hit ? _GEN_4524 : _GEN_3030; // @[ICache.scala 175:32]
  wire  _GEN_6592 = ~cache_hit ? _GEN_4525 : _GEN_2519; // @[ICache.scala 175:32]
  wire  _GEN_6593 = ~cache_hit ? _GEN_4526 : _GEN_3031; // @[ICache.scala 175:32]
  wire  _GEN_6594 = ~cache_hit ? _GEN_4527 : _GEN_2520; // @[ICache.scala 175:32]
  wire  _GEN_6595 = ~cache_hit ? _GEN_4528 : _GEN_3032; // @[ICache.scala 175:32]
  wire  _GEN_6596 = ~cache_hit ? _GEN_4529 : _GEN_2521; // @[ICache.scala 175:32]
  wire  _GEN_6597 = ~cache_hit ? _GEN_4530 : _GEN_3033; // @[ICache.scala 175:32]
  wire  _GEN_6598 = ~cache_hit ? _GEN_4531 : _GEN_2522; // @[ICache.scala 175:32]
  wire  _GEN_6599 = ~cache_hit ? _GEN_4532 : _GEN_3034; // @[ICache.scala 175:32]
  wire  _GEN_6600 = ~cache_hit ? _GEN_4533 : _GEN_2523; // @[ICache.scala 175:32]
  wire  _GEN_6601 = ~cache_hit ? _GEN_4534 : _GEN_3035; // @[ICache.scala 175:32]
  wire  _GEN_6602 = ~cache_hit ? _GEN_4535 : _GEN_2524; // @[ICache.scala 175:32]
  wire  _GEN_6603 = ~cache_hit ? _GEN_4536 : _GEN_3036; // @[ICache.scala 175:32]
  wire  _GEN_6604 = ~cache_hit ? _GEN_4537 : _GEN_2525; // @[ICache.scala 175:32]
  wire  _GEN_6605 = ~cache_hit ? _GEN_4538 : _GEN_3037; // @[ICache.scala 175:32]
  wire  _GEN_6606 = ~cache_hit ? _GEN_4539 : _GEN_2526; // @[ICache.scala 175:32]
  wire  _GEN_6607 = ~cache_hit ? _GEN_4540 : _GEN_3038; // @[ICache.scala 175:32]
  wire  _GEN_6608 = ~cache_hit ? _GEN_4541 : _GEN_2527; // @[ICache.scala 175:32]
  wire  _GEN_6609 = ~cache_hit ? _GEN_4542 : _GEN_3039; // @[ICache.scala 175:32]
  wire  _GEN_6610 = ~cache_hit ? _GEN_4543 : _GEN_2528; // @[ICache.scala 175:32]
  wire  _GEN_6611 = ~cache_hit ? _GEN_4544 : _GEN_3040; // @[ICache.scala 175:32]
  wire  _GEN_6612 = ~cache_hit ? _GEN_4545 : _GEN_2529; // @[ICache.scala 175:32]
  wire  _GEN_6613 = ~cache_hit ? _GEN_4546 : _GEN_3041; // @[ICache.scala 175:32]
  wire  _GEN_6614 = ~cache_hit ? _GEN_4547 : _GEN_2530; // @[ICache.scala 175:32]
  wire  _GEN_6615 = ~cache_hit ? _GEN_4548 : _GEN_3042; // @[ICache.scala 175:32]
  wire  _GEN_6616 = ~cache_hit ? _GEN_4549 : _GEN_2531; // @[ICache.scala 175:32]
  wire  _GEN_6617 = ~cache_hit ? _GEN_4550 : _GEN_3043; // @[ICache.scala 175:32]
  wire  _GEN_6618 = ~cache_hit ? _GEN_4551 : _GEN_2532; // @[ICache.scala 175:32]
  wire  _GEN_6619 = ~cache_hit ? _GEN_4552 : _GEN_3044; // @[ICache.scala 175:32]
  wire  _GEN_6620 = ~cache_hit ? _GEN_4553 : _GEN_2533; // @[ICache.scala 175:32]
  wire  _GEN_6621 = ~cache_hit ? _GEN_4554 : _GEN_3045; // @[ICache.scala 175:32]
  wire  _GEN_6622 = ~cache_hit ? _GEN_4555 : _GEN_2534; // @[ICache.scala 175:32]
  wire  _GEN_6623 = ~cache_hit ? _GEN_4556 : _GEN_3046; // @[ICache.scala 175:32]
  wire  _GEN_6624 = ~cache_hit ? _GEN_4557 : _GEN_2535; // @[ICache.scala 175:32]
  wire  _GEN_6625 = ~cache_hit ? _GEN_4558 : _GEN_3047; // @[ICache.scala 175:32]
  wire  _GEN_6626 = ~cache_hit ? _GEN_4559 : _GEN_2536; // @[ICache.scala 175:32]
  wire  _GEN_6627 = ~cache_hit ? _GEN_4560 : _GEN_3048; // @[ICache.scala 175:32]
  wire  _GEN_6628 = ~cache_hit ? _GEN_4561 : _GEN_2537; // @[ICache.scala 175:32]
  wire  _GEN_6629 = ~cache_hit ? _GEN_4562 : _GEN_3049; // @[ICache.scala 175:32]
  wire  _GEN_6630 = ~cache_hit ? _GEN_4563 : _GEN_2538; // @[ICache.scala 175:32]
  wire  _GEN_6631 = ~cache_hit ? _GEN_4564 : _GEN_3050; // @[ICache.scala 175:32]
  wire  _GEN_6632 = ~cache_hit ? _GEN_4565 : _GEN_2539; // @[ICache.scala 175:32]
  wire  _GEN_6633 = ~cache_hit ? _GEN_4566 : _GEN_3051; // @[ICache.scala 175:32]
  wire  _GEN_6634 = ~cache_hit ? _GEN_4567 : _GEN_2540; // @[ICache.scala 175:32]
  wire  _GEN_6635 = ~cache_hit ? _GEN_4568 : _GEN_3052; // @[ICache.scala 175:32]
  wire  _GEN_6636 = ~cache_hit ? _GEN_4569 : _GEN_2541; // @[ICache.scala 175:32]
  wire  _GEN_6637 = ~cache_hit ? _GEN_4570 : _GEN_3053; // @[ICache.scala 175:32]
  wire  _GEN_6638 = ~cache_hit ? _GEN_4571 : _GEN_2542; // @[ICache.scala 175:32]
  wire  _GEN_6639 = ~cache_hit ? _GEN_4572 : _GEN_3054; // @[ICache.scala 175:32]
  wire  _GEN_6640 = ~cache_hit ? _GEN_4573 : _GEN_2543; // @[ICache.scala 175:32]
  wire  _GEN_6641 = ~cache_hit ? _GEN_4574 : _GEN_3055; // @[ICache.scala 175:32]
  wire  _GEN_6642 = ~cache_hit ? _GEN_4575 : _GEN_2544; // @[ICache.scala 175:32]
  wire  _GEN_6643 = ~cache_hit ? _GEN_4576 : _GEN_3056; // @[ICache.scala 175:32]
  wire  _GEN_6644 = ~cache_hit ? _GEN_4577 : _GEN_2545; // @[ICache.scala 175:32]
  wire  _GEN_6645 = ~cache_hit ? _GEN_4578 : _GEN_3057; // @[ICache.scala 175:32]
  wire  _GEN_6646 = ~cache_hit ? _GEN_4579 : _GEN_2546; // @[ICache.scala 175:32]
  wire  _GEN_6647 = ~cache_hit ? _GEN_4580 : _GEN_3058; // @[ICache.scala 175:32]
  wire  _GEN_6648 = ~cache_hit ? _GEN_4581 : _GEN_2547; // @[ICache.scala 175:32]
  wire  _GEN_6649 = ~cache_hit ? _GEN_4582 : _GEN_3059; // @[ICache.scala 175:32]
  wire  _GEN_6650 = ~cache_hit ? _GEN_4583 : _GEN_2548; // @[ICache.scala 175:32]
  wire  _GEN_6651 = ~cache_hit ? _GEN_4584 : _GEN_3060; // @[ICache.scala 175:32]
  wire  _GEN_6652 = ~cache_hit ? _GEN_4585 : _GEN_2549; // @[ICache.scala 175:32]
  wire  _GEN_6653 = ~cache_hit ? _GEN_4586 : _GEN_3061; // @[ICache.scala 175:32]
  wire  _GEN_6654 = ~cache_hit ? _GEN_4587 : _GEN_2550; // @[ICache.scala 175:32]
  wire  _GEN_6655 = ~cache_hit ? _GEN_4588 : _GEN_3062; // @[ICache.scala 175:32]
  wire  _GEN_6656 = ~cache_hit ? _GEN_4589 : _GEN_2551; // @[ICache.scala 175:32]
  wire  _GEN_6657 = ~cache_hit ? _GEN_4590 : _GEN_3063; // @[ICache.scala 175:32]
  wire  _GEN_6658 = ~cache_hit ? _GEN_4591 : _GEN_2552; // @[ICache.scala 175:32]
  wire  _GEN_6659 = ~cache_hit ? _GEN_4592 : _GEN_3064; // @[ICache.scala 175:32]
  wire  _GEN_6660 = ~cache_hit ? _GEN_4593 : _GEN_2553; // @[ICache.scala 175:32]
  wire  _GEN_6661 = ~cache_hit ? _GEN_4594 : _GEN_3065; // @[ICache.scala 175:32]
  wire  _GEN_6662 = ~cache_hit ? _GEN_4595 : _GEN_2554; // @[ICache.scala 175:32]
  wire  _GEN_6663 = ~cache_hit ? _GEN_4596 : _GEN_3066; // @[ICache.scala 175:32]
  wire  _GEN_6664 = ~cache_hit ? _GEN_4597 : _GEN_2555; // @[ICache.scala 175:32]
  wire  _GEN_6665 = ~cache_hit ? _GEN_4598 : _GEN_3067; // @[ICache.scala 175:32]
  wire  _GEN_6666 = ~cache_hit ? _GEN_4599 : _GEN_2556; // @[ICache.scala 175:32]
  wire  _GEN_6667 = ~cache_hit ? _GEN_4600 : _GEN_3068; // @[ICache.scala 175:32]
  wire  _GEN_6668 = ~cache_hit ? _GEN_4601 : _GEN_2557; // @[ICache.scala 175:32]
  wire  _GEN_6669 = ~cache_hit ? _GEN_4602 : _GEN_3069; // @[ICache.scala 175:32]
  wire  _GEN_6670 = ~cache_hit ? _GEN_4603 : _GEN_2558; // @[ICache.scala 175:32]
  wire  _GEN_6671 = ~cache_hit ? _GEN_4604 : _GEN_3070; // @[ICache.scala 175:32]
  wire  _GEN_6672 = ~cache_hit ? _GEN_4605 : _GEN_2559; // @[ICache.scala 175:32]
  wire  _GEN_6673 = ~cache_hit ? _GEN_4606 : _GEN_3071; // @[ICache.scala 175:32]
  wire  _GEN_6674 = ~cache_hit ? _GEN_4607 : _GEN_2560; // @[ICache.scala 175:32]
  wire  _GEN_6675 = ~cache_hit ? _GEN_4608 : _GEN_3072; // @[ICache.scala 175:32]
  wire  _GEN_6676 = ~cache_hit ? _GEN_4609 : _GEN_2561; // @[ICache.scala 175:32]
  wire  _GEN_6677 = ~cache_hit ? _GEN_4610 : _GEN_3073; // @[ICache.scala 175:32]
  wire  _GEN_6678 = ~cache_hit ? _GEN_4611 : _GEN_2562; // @[ICache.scala 175:32]
  wire  _GEN_6679 = ~cache_hit ? _GEN_4612 : _GEN_3074; // @[ICache.scala 175:32]
  wire  _GEN_6680 = ~cache_hit ? _GEN_4613 : _GEN_2563; // @[ICache.scala 175:32]
  wire  _GEN_6681 = ~cache_hit ? _GEN_4614 : _GEN_3075; // @[ICache.scala 175:32]
  wire  _GEN_6682 = ~cache_hit ? _GEN_4615 : _GEN_2564; // @[ICache.scala 175:32]
  wire  _GEN_6683 = ~cache_hit ? _GEN_4616 : _GEN_3076; // @[ICache.scala 175:32]
  wire [4:0] _GEN_6684 = ~cache_hit ? 5'h0 : axi_cnt; // @[ICache.scala 109:24 175:32 187:60]
  wire  _GEN_6685 = ~cache_hit ? meta_0_lru : _GEN_5133; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6686 = ~cache_hit ? meta_1_lru : _GEN_5134; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6687 = ~cache_hit ? meta_2_lru : _GEN_5135; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6688 = ~cache_hit ? meta_3_lru : _GEN_5136; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6689 = ~cache_hit ? meta_4_lru : _GEN_5137; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6690 = ~cache_hit ? meta_5_lru : _GEN_5138; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6691 = ~cache_hit ? meta_6_lru : _GEN_5139; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6692 = ~cache_hit ? meta_7_lru : _GEN_5140; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6693 = ~cache_hit ? meta_8_lru : _GEN_5141; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6694 = ~cache_hit ? meta_9_lru : _GEN_5142; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6695 = ~cache_hit ? meta_10_lru : _GEN_5143; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6696 = ~cache_hit ? meta_11_lru : _GEN_5144; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6697 = ~cache_hit ? meta_12_lru : _GEN_5145; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6698 = ~cache_hit ? meta_13_lru : _GEN_5146; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6699 = ~cache_hit ? meta_14_lru : _GEN_5147; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6700 = ~cache_hit ? meta_15_lru : _GEN_5148; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6701 = ~cache_hit ? meta_16_lru : _GEN_5149; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6702 = ~cache_hit ? meta_17_lru : _GEN_5150; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6703 = ~cache_hit ? meta_18_lru : _GEN_5151; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6704 = ~cache_hit ? meta_19_lru : _GEN_5152; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6705 = ~cache_hit ? meta_20_lru : _GEN_5153; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6706 = ~cache_hit ? meta_21_lru : _GEN_5154; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6707 = ~cache_hit ? meta_22_lru : _GEN_5155; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6708 = ~cache_hit ? meta_23_lru : _GEN_5156; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6709 = ~cache_hit ? meta_24_lru : _GEN_5157; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6710 = ~cache_hit ? meta_25_lru : _GEN_5158; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6711 = ~cache_hit ? meta_26_lru : _GEN_5159; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6712 = ~cache_hit ? meta_27_lru : _GEN_5160; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6713 = ~cache_hit ? meta_28_lru : _GEN_5161; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6714 = ~cache_hit ? meta_29_lru : _GEN_5162; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6715 = ~cache_hit ? meta_30_lru : _GEN_5163; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6716 = ~cache_hit ? meta_31_lru : _GEN_5164; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6717 = ~cache_hit ? meta_32_lru : _GEN_5165; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6718 = ~cache_hit ? meta_33_lru : _GEN_5166; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6719 = ~cache_hit ? meta_34_lru : _GEN_5167; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6720 = ~cache_hit ? meta_35_lru : _GEN_5168; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6721 = ~cache_hit ? meta_36_lru : _GEN_5169; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6722 = ~cache_hit ? meta_37_lru : _GEN_5170; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6723 = ~cache_hit ? meta_38_lru : _GEN_5171; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6724 = ~cache_hit ? meta_39_lru : _GEN_5172; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6725 = ~cache_hit ? meta_40_lru : _GEN_5173; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6726 = ~cache_hit ? meta_41_lru : _GEN_5174; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6727 = ~cache_hit ? meta_42_lru : _GEN_5175; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6728 = ~cache_hit ? meta_43_lru : _GEN_5176; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6729 = ~cache_hit ? meta_44_lru : _GEN_5177; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6730 = ~cache_hit ? meta_45_lru : _GEN_5178; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6731 = ~cache_hit ? meta_46_lru : _GEN_5179; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6732 = ~cache_hit ? meta_47_lru : _GEN_5180; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6733 = ~cache_hit ? meta_48_lru : _GEN_5181; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6734 = ~cache_hit ? meta_49_lru : _GEN_5182; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6735 = ~cache_hit ? meta_50_lru : _GEN_5183; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6736 = ~cache_hit ? meta_51_lru : _GEN_5184; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6737 = ~cache_hit ? meta_52_lru : _GEN_5185; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6738 = ~cache_hit ? meta_53_lru : _GEN_5186; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6739 = ~cache_hit ? meta_54_lru : _GEN_5187; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6740 = ~cache_hit ? meta_55_lru : _GEN_5188; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6741 = ~cache_hit ? meta_56_lru : _GEN_5189; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6742 = ~cache_hit ? meta_57_lru : _GEN_5190; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6743 = ~cache_hit ? meta_58_lru : _GEN_5191; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6744 = ~cache_hit ? meta_59_lru : _GEN_5192; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6745 = ~cache_hit ? meta_60_lru : _GEN_5193; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6746 = ~cache_hit ? meta_61_lru : _GEN_5194; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6747 = ~cache_hit ? meta_62_lru : _GEN_5195; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6748 = ~cache_hit ? meta_63_lru : _GEN_5196; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6749 = ~cache_hit ? meta_64_lru : _GEN_5197; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6750 = ~cache_hit ? meta_65_lru : _GEN_5198; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6751 = ~cache_hit ? meta_66_lru : _GEN_5199; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6752 = ~cache_hit ? meta_67_lru : _GEN_5200; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6753 = ~cache_hit ? meta_68_lru : _GEN_5201; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6754 = ~cache_hit ? meta_69_lru : _GEN_5202; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6755 = ~cache_hit ? meta_70_lru : _GEN_5203; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6756 = ~cache_hit ? meta_71_lru : _GEN_5204; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6757 = ~cache_hit ? meta_72_lru : _GEN_5205; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6758 = ~cache_hit ? meta_73_lru : _GEN_5206; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6759 = ~cache_hit ? meta_74_lru : _GEN_5207; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6760 = ~cache_hit ? meta_75_lru : _GEN_5208; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6761 = ~cache_hit ? meta_76_lru : _GEN_5209; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6762 = ~cache_hit ? meta_77_lru : _GEN_5210; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6763 = ~cache_hit ? meta_78_lru : _GEN_5211; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6764 = ~cache_hit ? meta_79_lru : _GEN_5212; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6765 = ~cache_hit ? meta_80_lru : _GEN_5213; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6766 = ~cache_hit ? meta_81_lru : _GEN_5214; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6767 = ~cache_hit ? meta_82_lru : _GEN_5215; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6768 = ~cache_hit ? meta_83_lru : _GEN_5216; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6769 = ~cache_hit ? meta_84_lru : _GEN_5217; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6770 = ~cache_hit ? meta_85_lru : _GEN_5218; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6771 = ~cache_hit ? meta_86_lru : _GEN_5219; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6772 = ~cache_hit ? meta_87_lru : _GEN_5220; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6773 = ~cache_hit ? meta_88_lru : _GEN_5221; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6774 = ~cache_hit ? meta_89_lru : _GEN_5222; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6775 = ~cache_hit ? meta_90_lru : _GEN_5223; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6776 = ~cache_hit ? meta_91_lru : _GEN_5224; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6777 = ~cache_hit ? meta_92_lru : _GEN_5225; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6778 = ~cache_hit ? meta_93_lru : _GEN_5226; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6779 = ~cache_hit ? meta_94_lru : _GEN_5227; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6780 = ~cache_hit ? meta_95_lru : _GEN_5228; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6781 = ~cache_hit ? meta_96_lru : _GEN_5229; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6782 = ~cache_hit ? meta_97_lru : _GEN_5230; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6783 = ~cache_hit ? meta_98_lru : _GEN_5231; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6784 = ~cache_hit ? meta_99_lru : _GEN_5232; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6785 = ~cache_hit ? meta_100_lru : _GEN_5233; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6786 = ~cache_hit ? meta_101_lru : _GEN_5234; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6787 = ~cache_hit ? meta_102_lru : _GEN_5235; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6788 = ~cache_hit ? meta_103_lru : _GEN_5236; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6789 = ~cache_hit ? meta_104_lru : _GEN_5237; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6790 = ~cache_hit ? meta_105_lru : _GEN_5238; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6791 = ~cache_hit ? meta_106_lru : _GEN_5239; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6792 = ~cache_hit ? meta_107_lru : _GEN_5240; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6793 = ~cache_hit ? meta_108_lru : _GEN_5241; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6794 = ~cache_hit ? meta_109_lru : _GEN_5242; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6795 = ~cache_hit ? meta_110_lru : _GEN_5243; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6796 = ~cache_hit ? meta_111_lru : _GEN_5244; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6797 = ~cache_hit ? meta_112_lru : _GEN_5245; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6798 = ~cache_hit ? meta_113_lru : _GEN_5246; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6799 = ~cache_hit ? meta_114_lru : _GEN_5247; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6800 = ~cache_hit ? meta_115_lru : _GEN_5248; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6801 = ~cache_hit ? meta_116_lru : _GEN_5249; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6802 = ~cache_hit ? meta_117_lru : _GEN_5250; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6803 = ~cache_hit ? meta_118_lru : _GEN_5251; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6804 = ~cache_hit ? meta_119_lru : _GEN_5252; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6805 = ~cache_hit ? meta_120_lru : _GEN_5253; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6806 = ~cache_hit ? meta_121_lru : _GEN_5254; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6807 = ~cache_hit ? meta_122_lru : _GEN_5255; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6808 = ~cache_hit ? meta_123_lru : _GEN_5256; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6809 = ~cache_hit ? meta_124_lru : _GEN_5257; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6810 = ~cache_hit ? meta_125_lru : _GEN_5258; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6811 = ~cache_hit ? meta_126_lru : _GEN_5259; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6812 = ~cache_hit ? meta_127_lru : _GEN_5260; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6813 = ~cache_hit ? meta_128_lru : _GEN_5261; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6814 = ~cache_hit ? meta_129_lru : _GEN_5262; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6815 = ~cache_hit ? meta_130_lru : _GEN_5263; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6816 = ~cache_hit ? meta_131_lru : _GEN_5264; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6817 = ~cache_hit ? meta_132_lru : _GEN_5265; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6818 = ~cache_hit ? meta_133_lru : _GEN_5266; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6819 = ~cache_hit ? meta_134_lru : _GEN_5267; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6820 = ~cache_hit ? meta_135_lru : _GEN_5268; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6821 = ~cache_hit ? meta_136_lru : _GEN_5269; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6822 = ~cache_hit ? meta_137_lru : _GEN_5270; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6823 = ~cache_hit ? meta_138_lru : _GEN_5271; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6824 = ~cache_hit ? meta_139_lru : _GEN_5272; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6825 = ~cache_hit ? meta_140_lru : _GEN_5273; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6826 = ~cache_hit ? meta_141_lru : _GEN_5274; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6827 = ~cache_hit ? meta_142_lru : _GEN_5275; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6828 = ~cache_hit ? meta_143_lru : _GEN_5276; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6829 = ~cache_hit ? meta_144_lru : _GEN_5277; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6830 = ~cache_hit ? meta_145_lru : _GEN_5278; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6831 = ~cache_hit ? meta_146_lru : _GEN_5279; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6832 = ~cache_hit ? meta_147_lru : _GEN_5280; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6833 = ~cache_hit ? meta_148_lru : _GEN_5281; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6834 = ~cache_hit ? meta_149_lru : _GEN_5282; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6835 = ~cache_hit ? meta_150_lru : _GEN_5283; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6836 = ~cache_hit ? meta_151_lru : _GEN_5284; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6837 = ~cache_hit ? meta_152_lru : _GEN_5285; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6838 = ~cache_hit ? meta_153_lru : _GEN_5286; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6839 = ~cache_hit ? meta_154_lru : _GEN_5287; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6840 = ~cache_hit ? meta_155_lru : _GEN_5288; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6841 = ~cache_hit ? meta_156_lru : _GEN_5289; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6842 = ~cache_hit ? meta_157_lru : _GEN_5290; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6843 = ~cache_hit ? meta_158_lru : _GEN_5291; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6844 = ~cache_hit ? meta_159_lru : _GEN_5292; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6845 = ~cache_hit ? meta_160_lru : _GEN_5293; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6846 = ~cache_hit ? meta_161_lru : _GEN_5294; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6847 = ~cache_hit ? meta_162_lru : _GEN_5295; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6848 = ~cache_hit ? meta_163_lru : _GEN_5296; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6849 = ~cache_hit ? meta_164_lru : _GEN_5297; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6850 = ~cache_hit ? meta_165_lru : _GEN_5298; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6851 = ~cache_hit ? meta_166_lru : _GEN_5299; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6852 = ~cache_hit ? meta_167_lru : _GEN_5300; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6853 = ~cache_hit ? meta_168_lru : _GEN_5301; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6854 = ~cache_hit ? meta_169_lru : _GEN_5302; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6855 = ~cache_hit ? meta_170_lru : _GEN_5303; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6856 = ~cache_hit ? meta_171_lru : _GEN_5304; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6857 = ~cache_hit ? meta_172_lru : _GEN_5305; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6858 = ~cache_hit ? meta_173_lru : _GEN_5306; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6859 = ~cache_hit ? meta_174_lru : _GEN_5307; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6860 = ~cache_hit ? meta_175_lru : _GEN_5308; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6861 = ~cache_hit ? meta_176_lru : _GEN_5309; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6862 = ~cache_hit ? meta_177_lru : _GEN_5310; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6863 = ~cache_hit ? meta_178_lru : _GEN_5311; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6864 = ~cache_hit ? meta_179_lru : _GEN_5312; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6865 = ~cache_hit ? meta_180_lru : _GEN_5313; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6866 = ~cache_hit ? meta_181_lru : _GEN_5314; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6867 = ~cache_hit ? meta_182_lru : _GEN_5315; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6868 = ~cache_hit ? meta_183_lru : _GEN_5316; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6869 = ~cache_hit ? meta_184_lru : _GEN_5317; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6870 = ~cache_hit ? meta_185_lru : _GEN_5318; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6871 = ~cache_hit ? meta_186_lru : _GEN_5319; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6872 = ~cache_hit ? meta_187_lru : _GEN_5320; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6873 = ~cache_hit ? meta_188_lru : _GEN_5321; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6874 = ~cache_hit ? meta_189_lru : _GEN_5322; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6875 = ~cache_hit ? meta_190_lru : _GEN_5323; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6876 = ~cache_hit ? meta_191_lru : _GEN_5324; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6877 = ~cache_hit ? meta_192_lru : _GEN_5325; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6878 = ~cache_hit ? meta_193_lru : _GEN_5326; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6879 = ~cache_hit ? meta_194_lru : _GEN_5327; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6880 = ~cache_hit ? meta_195_lru : _GEN_5328; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6881 = ~cache_hit ? meta_196_lru : _GEN_5329; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6882 = ~cache_hit ? meta_197_lru : _GEN_5330; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6883 = ~cache_hit ? meta_198_lru : _GEN_5331; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6884 = ~cache_hit ? meta_199_lru : _GEN_5332; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6885 = ~cache_hit ? meta_200_lru : _GEN_5333; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6886 = ~cache_hit ? meta_201_lru : _GEN_5334; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6887 = ~cache_hit ? meta_202_lru : _GEN_5335; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6888 = ~cache_hit ? meta_203_lru : _GEN_5336; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6889 = ~cache_hit ? meta_204_lru : _GEN_5337; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6890 = ~cache_hit ? meta_205_lru : _GEN_5338; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6891 = ~cache_hit ? meta_206_lru : _GEN_5339; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6892 = ~cache_hit ? meta_207_lru : _GEN_5340; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6893 = ~cache_hit ? meta_208_lru : _GEN_5341; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6894 = ~cache_hit ? meta_209_lru : _GEN_5342; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6895 = ~cache_hit ? meta_210_lru : _GEN_5343; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6896 = ~cache_hit ? meta_211_lru : _GEN_5344; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6897 = ~cache_hit ? meta_212_lru : _GEN_5345; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6898 = ~cache_hit ? meta_213_lru : _GEN_5346; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6899 = ~cache_hit ? meta_214_lru : _GEN_5347; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6900 = ~cache_hit ? meta_215_lru : _GEN_5348; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6901 = ~cache_hit ? meta_216_lru : _GEN_5349; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6902 = ~cache_hit ? meta_217_lru : _GEN_5350; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6903 = ~cache_hit ? meta_218_lru : _GEN_5351; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6904 = ~cache_hit ? meta_219_lru : _GEN_5352; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6905 = ~cache_hit ? meta_220_lru : _GEN_5353; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6906 = ~cache_hit ? meta_221_lru : _GEN_5354; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6907 = ~cache_hit ? meta_222_lru : _GEN_5355; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6908 = ~cache_hit ? meta_223_lru : _GEN_5356; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6909 = ~cache_hit ? meta_224_lru : _GEN_5357; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6910 = ~cache_hit ? meta_225_lru : _GEN_5358; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6911 = ~cache_hit ? meta_226_lru : _GEN_5359; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6912 = ~cache_hit ? meta_227_lru : _GEN_5360; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6913 = ~cache_hit ? meta_228_lru : _GEN_5361; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6914 = ~cache_hit ? meta_229_lru : _GEN_5362; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6915 = ~cache_hit ? meta_230_lru : _GEN_5363; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6916 = ~cache_hit ? meta_231_lru : _GEN_5364; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6917 = ~cache_hit ? meta_232_lru : _GEN_5365; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6918 = ~cache_hit ? meta_233_lru : _GEN_5366; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6919 = ~cache_hit ? meta_234_lru : _GEN_5367; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6920 = ~cache_hit ? meta_235_lru : _GEN_5368; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6921 = ~cache_hit ? meta_236_lru : _GEN_5369; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6922 = ~cache_hit ? meta_237_lru : _GEN_5370; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6923 = ~cache_hit ? meta_238_lru : _GEN_5371; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6924 = ~cache_hit ? meta_239_lru : _GEN_5372; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6925 = ~cache_hit ? meta_240_lru : _GEN_5373; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6926 = ~cache_hit ? meta_241_lru : _GEN_5374; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6927 = ~cache_hit ? meta_242_lru : _GEN_5375; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6928 = ~cache_hit ? meta_243_lru : _GEN_5376; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6929 = ~cache_hit ? meta_244_lru : _GEN_5377; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6930 = ~cache_hit ? meta_245_lru : _GEN_5378; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6931 = ~cache_hit ? meta_246_lru : _GEN_5379; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6932 = ~cache_hit ? meta_247_lru : _GEN_5380; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6933 = ~cache_hit ? meta_248_lru : _GEN_5381; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6934 = ~cache_hit ? meta_249_lru : _GEN_5382; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6935 = ~cache_hit ? meta_250_lru : _GEN_5383; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6936 = ~cache_hit ? meta_251_lru : _GEN_5384; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6937 = ~cache_hit ? meta_252_lru : _GEN_5385; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6938 = ~cache_hit ? meta_253_lru : _GEN_5386; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6939 = ~cache_hit ? meta_254_lru : _GEN_5387; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6940 = ~cache_hit ? meta_255_lru : _GEN_5388; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6941 = ~cache_hit ? meta_256_lru : _GEN_5389; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6942 = ~cache_hit ? meta_257_lru : _GEN_5390; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6943 = ~cache_hit ? meta_258_lru : _GEN_5391; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6944 = ~cache_hit ? meta_259_lru : _GEN_5392; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6945 = ~cache_hit ? meta_260_lru : _GEN_5393; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6946 = ~cache_hit ? meta_261_lru : _GEN_5394; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6947 = ~cache_hit ? meta_262_lru : _GEN_5395; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6948 = ~cache_hit ? meta_263_lru : _GEN_5396; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6949 = ~cache_hit ? meta_264_lru : _GEN_5397; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6950 = ~cache_hit ? meta_265_lru : _GEN_5398; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6951 = ~cache_hit ? meta_266_lru : _GEN_5399; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6952 = ~cache_hit ? meta_267_lru : _GEN_5400; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6953 = ~cache_hit ? meta_268_lru : _GEN_5401; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6954 = ~cache_hit ? meta_269_lru : _GEN_5402; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6955 = ~cache_hit ? meta_270_lru : _GEN_5403; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6956 = ~cache_hit ? meta_271_lru : _GEN_5404; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6957 = ~cache_hit ? meta_272_lru : _GEN_5405; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6958 = ~cache_hit ? meta_273_lru : _GEN_5406; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6959 = ~cache_hit ? meta_274_lru : _GEN_5407; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6960 = ~cache_hit ? meta_275_lru : _GEN_5408; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6961 = ~cache_hit ? meta_276_lru : _GEN_5409; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6962 = ~cache_hit ? meta_277_lru : _GEN_5410; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6963 = ~cache_hit ? meta_278_lru : _GEN_5411; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6964 = ~cache_hit ? meta_279_lru : _GEN_5412; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6965 = ~cache_hit ? meta_280_lru : _GEN_5413; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6966 = ~cache_hit ? meta_281_lru : _GEN_5414; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6967 = ~cache_hit ? meta_282_lru : _GEN_5415; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6968 = ~cache_hit ? meta_283_lru : _GEN_5416; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6969 = ~cache_hit ? meta_284_lru : _GEN_5417; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6970 = ~cache_hit ? meta_285_lru : _GEN_5418; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6971 = ~cache_hit ? meta_286_lru : _GEN_5419; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6972 = ~cache_hit ? meta_287_lru : _GEN_5420; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6973 = ~cache_hit ? meta_288_lru : _GEN_5421; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6974 = ~cache_hit ? meta_289_lru : _GEN_5422; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6975 = ~cache_hit ? meta_290_lru : _GEN_5423; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6976 = ~cache_hit ? meta_291_lru : _GEN_5424; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6977 = ~cache_hit ? meta_292_lru : _GEN_5425; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6978 = ~cache_hit ? meta_293_lru : _GEN_5426; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6979 = ~cache_hit ? meta_294_lru : _GEN_5427; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6980 = ~cache_hit ? meta_295_lru : _GEN_5428; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6981 = ~cache_hit ? meta_296_lru : _GEN_5429; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6982 = ~cache_hit ? meta_297_lru : _GEN_5430; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6983 = ~cache_hit ? meta_298_lru : _GEN_5431; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6984 = ~cache_hit ? meta_299_lru : _GEN_5432; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6985 = ~cache_hit ? meta_300_lru : _GEN_5433; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6986 = ~cache_hit ? meta_301_lru : _GEN_5434; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6987 = ~cache_hit ? meta_302_lru : _GEN_5435; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6988 = ~cache_hit ? meta_303_lru : _GEN_5436; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6989 = ~cache_hit ? meta_304_lru : _GEN_5437; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6990 = ~cache_hit ? meta_305_lru : _GEN_5438; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6991 = ~cache_hit ? meta_306_lru : _GEN_5439; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6992 = ~cache_hit ? meta_307_lru : _GEN_5440; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6993 = ~cache_hit ? meta_308_lru : _GEN_5441; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6994 = ~cache_hit ? meta_309_lru : _GEN_5442; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6995 = ~cache_hit ? meta_310_lru : _GEN_5443; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6996 = ~cache_hit ? meta_311_lru : _GEN_5444; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6997 = ~cache_hit ? meta_312_lru : _GEN_5445; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6998 = ~cache_hit ? meta_313_lru : _GEN_5446; // @[ICache.scala 175:32 34:21]
  wire  _GEN_6999 = ~cache_hit ? meta_314_lru : _GEN_5447; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7000 = ~cache_hit ? meta_315_lru : _GEN_5448; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7001 = ~cache_hit ? meta_316_lru : _GEN_5449; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7002 = ~cache_hit ? meta_317_lru : _GEN_5450; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7003 = ~cache_hit ? meta_318_lru : _GEN_5451; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7004 = ~cache_hit ? meta_319_lru : _GEN_5452; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7005 = ~cache_hit ? meta_320_lru : _GEN_5453; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7006 = ~cache_hit ? meta_321_lru : _GEN_5454; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7007 = ~cache_hit ? meta_322_lru : _GEN_5455; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7008 = ~cache_hit ? meta_323_lru : _GEN_5456; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7009 = ~cache_hit ? meta_324_lru : _GEN_5457; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7010 = ~cache_hit ? meta_325_lru : _GEN_5458; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7011 = ~cache_hit ? meta_326_lru : _GEN_5459; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7012 = ~cache_hit ? meta_327_lru : _GEN_5460; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7013 = ~cache_hit ? meta_328_lru : _GEN_5461; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7014 = ~cache_hit ? meta_329_lru : _GEN_5462; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7015 = ~cache_hit ? meta_330_lru : _GEN_5463; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7016 = ~cache_hit ? meta_331_lru : _GEN_5464; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7017 = ~cache_hit ? meta_332_lru : _GEN_5465; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7018 = ~cache_hit ? meta_333_lru : _GEN_5466; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7019 = ~cache_hit ? meta_334_lru : _GEN_5467; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7020 = ~cache_hit ? meta_335_lru : _GEN_5468; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7021 = ~cache_hit ? meta_336_lru : _GEN_5469; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7022 = ~cache_hit ? meta_337_lru : _GEN_5470; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7023 = ~cache_hit ? meta_338_lru : _GEN_5471; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7024 = ~cache_hit ? meta_339_lru : _GEN_5472; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7025 = ~cache_hit ? meta_340_lru : _GEN_5473; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7026 = ~cache_hit ? meta_341_lru : _GEN_5474; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7027 = ~cache_hit ? meta_342_lru : _GEN_5475; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7028 = ~cache_hit ? meta_343_lru : _GEN_5476; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7029 = ~cache_hit ? meta_344_lru : _GEN_5477; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7030 = ~cache_hit ? meta_345_lru : _GEN_5478; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7031 = ~cache_hit ? meta_346_lru : _GEN_5479; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7032 = ~cache_hit ? meta_347_lru : _GEN_5480; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7033 = ~cache_hit ? meta_348_lru : _GEN_5481; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7034 = ~cache_hit ? meta_349_lru : _GEN_5482; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7035 = ~cache_hit ? meta_350_lru : _GEN_5483; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7036 = ~cache_hit ? meta_351_lru : _GEN_5484; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7037 = ~cache_hit ? meta_352_lru : _GEN_5485; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7038 = ~cache_hit ? meta_353_lru : _GEN_5486; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7039 = ~cache_hit ? meta_354_lru : _GEN_5487; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7040 = ~cache_hit ? meta_355_lru : _GEN_5488; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7041 = ~cache_hit ? meta_356_lru : _GEN_5489; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7042 = ~cache_hit ? meta_357_lru : _GEN_5490; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7043 = ~cache_hit ? meta_358_lru : _GEN_5491; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7044 = ~cache_hit ? meta_359_lru : _GEN_5492; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7045 = ~cache_hit ? meta_360_lru : _GEN_5493; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7046 = ~cache_hit ? meta_361_lru : _GEN_5494; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7047 = ~cache_hit ? meta_362_lru : _GEN_5495; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7048 = ~cache_hit ? meta_363_lru : _GEN_5496; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7049 = ~cache_hit ? meta_364_lru : _GEN_5497; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7050 = ~cache_hit ? meta_365_lru : _GEN_5498; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7051 = ~cache_hit ? meta_366_lru : _GEN_5499; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7052 = ~cache_hit ? meta_367_lru : _GEN_5500; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7053 = ~cache_hit ? meta_368_lru : _GEN_5501; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7054 = ~cache_hit ? meta_369_lru : _GEN_5502; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7055 = ~cache_hit ? meta_370_lru : _GEN_5503; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7056 = ~cache_hit ? meta_371_lru : _GEN_5504; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7057 = ~cache_hit ? meta_372_lru : _GEN_5505; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7058 = ~cache_hit ? meta_373_lru : _GEN_5506; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7059 = ~cache_hit ? meta_374_lru : _GEN_5507; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7060 = ~cache_hit ? meta_375_lru : _GEN_5508; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7061 = ~cache_hit ? meta_376_lru : _GEN_5509; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7062 = ~cache_hit ? meta_377_lru : _GEN_5510; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7063 = ~cache_hit ? meta_378_lru : _GEN_5511; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7064 = ~cache_hit ? meta_379_lru : _GEN_5512; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7065 = ~cache_hit ? meta_380_lru : _GEN_5513; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7066 = ~cache_hit ? meta_381_lru : _GEN_5514; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7067 = ~cache_hit ? meta_382_lru : _GEN_5515; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7068 = ~cache_hit ? meta_383_lru : _GEN_5516; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7069 = ~cache_hit ? meta_384_lru : _GEN_5517; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7070 = ~cache_hit ? meta_385_lru : _GEN_5518; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7071 = ~cache_hit ? meta_386_lru : _GEN_5519; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7072 = ~cache_hit ? meta_387_lru : _GEN_5520; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7073 = ~cache_hit ? meta_388_lru : _GEN_5521; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7074 = ~cache_hit ? meta_389_lru : _GEN_5522; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7075 = ~cache_hit ? meta_390_lru : _GEN_5523; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7076 = ~cache_hit ? meta_391_lru : _GEN_5524; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7077 = ~cache_hit ? meta_392_lru : _GEN_5525; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7078 = ~cache_hit ? meta_393_lru : _GEN_5526; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7079 = ~cache_hit ? meta_394_lru : _GEN_5527; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7080 = ~cache_hit ? meta_395_lru : _GEN_5528; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7081 = ~cache_hit ? meta_396_lru : _GEN_5529; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7082 = ~cache_hit ? meta_397_lru : _GEN_5530; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7083 = ~cache_hit ? meta_398_lru : _GEN_5531; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7084 = ~cache_hit ? meta_399_lru : _GEN_5532; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7085 = ~cache_hit ? meta_400_lru : _GEN_5533; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7086 = ~cache_hit ? meta_401_lru : _GEN_5534; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7087 = ~cache_hit ? meta_402_lru : _GEN_5535; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7088 = ~cache_hit ? meta_403_lru : _GEN_5536; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7089 = ~cache_hit ? meta_404_lru : _GEN_5537; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7090 = ~cache_hit ? meta_405_lru : _GEN_5538; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7091 = ~cache_hit ? meta_406_lru : _GEN_5539; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7092 = ~cache_hit ? meta_407_lru : _GEN_5540; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7093 = ~cache_hit ? meta_408_lru : _GEN_5541; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7094 = ~cache_hit ? meta_409_lru : _GEN_5542; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7095 = ~cache_hit ? meta_410_lru : _GEN_5543; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7096 = ~cache_hit ? meta_411_lru : _GEN_5544; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7097 = ~cache_hit ? meta_412_lru : _GEN_5545; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7098 = ~cache_hit ? meta_413_lru : _GEN_5546; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7099 = ~cache_hit ? meta_414_lru : _GEN_5547; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7100 = ~cache_hit ? meta_415_lru : _GEN_5548; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7101 = ~cache_hit ? meta_416_lru : _GEN_5549; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7102 = ~cache_hit ? meta_417_lru : _GEN_5550; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7103 = ~cache_hit ? meta_418_lru : _GEN_5551; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7104 = ~cache_hit ? meta_419_lru : _GEN_5552; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7105 = ~cache_hit ? meta_420_lru : _GEN_5553; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7106 = ~cache_hit ? meta_421_lru : _GEN_5554; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7107 = ~cache_hit ? meta_422_lru : _GEN_5555; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7108 = ~cache_hit ? meta_423_lru : _GEN_5556; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7109 = ~cache_hit ? meta_424_lru : _GEN_5557; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7110 = ~cache_hit ? meta_425_lru : _GEN_5558; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7111 = ~cache_hit ? meta_426_lru : _GEN_5559; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7112 = ~cache_hit ? meta_427_lru : _GEN_5560; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7113 = ~cache_hit ? meta_428_lru : _GEN_5561; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7114 = ~cache_hit ? meta_429_lru : _GEN_5562; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7115 = ~cache_hit ? meta_430_lru : _GEN_5563; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7116 = ~cache_hit ? meta_431_lru : _GEN_5564; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7117 = ~cache_hit ? meta_432_lru : _GEN_5565; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7118 = ~cache_hit ? meta_433_lru : _GEN_5566; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7119 = ~cache_hit ? meta_434_lru : _GEN_5567; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7120 = ~cache_hit ? meta_435_lru : _GEN_5568; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7121 = ~cache_hit ? meta_436_lru : _GEN_5569; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7122 = ~cache_hit ? meta_437_lru : _GEN_5570; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7123 = ~cache_hit ? meta_438_lru : _GEN_5571; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7124 = ~cache_hit ? meta_439_lru : _GEN_5572; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7125 = ~cache_hit ? meta_440_lru : _GEN_5573; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7126 = ~cache_hit ? meta_441_lru : _GEN_5574; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7127 = ~cache_hit ? meta_442_lru : _GEN_5575; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7128 = ~cache_hit ? meta_443_lru : _GEN_5576; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7129 = ~cache_hit ? meta_444_lru : _GEN_5577; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7130 = ~cache_hit ? meta_445_lru : _GEN_5578; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7131 = ~cache_hit ? meta_446_lru : _GEN_5579; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7132 = ~cache_hit ? meta_447_lru : _GEN_5580; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7133 = ~cache_hit ? meta_448_lru : _GEN_5581; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7134 = ~cache_hit ? meta_449_lru : _GEN_5582; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7135 = ~cache_hit ? meta_450_lru : _GEN_5583; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7136 = ~cache_hit ? meta_451_lru : _GEN_5584; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7137 = ~cache_hit ? meta_452_lru : _GEN_5585; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7138 = ~cache_hit ? meta_453_lru : _GEN_5586; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7139 = ~cache_hit ? meta_454_lru : _GEN_5587; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7140 = ~cache_hit ? meta_455_lru : _GEN_5588; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7141 = ~cache_hit ? meta_456_lru : _GEN_5589; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7142 = ~cache_hit ? meta_457_lru : _GEN_5590; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7143 = ~cache_hit ? meta_458_lru : _GEN_5591; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7144 = ~cache_hit ? meta_459_lru : _GEN_5592; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7145 = ~cache_hit ? meta_460_lru : _GEN_5593; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7146 = ~cache_hit ? meta_461_lru : _GEN_5594; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7147 = ~cache_hit ? meta_462_lru : _GEN_5595; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7148 = ~cache_hit ? meta_463_lru : _GEN_5596; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7149 = ~cache_hit ? meta_464_lru : _GEN_5597; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7150 = ~cache_hit ? meta_465_lru : _GEN_5598; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7151 = ~cache_hit ? meta_466_lru : _GEN_5599; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7152 = ~cache_hit ? meta_467_lru : _GEN_5600; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7153 = ~cache_hit ? meta_468_lru : _GEN_5601; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7154 = ~cache_hit ? meta_469_lru : _GEN_5602; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7155 = ~cache_hit ? meta_470_lru : _GEN_5603; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7156 = ~cache_hit ? meta_471_lru : _GEN_5604; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7157 = ~cache_hit ? meta_472_lru : _GEN_5605; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7158 = ~cache_hit ? meta_473_lru : _GEN_5606; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7159 = ~cache_hit ? meta_474_lru : _GEN_5607; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7160 = ~cache_hit ? meta_475_lru : _GEN_5608; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7161 = ~cache_hit ? meta_476_lru : _GEN_5609; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7162 = ~cache_hit ? meta_477_lru : _GEN_5610; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7163 = ~cache_hit ? meta_478_lru : _GEN_5611; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7164 = ~cache_hit ? meta_479_lru : _GEN_5612; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7165 = ~cache_hit ? meta_480_lru : _GEN_5613; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7166 = ~cache_hit ? meta_481_lru : _GEN_5614; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7167 = ~cache_hit ? meta_482_lru : _GEN_5615; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7168 = ~cache_hit ? meta_483_lru : _GEN_5616; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7169 = ~cache_hit ? meta_484_lru : _GEN_5617; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7170 = ~cache_hit ? meta_485_lru : _GEN_5618; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7171 = ~cache_hit ? meta_486_lru : _GEN_5619; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7172 = ~cache_hit ? meta_487_lru : _GEN_5620; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7173 = ~cache_hit ? meta_488_lru : _GEN_5621; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7174 = ~cache_hit ? meta_489_lru : _GEN_5622; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7175 = ~cache_hit ? meta_490_lru : _GEN_5623; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7176 = ~cache_hit ? meta_491_lru : _GEN_5624; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7177 = ~cache_hit ? meta_492_lru : _GEN_5625; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7178 = ~cache_hit ? meta_493_lru : _GEN_5626; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7179 = ~cache_hit ? meta_494_lru : _GEN_5627; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7180 = ~cache_hit ? meta_495_lru : _GEN_5628; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7181 = ~cache_hit ? meta_496_lru : _GEN_5629; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7182 = ~cache_hit ? meta_497_lru : _GEN_5630; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7183 = ~cache_hit ? meta_498_lru : _GEN_5631; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7184 = ~cache_hit ? meta_499_lru : _GEN_5632; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7185 = ~cache_hit ? meta_500_lru : _GEN_5633; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7186 = ~cache_hit ? meta_501_lru : _GEN_5634; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7187 = ~cache_hit ? meta_502_lru : _GEN_5635; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7188 = ~cache_hit ? meta_503_lru : _GEN_5636; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7189 = ~cache_hit ? meta_504_lru : _GEN_5637; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7190 = ~cache_hit ? meta_505_lru : _GEN_5638; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7191 = ~cache_hit ? meta_506_lru : _GEN_5639; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7192 = ~cache_hit ? meta_507_lru : _GEN_5640; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7193 = ~cache_hit ? meta_508_lru : _GEN_5641; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7194 = ~cache_hit ? meta_509_lru : _GEN_5642; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7195 = ~cache_hit ? meta_510_lru : _GEN_5643; // @[ICache.scala 175:32 34:21]
  wire  _GEN_7196 = ~cache_hit ? meta_511_lru : _GEN_5644; // @[ICache.scala 175:32 34:21]
  wire [63:0] _GEN_7197 = ~cache_hit ? {{32'd0}, saved_1_inst} : _GEN_5646; // @[ICache.scala 175:32 91:22]
  wire  _GEN_7198 = ~cache_hit ? saved_0_valid : _GEN_5647; // @[ICache.scala 175:32 91:22]
  wire  _GEN_7199 = ~cache_hit ? saved_1_valid : _GEN_5648; // @[ICache.scala 175:32 91:22]
  wire [2:0] _GEN_7200 = uncached ? 3'h2 : _GEN_5649; // @[ICache.scala 169:30 170:19]
  wire [31:0] _GEN_7201 = uncached ? inst_pa : _GEN_5650; // @[ICache.scala 169:30 171:19]
  wire [7:0] _GEN_7202 = uncached ? 8'h0 : _GEN_5651; // @[ICache.scala 169:30 172:19]
  wire [2:0] _GEN_7203 = uncached ? 3'h2 : _GEN_5652; // @[ICache.scala 169:30 173:19]
  wire  _GEN_7204 = uncached | _GEN_5653; // @[ICache.scala 169:30 174:19]
  wire [5:0] _GEN_7205 = uncached ? replace_line_addr : _GEN_5654; // @[ICache.scala 169:30 58:38]
  wire [7:0] _GEN_7206 = uncached ? data_wen_0 : _GEN_5655; // @[ICache.scala 169:30 66:30]
  wire [7:0] _GEN_7207 = uncached ? data_wen_1 : _GEN_5656; // @[ICache.scala 169:30 66:30]
  wire  _GEN_7208 = uncached ? tag_wen_0 : _GEN_5657; // @[ICache.scala 169:30 67:30]
  wire  _GEN_7209 = uncached ? tag_wen_1 : _GEN_5658; // @[ICache.scala 169:30 67:30]
  wire [19:0] _GEN_7210 = uncached ? {{3'd0}, tag_ram_wdata} : _GEN_5659; // @[ICache.scala 169:30 68:30]
  wire  _GEN_7211 = uncached ? _GEN_2053 : _GEN_5660; // @[ICache.scala 169:30]
  wire  _GEN_7212 = uncached ? _GEN_2565 : _GEN_5661; // @[ICache.scala 169:30]
  wire  _GEN_7213 = uncached ? _GEN_2054 : _GEN_5662; // @[ICache.scala 169:30]
  wire  _GEN_7214 = uncached ? _GEN_2566 : _GEN_5663; // @[ICache.scala 169:30]
  wire  _GEN_7215 = uncached ? _GEN_2055 : _GEN_5664; // @[ICache.scala 169:30]
  wire  _GEN_7216 = uncached ? _GEN_2567 : _GEN_5665; // @[ICache.scala 169:30]
  wire  _GEN_7217 = uncached ? _GEN_2056 : _GEN_5666; // @[ICache.scala 169:30]
  wire  _GEN_7218 = uncached ? _GEN_2568 : _GEN_5667; // @[ICache.scala 169:30]
  wire  _GEN_7219 = uncached ? _GEN_2057 : _GEN_5668; // @[ICache.scala 169:30]
  wire  _GEN_7220 = uncached ? _GEN_2569 : _GEN_5669; // @[ICache.scala 169:30]
  wire  _GEN_7221 = uncached ? _GEN_2058 : _GEN_5670; // @[ICache.scala 169:30]
  wire  _GEN_7222 = uncached ? _GEN_2570 : _GEN_5671; // @[ICache.scala 169:30]
  wire  _GEN_7223 = uncached ? _GEN_2059 : _GEN_5672; // @[ICache.scala 169:30]
  wire  _GEN_7224 = uncached ? _GEN_2571 : _GEN_5673; // @[ICache.scala 169:30]
  wire  _GEN_7225 = uncached ? _GEN_2060 : _GEN_5674; // @[ICache.scala 169:30]
  wire  _GEN_7226 = uncached ? _GEN_2572 : _GEN_5675; // @[ICache.scala 169:30]
  wire  _GEN_7227 = uncached ? _GEN_2061 : _GEN_5676; // @[ICache.scala 169:30]
  wire  _GEN_7228 = uncached ? _GEN_2573 : _GEN_5677; // @[ICache.scala 169:30]
  wire  _GEN_7229 = uncached ? _GEN_2062 : _GEN_5678; // @[ICache.scala 169:30]
  wire  _GEN_7230 = uncached ? _GEN_2574 : _GEN_5679; // @[ICache.scala 169:30]
  wire  _GEN_7231 = uncached ? _GEN_2063 : _GEN_5680; // @[ICache.scala 169:30]
  wire  _GEN_7232 = uncached ? _GEN_2575 : _GEN_5681; // @[ICache.scala 169:30]
  wire  _GEN_7233 = uncached ? _GEN_2064 : _GEN_5682; // @[ICache.scala 169:30]
  wire  _GEN_7234 = uncached ? _GEN_2576 : _GEN_5683; // @[ICache.scala 169:30]
  wire  _GEN_7235 = uncached ? _GEN_2065 : _GEN_5684; // @[ICache.scala 169:30]
  wire  _GEN_7236 = uncached ? _GEN_2577 : _GEN_5685; // @[ICache.scala 169:30]
  wire  _GEN_7237 = uncached ? _GEN_2066 : _GEN_5686; // @[ICache.scala 169:30]
  wire  _GEN_7238 = uncached ? _GEN_2578 : _GEN_5687; // @[ICache.scala 169:30]
  wire  _GEN_7239 = uncached ? _GEN_2067 : _GEN_5688; // @[ICache.scala 169:30]
  wire  _GEN_7240 = uncached ? _GEN_2579 : _GEN_5689; // @[ICache.scala 169:30]
  wire  _GEN_7241 = uncached ? _GEN_2068 : _GEN_5690; // @[ICache.scala 169:30]
  wire  _GEN_7242 = uncached ? _GEN_2580 : _GEN_5691; // @[ICache.scala 169:30]
  wire  _GEN_7243 = uncached ? _GEN_2069 : _GEN_5692; // @[ICache.scala 169:30]
  wire  _GEN_7244 = uncached ? _GEN_2581 : _GEN_5693; // @[ICache.scala 169:30]
  wire  _GEN_7245 = uncached ? _GEN_2070 : _GEN_5694; // @[ICache.scala 169:30]
  wire  _GEN_7246 = uncached ? _GEN_2582 : _GEN_5695; // @[ICache.scala 169:30]
  wire  _GEN_7247 = uncached ? _GEN_2071 : _GEN_5696; // @[ICache.scala 169:30]
  wire  _GEN_7248 = uncached ? _GEN_2583 : _GEN_5697; // @[ICache.scala 169:30]
  wire  _GEN_7249 = uncached ? _GEN_2072 : _GEN_5698; // @[ICache.scala 169:30]
  wire  _GEN_7250 = uncached ? _GEN_2584 : _GEN_5699; // @[ICache.scala 169:30]
  wire  _GEN_7251 = uncached ? _GEN_2073 : _GEN_5700; // @[ICache.scala 169:30]
  wire  _GEN_7252 = uncached ? _GEN_2585 : _GEN_5701; // @[ICache.scala 169:30]
  wire  _GEN_7253 = uncached ? _GEN_2074 : _GEN_5702; // @[ICache.scala 169:30]
  wire  _GEN_7254 = uncached ? _GEN_2586 : _GEN_5703; // @[ICache.scala 169:30]
  wire  _GEN_7255 = uncached ? _GEN_2075 : _GEN_5704; // @[ICache.scala 169:30]
  wire  _GEN_7256 = uncached ? _GEN_2587 : _GEN_5705; // @[ICache.scala 169:30]
  wire  _GEN_7257 = uncached ? _GEN_2076 : _GEN_5706; // @[ICache.scala 169:30]
  wire  _GEN_7258 = uncached ? _GEN_2588 : _GEN_5707; // @[ICache.scala 169:30]
  wire  _GEN_7259 = uncached ? _GEN_2077 : _GEN_5708; // @[ICache.scala 169:30]
  wire  _GEN_7260 = uncached ? _GEN_2589 : _GEN_5709; // @[ICache.scala 169:30]
  wire  _GEN_7261 = uncached ? _GEN_2078 : _GEN_5710; // @[ICache.scala 169:30]
  wire  _GEN_7262 = uncached ? _GEN_2590 : _GEN_5711; // @[ICache.scala 169:30]
  wire  _GEN_7263 = uncached ? _GEN_2079 : _GEN_5712; // @[ICache.scala 169:30]
  wire  _GEN_7264 = uncached ? _GEN_2591 : _GEN_5713; // @[ICache.scala 169:30]
  wire  _GEN_7265 = uncached ? _GEN_2080 : _GEN_5714; // @[ICache.scala 169:30]
  wire  _GEN_7266 = uncached ? _GEN_2592 : _GEN_5715; // @[ICache.scala 169:30]
  wire  _GEN_7267 = uncached ? _GEN_2081 : _GEN_5716; // @[ICache.scala 169:30]
  wire  _GEN_7268 = uncached ? _GEN_2593 : _GEN_5717; // @[ICache.scala 169:30]
  wire  _GEN_7269 = uncached ? _GEN_2082 : _GEN_5718; // @[ICache.scala 169:30]
  wire  _GEN_7270 = uncached ? _GEN_2594 : _GEN_5719; // @[ICache.scala 169:30]
  wire  _GEN_7271 = uncached ? _GEN_2083 : _GEN_5720; // @[ICache.scala 169:30]
  wire  _GEN_7272 = uncached ? _GEN_2595 : _GEN_5721; // @[ICache.scala 169:30]
  wire  _GEN_7273 = uncached ? _GEN_2084 : _GEN_5722; // @[ICache.scala 169:30]
  wire  _GEN_7274 = uncached ? _GEN_2596 : _GEN_5723; // @[ICache.scala 169:30]
  wire  _GEN_7275 = uncached ? _GEN_2085 : _GEN_5724; // @[ICache.scala 169:30]
  wire  _GEN_7276 = uncached ? _GEN_2597 : _GEN_5725; // @[ICache.scala 169:30]
  wire  _GEN_7277 = uncached ? _GEN_2086 : _GEN_5726; // @[ICache.scala 169:30]
  wire  _GEN_7278 = uncached ? _GEN_2598 : _GEN_5727; // @[ICache.scala 169:30]
  wire  _GEN_7279 = uncached ? _GEN_2087 : _GEN_5728; // @[ICache.scala 169:30]
  wire  _GEN_7280 = uncached ? _GEN_2599 : _GEN_5729; // @[ICache.scala 169:30]
  wire  _GEN_7281 = uncached ? _GEN_2088 : _GEN_5730; // @[ICache.scala 169:30]
  wire  _GEN_7282 = uncached ? _GEN_2600 : _GEN_5731; // @[ICache.scala 169:30]
  wire  _GEN_7283 = uncached ? _GEN_2089 : _GEN_5732; // @[ICache.scala 169:30]
  wire  _GEN_7284 = uncached ? _GEN_2601 : _GEN_5733; // @[ICache.scala 169:30]
  wire  _GEN_7285 = uncached ? _GEN_2090 : _GEN_5734; // @[ICache.scala 169:30]
  wire  _GEN_7286 = uncached ? _GEN_2602 : _GEN_5735; // @[ICache.scala 169:30]
  wire  _GEN_7287 = uncached ? _GEN_2091 : _GEN_5736; // @[ICache.scala 169:30]
  wire  _GEN_7288 = uncached ? _GEN_2603 : _GEN_5737; // @[ICache.scala 169:30]
  wire  _GEN_7289 = uncached ? _GEN_2092 : _GEN_5738; // @[ICache.scala 169:30]
  wire  _GEN_7290 = uncached ? _GEN_2604 : _GEN_5739; // @[ICache.scala 169:30]
  wire  _GEN_7291 = uncached ? _GEN_2093 : _GEN_5740; // @[ICache.scala 169:30]
  wire  _GEN_7292 = uncached ? _GEN_2605 : _GEN_5741; // @[ICache.scala 169:30]
  wire  _GEN_7293 = uncached ? _GEN_2094 : _GEN_5742; // @[ICache.scala 169:30]
  wire  _GEN_7294 = uncached ? _GEN_2606 : _GEN_5743; // @[ICache.scala 169:30]
  wire  _GEN_7295 = uncached ? _GEN_2095 : _GEN_5744; // @[ICache.scala 169:30]
  wire  _GEN_7296 = uncached ? _GEN_2607 : _GEN_5745; // @[ICache.scala 169:30]
  wire  _GEN_7297 = uncached ? _GEN_2096 : _GEN_5746; // @[ICache.scala 169:30]
  wire  _GEN_7298 = uncached ? _GEN_2608 : _GEN_5747; // @[ICache.scala 169:30]
  wire  _GEN_7299 = uncached ? _GEN_2097 : _GEN_5748; // @[ICache.scala 169:30]
  wire  _GEN_7300 = uncached ? _GEN_2609 : _GEN_5749; // @[ICache.scala 169:30]
  wire  _GEN_7301 = uncached ? _GEN_2098 : _GEN_5750; // @[ICache.scala 169:30]
  wire  _GEN_7302 = uncached ? _GEN_2610 : _GEN_5751; // @[ICache.scala 169:30]
  wire  _GEN_7303 = uncached ? _GEN_2099 : _GEN_5752; // @[ICache.scala 169:30]
  wire  _GEN_7304 = uncached ? _GEN_2611 : _GEN_5753; // @[ICache.scala 169:30]
  wire  _GEN_7305 = uncached ? _GEN_2100 : _GEN_5754; // @[ICache.scala 169:30]
  wire  _GEN_7306 = uncached ? _GEN_2612 : _GEN_5755; // @[ICache.scala 169:30]
  wire  _GEN_7307 = uncached ? _GEN_2101 : _GEN_5756; // @[ICache.scala 169:30]
  wire  _GEN_7308 = uncached ? _GEN_2613 : _GEN_5757; // @[ICache.scala 169:30]
  wire  _GEN_7309 = uncached ? _GEN_2102 : _GEN_5758; // @[ICache.scala 169:30]
  wire  _GEN_7310 = uncached ? _GEN_2614 : _GEN_5759; // @[ICache.scala 169:30]
  wire  _GEN_7311 = uncached ? _GEN_2103 : _GEN_5760; // @[ICache.scala 169:30]
  wire  _GEN_7312 = uncached ? _GEN_2615 : _GEN_5761; // @[ICache.scala 169:30]
  wire  _GEN_7313 = uncached ? _GEN_2104 : _GEN_5762; // @[ICache.scala 169:30]
  wire  _GEN_7314 = uncached ? _GEN_2616 : _GEN_5763; // @[ICache.scala 169:30]
  wire  _GEN_7315 = uncached ? _GEN_2105 : _GEN_5764; // @[ICache.scala 169:30]
  wire  _GEN_7316 = uncached ? _GEN_2617 : _GEN_5765; // @[ICache.scala 169:30]
  wire  _GEN_7317 = uncached ? _GEN_2106 : _GEN_5766; // @[ICache.scala 169:30]
  wire  _GEN_7318 = uncached ? _GEN_2618 : _GEN_5767; // @[ICache.scala 169:30]
  wire  _GEN_7319 = uncached ? _GEN_2107 : _GEN_5768; // @[ICache.scala 169:30]
  wire  _GEN_7320 = uncached ? _GEN_2619 : _GEN_5769; // @[ICache.scala 169:30]
  wire  _GEN_7321 = uncached ? _GEN_2108 : _GEN_5770; // @[ICache.scala 169:30]
  wire  _GEN_7322 = uncached ? _GEN_2620 : _GEN_5771; // @[ICache.scala 169:30]
  wire  _GEN_7323 = uncached ? _GEN_2109 : _GEN_5772; // @[ICache.scala 169:30]
  wire  _GEN_7324 = uncached ? _GEN_2621 : _GEN_5773; // @[ICache.scala 169:30]
  wire  _GEN_7325 = uncached ? _GEN_2110 : _GEN_5774; // @[ICache.scala 169:30]
  wire  _GEN_7326 = uncached ? _GEN_2622 : _GEN_5775; // @[ICache.scala 169:30]
  wire  _GEN_7327 = uncached ? _GEN_2111 : _GEN_5776; // @[ICache.scala 169:30]
  wire  _GEN_7328 = uncached ? _GEN_2623 : _GEN_5777; // @[ICache.scala 169:30]
  wire  _GEN_7329 = uncached ? _GEN_2112 : _GEN_5778; // @[ICache.scala 169:30]
  wire  _GEN_7330 = uncached ? _GEN_2624 : _GEN_5779; // @[ICache.scala 169:30]
  wire  _GEN_7331 = uncached ? _GEN_2113 : _GEN_5780; // @[ICache.scala 169:30]
  wire  _GEN_7332 = uncached ? _GEN_2625 : _GEN_5781; // @[ICache.scala 169:30]
  wire  _GEN_7333 = uncached ? _GEN_2114 : _GEN_5782; // @[ICache.scala 169:30]
  wire  _GEN_7334 = uncached ? _GEN_2626 : _GEN_5783; // @[ICache.scala 169:30]
  wire  _GEN_7335 = uncached ? _GEN_2115 : _GEN_5784; // @[ICache.scala 169:30]
  wire  _GEN_7336 = uncached ? _GEN_2627 : _GEN_5785; // @[ICache.scala 169:30]
  wire  _GEN_7337 = uncached ? _GEN_2116 : _GEN_5786; // @[ICache.scala 169:30]
  wire  _GEN_7338 = uncached ? _GEN_2628 : _GEN_5787; // @[ICache.scala 169:30]
  wire  _GEN_7339 = uncached ? _GEN_2117 : _GEN_5788; // @[ICache.scala 169:30]
  wire  _GEN_7340 = uncached ? _GEN_2629 : _GEN_5789; // @[ICache.scala 169:30]
  wire  _GEN_7341 = uncached ? _GEN_2118 : _GEN_5790; // @[ICache.scala 169:30]
  wire  _GEN_7342 = uncached ? _GEN_2630 : _GEN_5791; // @[ICache.scala 169:30]
  wire  _GEN_7343 = uncached ? _GEN_2119 : _GEN_5792; // @[ICache.scala 169:30]
  wire  _GEN_7344 = uncached ? _GEN_2631 : _GEN_5793; // @[ICache.scala 169:30]
  wire  _GEN_7345 = uncached ? _GEN_2120 : _GEN_5794; // @[ICache.scala 169:30]
  wire  _GEN_7346 = uncached ? _GEN_2632 : _GEN_5795; // @[ICache.scala 169:30]
  wire  _GEN_7347 = uncached ? _GEN_2121 : _GEN_5796; // @[ICache.scala 169:30]
  wire  _GEN_7348 = uncached ? _GEN_2633 : _GEN_5797; // @[ICache.scala 169:30]
  wire  _GEN_7349 = uncached ? _GEN_2122 : _GEN_5798; // @[ICache.scala 169:30]
  wire  _GEN_7350 = uncached ? _GEN_2634 : _GEN_5799; // @[ICache.scala 169:30]
  wire  _GEN_7351 = uncached ? _GEN_2123 : _GEN_5800; // @[ICache.scala 169:30]
  wire  _GEN_7352 = uncached ? _GEN_2635 : _GEN_5801; // @[ICache.scala 169:30]
  wire  _GEN_7353 = uncached ? _GEN_2124 : _GEN_5802; // @[ICache.scala 169:30]
  wire  _GEN_7354 = uncached ? _GEN_2636 : _GEN_5803; // @[ICache.scala 169:30]
  wire  _GEN_7355 = uncached ? _GEN_2125 : _GEN_5804; // @[ICache.scala 169:30]
  wire  _GEN_7356 = uncached ? _GEN_2637 : _GEN_5805; // @[ICache.scala 169:30]
  wire  _GEN_7357 = uncached ? _GEN_2126 : _GEN_5806; // @[ICache.scala 169:30]
  wire  _GEN_7358 = uncached ? _GEN_2638 : _GEN_5807; // @[ICache.scala 169:30]
  wire  _GEN_7359 = uncached ? _GEN_2127 : _GEN_5808; // @[ICache.scala 169:30]
  wire  _GEN_7360 = uncached ? _GEN_2639 : _GEN_5809; // @[ICache.scala 169:30]
  wire  _GEN_7361 = uncached ? _GEN_2128 : _GEN_5810; // @[ICache.scala 169:30]
  wire  _GEN_7362 = uncached ? _GEN_2640 : _GEN_5811; // @[ICache.scala 169:30]
  wire  _GEN_7363 = uncached ? _GEN_2129 : _GEN_5812; // @[ICache.scala 169:30]
  wire  _GEN_7364 = uncached ? _GEN_2641 : _GEN_5813; // @[ICache.scala 169:30]
  wire  _GEN_7365 = uncached ? _GEN_2130 : _GEN_5814; // @[ICache.scala 169:30]
  wire  _GEN_7366 = uncached ? _GEN_2642 : _GEN_5815; // @[ICache.scala 169:30]
  wire  _GEN_7367 = uncached ? _GEN_2131 : _GEN_5816; // @[ICache.scala 169:30]
  wire  _GEN_7368 = uncached ? _GEN_2643 : _GEN_5817; // @[ICache.scala 169:30]
  wire  _GEN_7369 = uncached ? _GEN_2132 : _GEN_5818; // @[ICache.scala 169:30]
  wire  _GEN_7370 = uncached ? _GEN_2644 : _GEN_5819; // @[ICache.scala 169:30]
  wire  _GEN_7371 = uncached ? _GEN_2133 : _GEN_5820; // @[ICache.scala 169:30]
  wire  _GEN_7372 = uncached ? _GEN_2645 : _GEN_5821; // @[ICache.scala 169:30]
  wire  _GEN_7373 = uncached ? _GEN_2134 : _GEN_5822; // @[ICache.scala 169:30]
  wire  _GEN_7374 = uncached ? _GEN_2646 : _GEN_5823; // @[ICache.scala 169:30]
  wire  _GEN_7375 = uncached ? _GEN_2135 : _GEN_5824; // @[ICache.scala 169:30]
  wire  _GEN_7376 = uncached ? _GEN_2647 : _GEN_5825; // @[ICache.scala 169:30]
  wire  _GEN_7377 = uncached ? _GEN_2136 : _GEN_5826; // @[ICache.scala 169:30]
  wire  _GEN_7378 = uncached ? _GEN_2648 : _GEN_5827; // @[ICache.scala 169:30]
  wire  _GEN_7379 = uncached ? _GEN_2137 : _GEN_5828; // @[ICache.scala 169:30]
  wire  _GEN_7380 = uncached ? _GEN_2649 : _GEN_5829; // @[ICache.scala 169:30]
  wire  _GEN_7381 = uncached ? _GEN_2138 : _GEN_5830; // @[ICache.scala 169:30]
  wire  _GEN_7382 = uncached ? _GEN_2650 : _GEN_5831; // @[ICache.scala 169:30]
  wire  _GEN_7383 = uncached ? _GEN_2139 : _GEN_5832; // @[ICache.scala 169:30]
  wire  _GEN_7384 = uncached ? _GEN_2651 : _GEN_5833; // @[ICache.scala 169:30]
  wire  _GEN_7385 = uncached ? _GEN_2140 : _GEN_5834; // @[ICache.scala 169:30]
  wire  _GEN_7386 = uncached ? _GEN_2652 : _GEN_5835; // @[ICache.scala 169:30]
  wire  _GEN_7387 = uncached ? _GEN_2141 : _GEN_5836; // @[ICache.scala 169:30]
  wire  _GEN_7388 = uncached ? _GEN_2653 : _GEN_5837; // @[ICache.scala 169:30]
  wire  _GEN_7389 = uncached ? _GEN_2142 : _GEN_5838; // @[ICache.scala 169:30]
  wire  _GEN_7390 = uncached ? _GEN_2654 : _GEN_5839; // @[ICache.scala 169:30]
  wire  _GEN_7391 = uncached ? _GEN_2143 : _GEN_5840; // @[ICache.scala 169:30]
  wire  _GEN_7392 = uncached ? _GEN_2655 : _GEN_5841; // @[ICache.scala 169:30]
  wire  _GEN_7393 = uncached ? _GEN_2144 : _GEN_5842; // @[ICache.scala 169:30]
  wire  _GEN_7394 = uncached ? _GEN_2656 : _GEN_5843; // @[ICache.scala 169:30]
  wire  _GEN_7395 = uncached ? _GEN_2145 : _GEN_5844; // @[ICache.scala 169:30]
  wire  _GEN_7396 = uncached ? _GEN_2657 : _GEN_5845; // @[ICache.scala 169:30]
  wire  _GEN_7397 = uncached ? _GEN_2146 : _GEN_5846; // @[ICache.scala 169:30]
  wire  _GEN_7398 = uncached ? _GEN_2658 : _GEN_5847; // @[ICache.scala 169:30]
  wire  _GEN_7399 = uncached ? _GEN_2147 : _GEN_5848; // @[ICache.scala 169:30]
  wire  _GEN_7400 = uncached ? _GEN_2659 : _GEN_5849; // @[ICache.scala 169:30]
  wire  _GEN_7401 = uncached ? _GEN_2148 : _GEN_5850; // @[ICache.scala 169:30]
  wire  _GEN_7402 = uncached ? _GEN_2660 : _GEN_5851; // @[ICache.scala 169:30]
  wire  _GEN_7403 = uncached ? _GEN_2149 : _GEN_5852; // @[ICache.scala 169:30]
  wire  _GEN_7404 = uncached ? _GEN_2661 : _GEN_5853; // @[ICache.scala 169:30]
  wire  _GEN_7405 = uncached ? _GEN_2150 : _GEN_5854; // @[ICache.scala 169:30]
  wire  _GEN_7406 = uncached ? _GEN_2662 : _GEN_5855; // @[ICache.scala 169:30]
  wire  _GEN_7407 = uncached ? _GEN_2151 : _GEN_5856; // @[ICache.scala 169:30]
  wire  _GEN_7408 = uncached ? _GEN_2663 : _GEN_5857; // @[ICache.scala 169:30]
  wire  _GEN_7409 = uncached ? _GEN_2152 : _GEN_5858; // @[ICache.scala 169:30]
  wire  _GEN_7410 = uncached ? _GEN_2664 : _GEN_5859; // @[ICache.scala 169:30]
  wire  _GEN_7411 = uncached ? _GEN_2153 : _GEN_5860; // @[ICache.scala 169:30]
  wire  _GEN_7412 = uncached ? _GEN_2665 : _GEN_5861; // @[ICache.scala 169:30]
  wire  _GEN_7413 = uncached ? _GEN_2154 : _GEN_5862; // @[ICache.scala 169:30]
  wire  _GEN_7414 = uncached ? _GEN_2666 : _GEN_5863; // @[ICache.scala 169:30]
  wire  _GEN_7415 = uncached ? _GEN_2155 : _GEN_5864; // @[ICache.scala 169:30]
  wire  _GEN_7416 = uncached ? _GEN_2667 : _GEN_5865; // @[ICache.scala 169:30]
  wire  _GEN_7417 = uncached ? _GEN_2156 : _GEN_5866; // @[ICache.scala 169:30]
  wire  _GEN_7418 = uncached ? _GEN_2668 : _GEN_5867; // @[ICache.scala 169:30]
  wire  _GEN_7419 = uncached ? _GEN_2157 : _GEN_5868; // @[ICache.scala 169:30]
  wire  _GEN_7420 = uncached ? _GEN_2669 : _GEN_5869; // @[ICache.scala 169:30]
  wire  _GEN_7421 = uncached ? _GEN_2158 : _GEN_5870; // @[ICache.scala 169:30]
  wire  _GEN_7422 = uncached ? _GEN_2670 : _GEN_5871; // @[ICache.scala 169:30]
  wire  _GEN_7423 = uncached ? _GEN_2159 : _GEN_5872; // @[ICache.scala 169:30]
  wire  _GEN_7424 = uncached ? _GEN_2671 : _GEN_5873; // @[ICache.scala 169:30]
  wire  _GEN_7425 = uncached ? _GEN_2160 : _GEN_5874; // @[ICache.scala 169:30]
  wire  _GEN_7426 = uncached ? _GEN_2672 : _GEN_5875; // @[ICache.scala 169:30]
  wire  _GEN_7427 = uncached ? _GEN_2161 : _GEN_5876; // @[ICache.scala 169:30]
  wire  _GEN_7428 = uncached ? _GEN_2673 : _GEN_5877; // @[ICache.scala 169:30]
  wire  _GEN_7429 = uncached ? _GEN_2162 : _GEN_5878; // @[ICache.scala 169:30]
  wire  _GEN_7430 = uncached ? _GEN_2674 : _GEN_5879; // @[ICache.scala 169:30]
  wire  _GEN_7431 = uncached ? _GEN_2163 : _GEN_5880; // @[ICache.scala 169:30]
  wire  _GEN_7432 = uncached ? _GEN_2675 : _GEN_5881; // @[ICache.scala 169:30]
  wire  _GEN_7433 = uncached ? _GEN_2164 : _GEN_5882; // @[ICache.scala 169:30]
  wire  _GEN_7434 = uncached ? _GEN_2676 : _GEN_5883; // @[ICache.scala 169:30]
  wire  _GEN_7435 = uncached ? _GEN_2165 : _GEN_5884; // @[ICache.scala 169:30]
  wire  _GEN_7436 = uncached ? _GEN_2677 : _GEN_5885; // @[ICache.scala 169:30]
  wire  _GEN_7437 = uncached ? _GEN_2166 : _GEN_5886; // @[ICache.scala 169:30]
  wire  _GEN_7438 = uncached ? _GEN_2678 : _GEN_5887; // @[ICache.scala 169:30]
  wire  _GEN_7439 = uncached ? _GEN_2167 : _GEN_5888; // @[ICache.scala 169:30]
  wire  _GEN_7440 = uncached ? _GEN_2679 : _GEN_5889; // @[ICache.scala 169:30]
  wire  _GEN_7441 = uncached ? _GEN_2168 : _GEN_5890; // @[ICache.scala 169:30]
  wire  _GEN_7442 = uncached ? _GEN_2680 : _GEN_5891; // @[ICache.scala 169:30]
  wire  _GEN_7443 = uncached ? _GEN_2169 : _GEN_5892; // @[ICache.scala 169:30]
  wire  _GEN_7444 = uncached ? _GEN_2681 : _GEN_5893; // @[ICache.scala 169:30]
  wire  _GEN_7445 = uncached ? _GEN_2170 : _GEN_5894; // @[ICache.scala 169:30]
  wire  _GEN_7446 = uncached ? _GEN_2682 : _GEN_5895; // @[ICache.scala 169:30]
  wire  _GEN_7447 = uncached ? _GEN_2171 : _GEN_5896; // @[ICache.scala 169:30]
  wire  _GEN_7448 = uncached ? _GEN_2683 : _GEN_5897; // @[ICache.scala 169:30]
  wire  _GEN_7449 = uncached ? _GEN_2172 : _GEN_5898; // @[ICache.scala 169:30]
  wire  _GEN_7450 = uncached ? _GEN_2684 : _GEN_5899; // @[ICache.scala 169:30]
  wire  _GEN_7451 = uncached ? _GEN_2173 : _GEN_5900; // @[ICache.scala 169:30]
  wire  _GEN_7452 = uncached ? _GEN_2685 : _GEN_5901; // @[ICache.scala 169:30]
  wire  _GEN_7453 = uncached ? _GEN_2174 : _GEN_5902; // @[ICache.scala 169:30]
  wire  _GEN_7454 = uncached ? _GEN_2686 : _GEN_5903; // @[ICache.scala 169:30]
  wire  _GEN_7455 = uncached ? _GEN_2175 : _GEN_5904; // @[ICache.scala 169:30]
  wire  _GEN_7456 = uncached ? _GEN_2687 : _GEN_5905; // @[ICache.scala 169:30]
  wire  _GEN_7457 = uncached ? _GEN_2176 : _GEN_5906; // @[ICache.scala 169:30]
  wire  _GEN_7458 = uncached ? _GEN_2688 : _GEN_5907; // @[ICache.scala 169:30]
  wire  _GEN_7459 = uncached ? _GEN_2177 : _GEN_5908; // @[ICache.scala 169:30]
  wire  _GEN_7460 = uncached ? _GEN_2689 : _GEN_5909; // @[ICache.scala 169:30]
  wire  _GEN_7461 = uncached ? _GEN_2178 : _GEN_5910; // @[ICache.scala 169:30]
  wire  _GEN_7462 = uncached ? _GEN_2690 : _GEN_5911; // @[ICache.scala 169:30]
  wire  _GEN_7463 = uncached ? _GEN_2179 : _GEN_5912; // @[ICache.scala 169:30]
  wire  _GEN_7464 = uncached ? _GEN_2691 : _GEN_5913; // @[ICache.scala 169:30]
  wire  _GEN_7465 = uncached ? _GEN_2180 : _GEN_5914; // @[ICache.scala 169:30]
  wire  _GEN_7466 = uncached ? _GEN_2692 : _GEN_5915; // @[ICache.scala 169:30]
  wire  _GEN_7467 = uncached ? _GEN_2181 : _GEN_5916; // @[ICache.scala 169:30]
  wire  _GEN_7468 = uncached ? _GEN_2693 : _GEN_5917; // @[ICache.scala 169:30]
  wire  _GEN_7469 = uncached ? _GEN_2182 : _GEN_5918; // @[ICache.scala 169:30]
  wire  _GEN_7470 = uncached ? _GEN_2694 : _GEN_5919; // @[ICache.scala 169:30]
  wire  _GEN_7471 = uncached ? _GEN_2183 : _GEN_5920; // @[ICache.scala 169:30]
  wire  _GEN_7472 = uncached ? _GEN_2695 : _GEN_5921; // @[ICache.scala 169:30]
  wire  _GEN_7473 = uncached ? _GEN_2184 : _GEN_5922; // @[ICache.scala 169:30]
  wire  _GEN_7474 = uncached ? _GEN_2696 : _GEN_5923; // @[ICache.scala 169:30]
  wire  _GEN_7475 = uncached ? _GEN_2185 : _GEN_5924; // @[ICache.scala 169:30]
  wire  _GEN_7476 = uncached ? _GEN_2697 : _GEN_5925; // @[ICache.scala 169:30]
  wire  _GEN_7477 = uncached ? _GEN_2186 : _GEN_5926; // @[ICache.scala 169:30]
  wire  _GEN_7478 = uncached ? _GEN_2698 : _GEN_5927; // @[ICache.scala 169:30]
  wire  _GEN_7479 = uncached ? _GEN_2187 : _GEN_5928; // @[ICache.scala 169:30]
  wire  _GEN_7480 = uncached ? _GEN_2699 : _GEN_5929; // @[ICache.scala 169:30]
  wire  _GEN_7481 = uncached ? _GEN_2188 : _GEN_5930; // @[ICache.scala 169:30]
  wire  _GEN_7482 = uncached ? _GEN_2700 : _GEN_5931; // @[ICache.scala 169:30]
  wire  _GEN_7483 = uncached ? _GEN_2189 : _GEN_5932; // @[ICache.scala 169:30]
  wire  _GEN_7484 = uncached ? _GEN_2701 : _GEN_5933; // @[ICache.scala 169:30]
  wire  _GEN_7485 = uncached ? _GEN_2190 : _GEN_5934; // @[ICache.scala 169:30]
  wire  _GEN_7486 = uncached ? _GEN_2702 : _GEN_5935; // @[ICache.scala 169:30]
  wire  _GEN_7487 = uncached ? _GEN_2191 : _GEN_5936; // @[ICache.scala 169:30]
  wire  _GEN_7488 = uncached ? _GEN_2703 : _GEN_5937; // @[ICache.scala 169:30]
  wire  _GEN_7489 = uncached ? _GEN_2192 : _GEN_5938; // @[ICache.scala 169:30]
  wire  _GEN_7490 = uncached ? _GEN_2704 : _GEN_5939; // @[ICache.scala 169:30]
  wire  _GEN_7491 = uncached ? _GEN_2193 : _GEN_5940; // @[ICache.scala 169:30]
  wire  _GEN_7492 = uncached ? _GEN_2705 : _GEN_5941; // @[ICache.scala 169:30]
  wire  _GEN_7493 = uncached ? _GEN_2194 : _GEN_5942; // @[ICache.scala 169:30]
  wire  _GEN_7494 = uncached ? _GEN_2706 : _GEN_5943; // @[ICache.scala 169:30]
  wire  _GEN_7495 = uncached ? _GEN_2195 : _GEN_5944; // @[ICache.scala 169:30]
  wire  _GEN_7496 = uncached ? _GEN_2707 : _GEN_5945; // @[ICache.scala 169:30]
  wire  _GEN_7497 = uncached ? _GEN_2196 : _GEN_5946; // @[ICache.scala 169:30]
  wire  _GEN_7498 = uncached ? _GEN_2708 : _GEN_5947; // @[ICache.scala 169:30]
  wire  _GEN_7499 = uncached ? _GEN_2197 : _GEN_5948; // @[ICache.scala 169:30]
  wire  _GEN_7500 = uncached ? _GEN_2709 : _GEN_5949; // @[ICache.scala 169:30]
  wire  _GEN_7501 = uncached ? _GEN_2198 : _GEN_5950; // @[ICache.scala 169:30]
  wire  _GEN_7502 = uncached ? _GEN_2710 : _GEN_5951; // @[ICache.scala 169:30]
  wire  _GEN_7503 = uncached ? _GEN_2199 : _GEN_5952; // @[ICache.scala 169:30]
  wire  _GEN_7504 = uncached ? _GEN_2711 : _GEN_5953; // @[ICache.scala 169:30]
  wire  _GEN_7505 = uncached ? _GEN_2200 : _GEN_5954; // @[ICache.scala 169:30]
  wire  _GEN_7506 = uncached ? _GEN_2712 : _GEN_5955; // @[ICache.scala 169:30]
  wire  _GEN_7507 = uncached ? _GEN_2201 : _GEN_5956; // @[ICache.scala 169:30]
  wire  _GEN_7508 = uncached ? _GEN_2713 : _GEN_5957; // @[ICache.scala 169:30]
  wire  _GEN_7509 = uncached ? _GEN_2202 : _GEN_5958; // @[ICache.scala 169:30]
  wire  _GEN_7510 = uncached ? _GEN_2714 : _GEN_5959; // @[ICache.scala 169:30]
  wire  _GEN_7511 = uncached ? _GEN_2203 : _GEN_5960; // @[ICache.scala 169:30]
  wire  _GEN_7512 = uncached ? _GEN_2715 : _GEN_5961; // @[ICache.scala 169:30]
  wire  _GEN_7513 = uncached ? _GEN_2204 : _GEN_5962; // @[ICache.scala 169:30]
  wire  _GEN_7514 = uncached ? _GEN_2716 : _GEN_5963; // @[ICache.scala 169:30]
  wire  _GEN_7515 = uncached ? _GEN_2205 : _GEN_5964; // @[ICache.scala 169:30]
  wire  _GEN_7516 = uncached ? _GEN_2717 : _GEN_5965; // @[ICache.scala 169:30]
  wire  _GEN_7517 = uncached ? _GEN_2206 : _GEN_5966; // @[ICache.scala 169:30]
  wire  _GEN_7518 = uncached ? _GEN_2718 : _GEN_5967; // @[ICache.scala 169:30]
  wire  _GEN_7519 = uncached ? _GEN_2207 : _GEN_5968; // @[ICache.scala 169:30]
  wire  _GEN_7520 = uncached ? _GEN_2719 : _GEN_5969; // @[ICache.scala 169:30]
  wire  _GEN_7521 = uncached ? _GEN_2208 : _GEN_5970; // @[ICache.scala 169:30]
  wire  _GEN_7522 = uncached ? _GEN_2720 : _GEN_5971; // @[ICache.scala 169:30]
  wire  _GEN_7523 = uncached ? _GEN_2209 : _GEN_5972; // @[ICache.scala 169:30]
  wire  _GEN_7524 = uncached ? _GEN_2721 : _GEN_5973; // @[ICache.scala 169:30]
  wire  _GEN_7525 = uncached ? _GEN_2210 : _GEN_5974; // @[ICache.scala 169:30]
  wire  _GEN_7526 = uncached ? _GEN_2722 : _GEN_5975; // @[ICache.scala 169:30]
  wire  _GEN_7527 = uncached ? _GEN_2211 : _GEN_5976; // @[ICache.scala 169:30]
  wire  _GEN_7528 = uncached ? _GEN_2723 : _GEN_5977; // @[ICache.scala 169:30]
  wire  _GEN_7529 = uncached ? _GEN_2212 : _GEN_5978; // @[ICache.scala 169:30]
  wire  _GEN_7530 = uncached ? _GEN_2724 : _GEN_5979; // @[ICache.scala 169:30]
  wire  _GEN_7531 = uncached ? _GEN_2213 : _GEN_5980; // @[ICache.scala 169:30]
  wire  _GEN_7532 = uncached ? _GEN_2725 : _GEN_5981; // @[ICache.scala 169:30]
  wire  _GEN_7533 = uncached ? _GEN_2214 : _GEN_5982; // @[ICache.scala 169:30]
  wire  _GEN_7534 = uncached ? _GEN_2726 : _GEN_5983; // @[ICache.scala 169:30]
  wire  _GEN_7535 = uncached ? _GEN_2215 : _GEN_5984; // @[ICache.scala 169:30]
  wire  _GEN_7536 = uncached ? _GEN_2727 : _GEN_5985; // @[ICache.scala 169:30]
  wire  _GEN_7537 = uncached ? _GEN_2216 : _GEN_5986; // @[ICache.scala 169:30]
  wire  _GEN_7538 = uncached ? _GEN_2728 : _GEN_5987; // @[ICache.scala 169:30]
  wire  _GEN_7539 = uncached ? _GEN_2217 : _GEN_5988; // @[ICache.scala 169:30]
  wire  _GEN_7540 = uncached ? _GEN_2729 : _GEN_5989; // @[ICache.scala 169:30]
  wire  _GEN_7541 = uncached ? _GEN_2218 : _GEN_5990; // @[ICache.scala 169:30]
  wire  _GEN_7542 = uncached ? _GEN_2730 : _GEN_5991; // @[ICache.scala 169:30]
  wire  _GEN_7543 = uncached ? _GEN_2219 : _GEN_5992; // @[ICache.scala 169:30]
  wire  _GEN_7544 = uncached ? _GEN_2731 : _GEN_5993; // @[ICache.scala 169:30]
  wire  _GEN_7545 = uncached ? _GEN_2220 : _GEN_5994; // @[ICache.scala 169:30]
  wire  _GEN_7546 = uncached ? _GEN_2732 : _GEN_5995; // @[ICache.scala 169:30]
  wire  _GEN_7547 = uncached ? _GEN_2221 : _GEN_5996; // @[ICache.scala 169:30]
  wire  _GEN_7548 = uncached ? _GEN_2733 : _GEN_5997; // @[ICache.scala 169:30]
  wire  _GEN_7549 = uncached ? _GEN_2222 : _GEN_5998; // @[ICache.scala 169:30]
  wire  _GEN_7550 = uncached ? _GEN_2734 : _GEN_5999; // @[ICache.scala 169:30]
  wire  _GEN_7551 = uncached ? _GEN_2223 : _GEN_6000; // @[ICache.scala 169:30]
  wire  _GEN_7552 = uncached ? _GEN_2735 : _GEN_6001; // @[ICache.scala 169:30]
  wire  _GEN_7553 = uncached ? _GEN_2224 : _GEN_6002; // @[ICache.scala 169:30]
  wire  _GEN_7554 = uncached ? _GEN_2736 : _GEN_6003; // @[ICache.scala 169:30]
  wire  _GEN_7555 = uncached ? _GEN_2225 : _GEN_6004; // @[ICache.scala 169:30]
  wire  _GEN_7556 = uncached ? _GEN_2737 : _GEN_6005; // @[ICache.scala 169:30]
  wire  _GEN_7557 = uncached ? _GEN_2226 : _GEN_6006; // @[ICache.scala 169:30]
  wire  _GEN_7558 = uncached ? _GEN_2738 : _GEN_6007; // @[ICache.scala 169:30]
  wire  _GEN_7559 = uncached ? _GEN_2227 : _GEN_6008; // @[ICache.scala 169:30]
  wire  _GEN_7560 = uncached ? _GEN_2739 : _GEN_6009; // @[ICache.scala 169:30]
  wire  _GEN_7561 = uncached ? _GEN_2228 : _GEN_6010; // @[ICache.scala 169:30]
  wire  _GEN_7562 = uncached ? _GEN_2740 : _GEN_6011; // @[ICache.scala 169:30]
  wire  _GEN_7563 = uncached ? _GEN_2229 : _GEN_6012; // @[ICache.scala 169:30]
  wire  _GEN_7564 = uncached ? _GEN_2741 : _GEN_6013; // @[ICache.scala 169:30]
  wire  _GEN_7565 = uncached ? _GEN_2230 : _GEN_6014; // @[ICache.scala 169:30]
  wire  _GEN_7566 = uncached ? _GEN_2742 : _GEN_6015; // @[ICache.scala 169:30]
  wire  _GEN_7567 = uncached ? _GEN_2231 : _GEN_6016; // @[ICache.scala 169:30]
  wire  _GEN_7568 = uncached ? _GEN_2743 : _GEN_6017; // @[ICache.scala 169:30]
  wire  _GEN_7569 = uncached ? _GEN_2232 : _GEN_6018; // @[ICache.scala 169:30]
  wire  _GEN_7570 = uncached ? _GEN_2744 : _GEN_6019; // @[ICache.scala 169:30]
  wire  _GEN_7571 = uncached ? _GEN_2233 : _GEN_6020; // @[ICache.scala 169:30]
  wire  _GEN_7572 = uncached ? _GEN_2745 : _GEN_6021; // @[ICache.scala 169:30]
  wire  _GEN_7573 = uncached ? _GEN_2234 : _GEN_6022; // @[ICache.scala 169:30]
  wire  _GEN_7574 = uncached ? _GEN_2746 : _GEN_6023; // @[ICache.scala 169:30]
  wire  _GEN_7575 = uncached ? _GEN_2235 : _GEN_6024; // @[ICache.scala 169:30]
  wire  _GEN_7576 = uncached ? _GEN_2747 : _GEN_6025; // @[ICache.scala 169:30]
  wire  _GEN_7577 = uncached ? _GEN_2236 : _GEN_6026; // @[ICache.scala 169:30]
  wire  _GEN_7578 = uncached ? _GEN_2748 : _GEN_6027; // @[ICache.scala 169:30]
  wire  _GEN_7579 = uncached ? _GEN_2237 : _GEN_6028; // @[ICache.scala 169:30]
  wire  _GEN_7580 = uncached ? _GEN_2749 : _GEN_6029; // @[ICache.scala 169:30]
  wire  _GEN_7581 = uncached ? _GEN_2238 : _GEN_6030; // @[ICache.scala 169:30]
  wire  _GEN_7582 = uncached ? _GEN_2750 : _GEN_6031; // @[ICache.scala 169:30]
  wire  _GEN_7583 = uncached ? _GEN_2239 : _GEN_6032; // @[ICache.scala 169:30]
  wire  _GEN_7584 = uncached ? _GEN_2751 : _GEN_6033; // @[ICache.scala 169:30]
  wire  _GEN_7585 = uncached ? _GEN_2240 : _GEN_6034; // @[ICache.scala 169:30]
  wire  _GEN_7586 = uncached ? _GEN_2752 : _GEN_6035; // @[ICache.scala 169:30]
  wire  _GEN_7587 = uncached ? _GEN_2241 : _GEN_6036; // @[ICache.scala 169:30]
  wire  _GEN_7588 = uncached ? _GEN_2753 : _GEN_6037; // @[ICache.scala 169:30]
  wire  _GEN_7589 = uncached ? _GEN_2242 : _GEN_6038; // @[ICache.scala 169:30]
  wire  _GEN_7590 = uncached ? _GEN_2754 : _GEN_6039; // @[ICache.scala 169:30]
  wire  _GEN_7591 = uncached ? _GEN_2243 : _GEN_6040; // @[ICache.scala 169:30]
  wire  _GEN_7592 = uncached ? _GEN_2755 : _GEN_6041; // @[ICache.scala 169:30]
  wire  _GEN_7593 = uncached ? _GEN_2244 : _GEN_6042; // @[ICache.scala 169:30]
  wire  _GEN_7594 = uncached ? _GEN_2756 : _GEN_6043; // @[ICache.scala 169:30]
  wire  _GEN_7595 = uncached ? _GEN_2245 : _GEN_6044; // @[ICache.scala 169:30]
  wire  _GEN_7596 = uncached ? _GEN_2757 : _GEN_6045; // @[ICache.scala 169:30]
  wire  _GEN_7597 = uncached ? _GEN_2246 : _GEN_6046; // @[ICache.scala 169:30]
  wire  _GEN_7598 = uncached ? _GEN_2758 : _GEN_6047; // @[ICache.scala 169:30]
  wire  _GEN_7599 = uncached ? _GEN_2247 : _GEN_6048; // @[ICache.scala 169:30]
  wire  _GEN_7600 = uncached ? _GEN_2759 : _GEN_6049; // @[ICache.scala 169:30]
  wire  _GEN_7601 = uncached ? _GEN_2248 : _GEN_6050; // @[ICache.scala 169:30]
  wire  _GEN_7602 = uncached ? _GEN_2760 : _GEN_6051; // @[ICache.scala 169:30]
  wire  _GEN_7603 = uncached ? _GEN_2249 : _GEN_6052; // @[ICache.scala 169:30]
  wire  _GEN_7604 = uncached ? _GEN_2761 : _GEN_6053; // @[ICache.scala 169:30]
  wire  _GEN_7605 = uncached ? _GEN_2250 : _GEN_6054; // @[ICache.scala 169:30]
  wire  _GEN_7606 = uncached ? _GEN_2762 : _GEN_6055; // @[ICache.scala 169:30]
  wire  _GEN_7607 = uncached ? _GEN_2251 : _GEN_6056; // @[ICache.scala 169:30]
  wire  _GEN_7608 = uncached ? _GEN_2763 : _GEN_6057; // @[ICache.scala 169:30]
  wire  _GEN_7609 = uncached ? _GEN_2252 : _GEN_6058; // @[ICache.scala 169:30]
  wire  _GEN_7610 = uncached ? _GEN_2764 : _GEN_6059; // @[ICache.scala 169:30]
  wire  _GEN_7611 = uncached ? _GEN_2253 : _GEN_6060; // @[ICache.scala 169:30]
  wire  _GEN_7612 = uncached ? _GEN_2765 : _GEN_6061; // @[ICache.scala 169:30]
  wire  _GEN_7613 = uncached ? _GEN_2254 : _GEN_6062; // @[ICache.scala 169:30]
  wire  _GEN_7614 = uncached ? _GEN_2766 : _GEN_6063; // @[ICache.scala 169:30]
  wire  _GEN_7615 = uncached ? _GEN_2255 : _GEN_6064; // @[ICache.scala 169:30]
  wire  _GEN_7616 = uncached ? _GEN_2767 : _GEN_6065; // @[ICache.scala 169:30]
  wire  _GEN_7617 = uncached ? _GEN_2256 : _GEN_6066; // @[ICache.scala 169:30]
  wire  _GEN_7618 = uncached ? _GEN_2768 : _GEN_6067; // @[ICache.scala 169:30]
  wire  _GEN_7619 = uncached ? _GEN_2257 : _GEN_6068; // @[ICache.scala 169:30]
  wire  _GEN_7620 = uncached ? _GEN_2769 : _GEN_6069; // @[ICache.scala 169:30]
  wire  _GEN_7621 = uncached ? _GEN_2258 : _GEN_6070; // @[ICache.scala 169:30]
  wire  _GEN_7622 = uncached ? _GEN_2770 : _GEN_6071; // @[ICache.scala 169:30]
  wire  _GEN_7623 = uncached ? _GEN_2259 : _GEN_6072; // @[ICache.scala 169:30]
  wire  _GEN_7624 = uncached ? _GEN_2771 : _GEN_6073; // @[ICache.scala 169:30]
  wire  _GEN_7625 = uncached ? _GEN_2260 : _GEN_6074; // @[ICache.scala 169:30]
  wire  _GEN_7626 = uncached ? _GEN_2772 : _GEN_6075; // @[ICache.scala 169:30]
  wire  _GEN_7627 = uncached ? _GEN_2261 : _GEN_6076; // @[ICache.scala 169:30]
  wire  _GEN_7628 = uncached ? _GEN_2773 : _GEN_6077; // @[ICache.scala 169:30]
  wire  _GEN_7629 = uncached ? _GEN_2262 : _GEN_6078; // @[ICache.scala 169:30]
  wire  _GEN_7630 = uncached ? _GEN_2774 : _GEN_6079; // @[ICache.scala 169:30]
  wire  _GEN_7631 = uncached ? _GEN_2263 : _GEN_6080; // @[ICache.scala 169:30]
  wire  _GEN_7632 = uncached ? _GEN_2775 : _GEN_6081; // @[ICache.scala 169:30]
  wire  _GEN_7633 = uncached ? _GEN_2264 : _GEN_6082; // @[ICache.scala 169:30]
  wire  _GEN_7634 = uncached ? _GEN_2776 : _GEN_6083; // @[ICache.scala 169:30]
  wire  _GEN_7635 = uncached ? _GEN_2265 : _GEN_6084; // @[ICache.scala 169:30]
  wire  _GEN_7636 = uncached ? _GEN_2777 : _GEN_6085; // @[ICache.scala 169:30]
  wire  _GEN_7637 = uncached ? _GEN_2266 : _GEN_6086; // @[ICache.scala 169:30]
  wire  _GEN_7638 = uncached ? _GEN_2778 : _GEN_6087; // @[ICache.scala 169:30]
  wire  _GEN_7639 = uncached ? _GEN_2267 : _GEN_6088; // @[ICache.scala 169:30]
  wire  _GEN_7640 = uncached ? _GEN_2779 : _GEN_6089; // @[ICache.scala 169:30]
  wire  _GEN_7641 = uncached ? _GEN_2268 : _GEN_6090; // @[ICache.scala 169:30]
  wire  _GEN_7642 = uncached ? _GEN_2780 : _GEN_6091; // @[ICache.scala 169:30]
  wire  _GEN_7643 = uncached ? _GEN_2269 : _GEN_6092; // @[ICache.scala 169:30]
  wire  _GEN_7644 = uncached ? _GEN_2781 : _GEN_6093; // @[ICache.scala 169:30]
  wire  _GEN_7645 = uncached ? _GEN_2270 : _GEN_6094; // @[ICache.scala 169:30]
  wire  _GEN_7646 = uncached ? _GEN_2782 : _GEN_6095; // @[ICache.scala 169:30]
  wire  _GEN_7647 = uncached ? _GEN_2271 : _GEN_6096; // @[ICache.scala 169:30]
  wire  _GEN_7648 = uncached ? _GEN_2783 : _GEN_6097; // @[ICache.scala 169:30]
  wire  _GEN_7649 = uncached ? _GEN_2272 : _GEN_6098; // @[ICache.scala 169:30]
  wire  _GEN_7650 = uncached ? _GEN_2784 : _GEN_6099; // @[ICache.scala 169:30]
  wire  _GEN_7651 = uncached ? _GEN_2273 : _GEN_6100; // @[ICache.scala 169:30]
  wire  _GEN_7652 = uncached ? _GEN_2785 : _GEN_6101; // @[ICache.scala 169:30]
  wire  _GEN_7653 = uncached ? _GEN_2274 : _GEN_6102; // @[ICache.scala 169:30]
  wire  _GEN_7654 = uncached ? _GEN_2786 : _GEN_6103; // @[ICache.scala 169:30]
  wire  _GEN_7655 = uncached ? _GEN_2275 : _GEN_6104; // @[ICache.scala 169:30]
  wire  _GEN_7656 = uncached ? _GEN_2787 : _GEN_6105; // @[ICache.scala 169:30]
  wire  _GEN_7657 = uncached ? _GEN_2276 : _GEN_6106; // @[ICache.scala 169:30]
  wire  _GEN_7658 = uncached ? _GEN_2788 : _GEN_6107; // @[ICache.scala 169:30]
  wire  _GEN_7659 = uncached ? _GEN_2277 : _GEN_6108; // @[ICache.scala 169:30]
  wire  _GEN_7660 = uncached ? _GEN_2789 : _GEN_6109; // @[ICache.scala 169:30]
  wire  _GEN_7661 = uncached ? _GEN_2278 : _GEN_6110; // @[ICache.scala 169:30]
  wire  _GEN_7662 = uncached ? _GEN_2790 : _GEN_6111; // @[ICache.scala 169:30]
  wire  _GEN_7663 = uncached ? _GEN_2279 : _GEN_6112; // @[ICache.scala 169:30]
  wire  _GEN_7664 = uncached ? _GEN_2791 : _GEN_6113; // @[ICache.scala 169:30]
  wire  _GEN_7665 = uncached ? _GEN_2280 : _GEN_6114; // @[ICache.scala 169:30]
  wire  _GEN_7666 = uncached ? _GEN_2792 : _GEN_6115; // @[ICache.scala 169:30]
  wire  _GEN_7667 = uncached ? _GEN_2281 : _GEN_6116; // @[ICache.scala 169:30]
  wire  _GEN_7668 = uncached ? _GEN_2793 : _GEN_6117; // @[ICache.scala 169:30]
  wire  _GEN_7669 = uncached ? _GEN_2282 : _GEN_6118; // @[ICache.scala 169:30]
  wire  _GEN_7670 = uncached ? _GEN_2794 : _GEN_6119; // @[ICache.scala 169:30]
  wire  _GEN_7671 = uncached ? _GEN_2283 : _GEN_6120; // @[ICache.scala 169:30]
  wire  _GEN_7672 = uncached ? _GEN_2795 : _GEN_6121; // @[ICache.scala 169:30]
  wire  _GEN_7673 = uncached ? _GEN_2284 : _GEN_6122; // @[ICache.scala 169:30]
  wire  _GEN_7674 = uncached ? _GEN_2796 : _GEN_6123; // @[ICache.scala 169:30]
  wire  _GEN_7675 = uncached ? _GEN_2285 : _GEN_6124; // @[ICache.scala 169:30]
  wire  _GEN_7676 = uncached ? _GEN_2797 : _GEN_6125; // @[ICache.scala 169:30]
  wire  _GEN_7677 = uncached ? _GEN_2286 : _GEN_6126; // @[ICache.scala 169:30]
  wire  _GEN_7678 = uncached ? _GEN_2798 : _GEN_6127; // @[ICache.scala 169:30]
  wire  _GEN_7679 = uncached ? _GEN_2287 : _GEN_6128; // @[ICache.scala 169:30]
  wire  _GEN_7680 = uncached ? _GEN_2799 : _GEN_6129; // @[ICache.scala 169:30]
  wire  _GEN_7681 = uncached ? _GEN_2288 : _GEN_6130; // @[ICache.scala 169:30]
  wire  _GEN_7682 = uncached ? _GEN_2800 : _GEN_6131; // @[ICache.scala 169:30]
  wire  _GEN_7683 = uncached ? _GEN_2289 : _GEN_6132; // @[ICache.scala 169:30]
  wire  _GEN_7684 = uncached ? _GEN_2801 : _GEN_6133; // @[ICache.scala 169:30]
  wire  _GEN_7685 = uncached ? _GEN_2290 : _GEN_6134; // @[ICache.scala 169:30]
  wire  _GEN_7686 = uncached ? _GEN_2802 : _GEN_6135; // @[ICache.scala 169:30]
  wire  _GEN_7687 = uncached ? _GEN_2291 : _GEN_6136; // @[ICache.scala 169:30]
  wire  _GEN_7688 = uncached ? _GEN_2803 : _GEN_6137; // @[ICache.scala 169:30]
  wire  _GEN_7689 = uncached ? _GEN_2292 : _GEN_6138; // @[ICache.scala 169:30]
  wire  _GEN_7690 = uncached ? _GEN_2804 : _GEN_6139; // @[ICache.scala 169:30]
  wire  _GEN_7691 = uncached ? _GEN_2293 : _GEN_6140; // @[ICache.scala 169:30]
  wire  _GEN_7692 = uncached ? _GEN_2805 : _GEN_6141; // @[ICache.scala 169:30]
  wire  _GEN_7693 = uncached ? _GEN_2294 : _GEN_6142; // @[ICache.scala 169:30]
  wire  _GEN_7694 = uncached ? _GEN_2806 : _GEN_6143; // @[ICache.scala 169:30]
  wire  _GEN_7695 = uncached ? _GEN_2295 : _GEN_6144; // @[ICache.scala 169:30]
  wire  _GEN_7696 = uncached ? _GEN_2807 : _GEN_6145; // @[ICache.scala 169:30]
  wire  _GEN_7697 = uncached ? _GEN_2296 : _GEN_6146; // @[ICache.scala 169:30]
  wire  _GEN_7698 = uncached ? _GEN_2808 : _GEN_6147; // @[ICache.scala 169:30]
  wire  _GEN_7699 = uncached ? _GEN_2297 : _GEN_6148; // @[ICache.scala 169:30]
  wire  _GEN_7700 = uncached ? _GEN_2809 : _GEN_6149; // @[ICache.scala 169:30]
  wire  _GEN_7701 = uncached ? _GEN_2298 : _GEN_6150; // @[ICache.scala 169:30]
  wire  _GEN_7702 = uncached ? _GEN_2810 : _GEN_6151; // @[ICache.scala 169:30]
  wire  _GEN_7703 = uncached ? _GEN_2299 : _GEN_6152; // @[ICache.scala 169:30]
  wire  _GEN_7704 = uncached ? _GEN_2811 : _GEN_6153; // @[ICache.scala 169:30]
  wire  _GEN_7705 = uncached ? _GEN_2300 : _GEN_6154; // @[ICache.scala 169:30]
  wire  _GEN_7706 = uncached ? _GEN_2812 : _GEN_6155; // @[ICache.scala 169:30]
  wire  _GEN_7707 = uncached ? _GEN_2301 : _GEN_6156; // @[ICache.scala 169:30]
  wire  _GEN_7708 = uncached ? _GEN_2813 : _GEN_6157; // @[ICache.scala 169:30]
  wire  _GEN_7709 = uncached ? _GEN_2302 : _GEN_6158; // @[ICache.scala 169:30]
  wire  _GEN_7710 = uncached ? _GEN_2814 : _GEN_6159; // @[ICache.scala 169:30]
  wire  _GEN_7711 = uncached ? _GEN_2303 : _GEN_6160; // @[ICache.scala 169:30]
  wire  _GEN_7712 = uncached ? _GEN_2815 : _GEN_6161; // @[ICache.scala 169:30]
  wire  _GEN_7713 = uncached ? _GEN_2304 : _GEN_6162; // @[ICache.scala 169:30]
  wire  _GEN_7714 = uncached ? _GEN_2816 : _GEN_6163; // @[ICache.scala 169:30]
  wire  _GEN_7715 = uncached ? _GEN_2305 : _GEN_6164; // @[ICache.scala 169:30]
  wire  _GEN_7716 = uncached ? _GEN_2817 : _GEN_6165; // @[ICache.scala 169:30]
  wire  _GEN_7717 = uncached ? _GEN_2306 : _GEN_6166; // @[ICache.scala 169:30]
  wire  _GEN_7718 = uncached ? _GEN_2818 : _GEN_6167; // @[ICache.scala 169:30]
  wire  _GEN_7719 = uncached ? _GEN_2307 : _GEN_6168; // @[ICache.scala 169:30]
  wire  _GEN_7720 = uncached ? _GEN_2819 : _GEN_6169; // @[ICache.scala 169:30]
  wire  _GEN_7721 = uncached ? _GEN_2308 : _GEN_6170; // @[ICache.scala 169:30]
  wire  _GEN_7722 = uncached ? _GEN_2820 : _GEN_6171; // @[ICache.scala 169:30]
  wire  _GEN_7723 = uncached ? _GEN_2309 : _GEN_6172; // @[ICache.scala 169:30]
  wire  _GEN_7724 = uncached ? _GEN_2821 : _GEN_6173; // @[ICache.scala 169:30]
  wire  _GEN_7725 = uncached ? _GEN_2310 : _GEN_6174; // @[ICache.scala 169:30]
  wire  _GEN_7726 = uncached ? _GEN_2822 : _GEN_6175; // @[ICache.scala 169:30]
  wire  _GEN_7727 = uncached ? _GEN_2311 : _GEN_6176; // @[ICache.scala 169:30]
  wire  _GEN_7728 = uncached ? _GEN_2823 : _GEN_6177; // @[ICache.scala 169:30]
  wire  _GEN_7729 = uncached ? _GEN_2312 : _GEN_6178; // @[ICache.scala 169:30]
  wire  _GEN_7730 = uncached ? _GEN_2824 : _GEN_6179; // @[ICache.scala 169:30]
  wire  _GEN_7731 = uncached ? _GEN_2313 : _GEN_6180; // @[ICache.scala 169:30]
  wire  _GEN_7732 = uncached ? _GEN_2825 : _GEN_6181; // @[ICache.scala 169:30]
  wire  _GEN_7733 = uncached ? _GEN_2314 : _GEN_6182; // @[ICache.scala 169:30]
  wire  _GEN_7734 = uncached ? _GEN_2826 : _GEN_6183; // @[ICache.scala 169:30]
  wire  _GEN_7735 = uncached ? _GEN_2315 : _GEN_6184; // @[ICache.scala 169:30]
  wire  _GEN_7736 = uncached ? _GEN_2827 : _GEN_6185; // @[ICache.scala 169:30]
  wire  _GEN_7737 = uncached ? _GEN_2316 : _GEN_6186; // @[ICache.scala 169:30]
  wire  _GEN_7738 = uncached ? _GEN_2828 : _GEN_6187; // @[ICache.scala 169:30]
  wire  _GEN_7739 = uncached ? _GEN_2317 : _GEN_6188; // @[ICache.scala 169:30]
  wire  _GEN_7740 = uncached ? _GEN_2829 : _GEN_6189; // @[ICache.scala 169:30]
  wire  _GEN_7741 = uncached ? _GEN_2318 : _GEN_6190; // @[ICache.scala 169:30]
  wire  _GEN_7742 = uncached ? _GEN_2830 : _GEN_6191; // @[ICache.scala 169:30]
  wire  _GEN_7743 = uncached ? _GEN_2319 : _GEN_6192; // @[ICache.scala 169:30]
  wire  _GEN_7744 = uncached ? _GEN_2831 : _GEN_6193; // @[ICache.scala 169:30]
  wire  _GEN_7745 = uncached ? _GEN_2320 : _GEN_6194; // @[ICache.scala 169:30]
  wire  _GEN_7746 = uncached ? _GEN_2832 : _GEN_6195; // @[ICache.scala 169:30]
  wire  _GEN_7747 = uncached ? _GEN_2321 : _GEN_6196; // @[ICache.scala 169:30]
  wire  _GEN_7748 = uncached ? _GEN_2833 : _GEN_6197; // @[ICache.scala 169:30]
  wire  _GEN_7749 = uncached ? _GEN_2322 : _GEN_6198; // @[ICache.scala 169:30]
  wire  _GEN_7750 = uncached ? _GEN_2834 : _GEN_6199; // @[ICache.scala 169:30]
  wire  _GEN_7751 = uncached ? _GEN_2323 : _GEN_6200; // @[ICache.scala 169:30]
  wire  _GEN_7752 = uncached ? _GEN_2835 : _GEN_6201; // @[ICache.scala 169:30]
  wire  _GEN_7753 = uncached ? _GEN_2324 : _GEN_6202; // @[ICache.scala 169:30]
  wire  _GEN_7754 = uncached ? _GEN_2836 : _GEN_6203; // @[ICache.scala 169:30]
  wire  _GEN_7755 = uncached ? _GEN_2325 : _GEN_6204; // @[ICache.scala 169:30]
  wire  _GEN_7756 = uncached ? _GEN_2837 : _GEN_6205; // @[ICache.scala 169:30]
  wire  _GEN_7757 = uncached ? _GEN_2326 : _GEN_6206; // @[ICache.scala 169:30]
  wire  _GEN_7758 = uncached ? _GEN_2838 : _GEN_6207; // @[ICache.scala 169:30]
  wire  _GEN_7759 = uncached ? _GEN_2327 : _GEN_6208; // @[ICache.scala 169:30]
  wire  _GEN_7760 = uncached ? _GEN_2839 : _GEN_6209; // @[ICache.scala 169:30]
  wire  _GEN_7761 = uncached ? _GEN_2328 : _GEN_6210; // @[ICache.scala 169:30]
  wire  _GEN_7762 = uncached ? _GEN_2840 : _GEN_6211; // @[ICache.scala 169:30]
  wire  _GEN_7763 = uncached ? _GEN_2329 : _GEN_6212; // @[ICache.scala 169:30]
  wire  _GEN_7764 = uncached ? _GEN_2841 : _GEN_6213; // @[ICache.scala 169:30]
  wire  _GEN_7765 = uncached ? _GEN_2330 : _GEN_6214; // @[ICache.scala 169:30]
  wire  _GEN_7766 = uncached ? _GEN_2842 : _GEN_6215; // @[ICache.scala 169:30]
  wire  _GEN_7767 = uncached ? _GEN_2331 : _GEN_6216; // @[ICache.scala 169:30]
  wire  _GEN_7768 = uncached ? _GEN_2843 : _GEN_6217; // @[ICache.scala 169:30]
  wire  _GEN_7769 = uncached ? _GEN_2332 : _GEN_6218; // @[ICache.scala 169:30]
  wire  _GEN_7770 = uncached ? _GEN_2844 : _GEN_6219; // @[ICache.scala 169:30]
  wire  _GEN_7771 = uncached ? _GEN_2333 : _GEN_6220; // @[ICache.scala 169:30]
  wire  _GEN_7772 = uncached ? _GEN_2845 : _GEN_6221; // @[ICache.scala 169:30]
  wire  _GEN_7773 = uncached ? _GEN_2334 : _GEN_6222; // @[ICache.scala 169:30]
  wire  _GEN_7774 = uncached ? _GEN_2846 : _GEN_6223; // @[ICache.scala 169:30]
  wire  _GEN_7775 = uncached ? _GEN_2335 : _GEN_6224; // @[ICache.scala 169:30]
  wire  _GEN_7776 = uncached ? _GEN_2847 : _GEN_6225; // @[ICache.scala 169:30]
  wire  _GEN_7777 = uncached ? _GEN_2336 : _GEN_6226; // @[ICache.scala 169:30]
  wire  _GEN_7778 = uncached ? _GEN_2848 : _GEN_6227; // @[ICache.scala 169:30]
  wire  _GEN_7779 = uncached ? _GEN_2337 : _GEN_6228; // @[ICache.scala 169:30]
  wire  _GEN_7780 = uncached ? _GEN_2849 : _GEN_6229; // @[ICache.scala 169:30]
  wire  _GEN_7781 = uncached ? _GEN_2338 : _GEN_6230; // @[ICache.scala 169:30]
  wire  _GEN_7782 = uncached ? _GEN_2850 : _GEN_6231; // @[ICache.scala 169:30]
  wire  _GEN_7783 = uncached ? _GEN_2339 : _GEN_6232; // @[ICache.scala 169:30]
  wire  _GEN_7784 = uncached ? _GEN_2851 : _GEN_6233; // @[ICache.scala 169:30]
  wire  _GEN_7785 = uncached ? _GEN_2340 : _GEN_6234; // @[ICache.scala 169:30]
  wire  _GEN_7786 = uncached ? _GEN_2852 : _GEN_6235; // @[ICache.scala 169:30]
  wire  _GEN_7787 = uncached ? _GEN_2341 : _GEN_6236; // @[ICache.scala 169:30]
  wire  _GEN_7788 = uncached ? _GEN_2853 : _GEN_6237; // @[ICache.scala 169:30]
  wire  _GEN_7789 = uncached ? _GEN_2342 : _GEN_6238; // @[ICache.scala 169:30]
  wire  _GEN_7790 = uncached ? _GEN_2854 : _GEN_6239; // @[ICache.scala 169:30]
  wire  _GEN_7791 = uncached ? _GEN_2343 : _GEN_6240; // @[ICache.scala 169:30]
  wire  _GEN_7792 = uncached ? _GEN_2855 : _GEN_6241; // @[ICache.scala 169:30]
  wire  _GEN_7793 = uncached ? _GEN_2344 : _GEN_6242; // @[ICache.scala 169:30]
  wire  _GEN_7794 = uncached ? _GEN_2856 : _GEN_6243; // @[ICache.scala 169:30]
  wire  _GEN_7795 = uncached ? _GEN_2345 : _GEN_6244; // @[ICache.scala 169:30]
  wire  _GEN_7796 = uncached ? _GEN_2857 : _GEN_6245; // @[ICache.scala 169:30]
  wire  _GEN_7797 = uncached ? _GEN_2346 : _GEN_6246; // @[ICache.scala 169:30]
  wire  _GEN_7798 = uncached ? _GEN_2858 : _GEN_6247; // @[ICache.scala 169:30]
  wire  _GEN_7799 = uncached ? _GEN_2347 : _GEN_6248; // @[ICache.scala 169:30]
  wire  _GEN_7800 = uncached ? _GEN_2859 : _GEN_6249; // @[ICache.scala 169:30]
  wire  _GEN_7801 = uncached ? _GEN_2348 : _GEN_6250; // @[ICache.scala 169:30]
  wire  _GEN_7802 = uncached ? _GEN_2860 : _GEN_6251; // @[ICache.scala 169:30]
  wire  _GEN_7803 = uncached ? _GEN_2349 : _GEN_6252; // @[ICache.scala 169:30]
  wire  _GEN_7804 = uncached ? _GEN_2861 : _GEN_6253; // @[ICache.scala 169:30]
  wire  _GEN_7805 = uncached ? _GEN_2350 : _GEN_6254; // @[ICache.scala 169:30]
  wire  _GEN_7806 = uncached ? _GEN_2862 : _GEN_6255; // @[ICache.scala 169:30]
  wire  _GEN_7807 = uncached ? _GEN_2351 : _GEN_6256; // @[ICache.scala 169:30]
  wire  _GEN_7808 = uncached ? _GEN_2863 : _GEN_6257; // @[ICache.scala 169:30]
  wire  _GEN_7809 = uncached ? _GEN_2352 : _GEN_6258; // @[ICache.scala 169:30]
  wire  _GEN_7810 = uncached ? _GEN_2864 : _GEN_6259; // @[ICache.scala 169:30]
  wire  _GEN_7811 = uncached ? _GEN_2353 : _GEN_6260; // @[ICache.scala 169:30]
  wire  _GEN_7812 = uncached ? _GEN_2865 : _GEN_6261; // @[ICache.scala 169:30]
  wire  _GEN_7813 = uncached ? _GEN_2354 : _GEN_6262; // @[ICache.scala 169:30]
  wire  _GEN_7814 = uncached ? _GEN_2866 : _GEN_6263; // @[ICache.scala 169:30]
  wire  _GEN_7815 = uncached ? _GEN_2355 : _GEN_6264; // @[ICache.scala 169:30]
  wire  _GEN_7816 = uncached ? _GEN_2867 : _GEN_6265; // @[ICache.scala 169:30]
  wire  _GEN_7817 = uncached ? _GEN_2356 : _GEN_6266; // @[ICache.scala 169:30]
  wire  _GEN_7818 = uncached ? _GEN_2868 : _GEN_6267; // @[ICache.scala 169:30]
  wire  _GEN_7819 = uncached ? _GEN_2357 : _GEN_6268; // @[ICache.scala 169:30]
  wire  _GEN_7820 = uncached ? _GEN_2869 : _GEN_6269; // @[ICache.scala 169:30]
  wire  _GEN_7821 = uncached ? _GEN_2358 : _GEN_6270; // @[ICache.scala 169:30]
  wire  _GEN_7822 = uncached ? _GEN_2870 : _GEN_6271; // @[ICache.scala 169:30]
  wire  _GEN_7823 = uncached ? _GEN_2359 : _GEN_6272; // @[ICache.scala 169:30]
  wire  _GEN_7824 = uncached ? _GEN_2871 : _GEN_6273; // @[ICache.scala 169:30]
  wire  _GEN_7825 = uncached ? _GEN_2360 : _GEN_6274; // @[ICache.scala 169:30]
  wire  _GEN_7826 = uncached ? _GEN_2872 : _GEN_6275; // @[ICache.scala 169:30]
  wire  _GEN_7827 = uncached ? _GEN_2361 : _GEN_6276; // @[ICache.scala 169:30]
  wire  _GEN_7828 = uncached ? _GEN_2873 : _GEN_6277; // @[ICache.scala 169:30]
  wire  _GEN_7829 = uncached ? _GEN_2362 : _GEN_6278; // @[ICache.scala 169:30]
  wire  _GEN_7830 = uncached ? _GEN_2874 : _GEN_6279; // @[ICache.scala 169:30]
  wire  _GEN_7831 = uncached ? _GEN_2363 : _GEN_6280; // @[ICache.scala 169:30]
  wire  _GEN_7832 = uncached ? _GEN_2875 : _GEN_6281; // @[ICache.scala 169:30]
  wire  _GEN_7833 = uncached ? _GEN_2364 : _GEN_6282; // @[ICache.scala 169:30]
  wire  _GEN_7834 = uncached ? _GEN_2876 : _GEN_6283; // @[ICache.scala 169:30]
  wire  _GEN_7835 = uncached ? _GEN_2365 : _GEN_6284; // @[ICache.scala 169:30]
  wire  _GEN_7836 = uncached ? _GEN_2877 : _GEN_6285; // @[ICache.scala 169:30]
  wire  _GEN_7837 = uncached ? _GEN_2366 : _GEN_6286; // @[ICache.scala 169:30]
  wire  _GEN_7838 = uncached ? _GEN_2878 : _GEN_6287; // @[ICache.scala 169:30]
  wire  _GEN_7839 = uncached ? _GEN_2367 : _GEN_6288; // @[ICache.scala 169:30]
  wire  _GEN_7840 = uncached ? _GEN_2879 : _GEN_6289; // @[ICache.scala 169:30]
  wire  _GEN_7841 = uncached ? _GEN_2368 : _GEN_6290; // @[ICache.scala 169:30]
  wire  _GEN_7842 = uncached ? _GEN_2880 : _GEN_6291; // @[ICache.scala 169:30]
  wire  _GEN_7843 = uncached ? _GEN_2369 : _GEN_6292; // @[ICache.scala 169:30]
  wire  _GEN_7844 = uncached ? _GEN_2881 : _GEN_6293; // @[ICache.scala 169:30]
  wire  _GEN_7845 = uncached ? _GEN_2370 : _GEN_6294; // @[ICache.scala 169:30]
  wire  _GEN_7846 = uncached ? _GEN_2882 : _GEN_6295; // @[ICache.scala 169:30]
  wire  _GEN_7847 = uncached ? _GEN_2371 : _GEN_6296; // @[ICache.scala 169:30]
  wire  _GEN_7848 = uncached ? _GEN_2883 : _GEN_6297; // @[ICache.scala 169:30]
  wire  _GEN_7849 = uncached ? _GEN_2372 : _GEN_6298; // @[ICache.scala 169:30]
  wire  _GEN_7850 = uncached ? _GEN_2884 : _GEN_6299; // @[ICache.scala 169:30]
  wire  _GEN_7851 = uncached ? _GEN_2373 : _GEN_6300; // @[ICache.scala 169:30]
  wire  _GEN_7852 = uncached ? _GEN_2885 : _GEN_6301; // @[ICache.scala 169:30]
  wire  _GEN_7853 = uncached ? _GEN_2374 : _GEN_6302; // @[ICache.scala 169:30]
  wire  _GEN_7854 = uncached ? _GEN_2886 : _GEN_6303; // @[ICache.scala 169:30]
  wire  _GEN_7855 = uncached ? _GEN_2375 : _GEN_6304; // @[ICache.scala 169:30]
  wire  _GEN_7856 = uncached ? _GEN_2887 : _GEN_6305; // @[ICache.scala 169:30]
  wire  _GEN_7857 = uncached ? _GEN_2376 : _GEN_6306; // @[ICache.scala 169:30]
  wire  _GEN_7858 = uncached ? _GEN_2888 : _GEN_6307; // @[ICache.scala 169:30]
  wire  _GEN_7859 = uncached ? _GEN_2377 : _GEN_6308; // @[ICache.scala 169:30]
  wire  _GEN_7860 = uncached ? _GEN_2889 : _GEN_6309; // @[ICache.scala 169:30]
  wire  _GEN_7861 = uncached ? _GEN_2378 : _GEN_6310; // @[ICache.scala 169:30]
  wire  _GEN_7862 = uncached ? _GEN_2890 : _GEN_6311; // @[ICache.scala 169:30]
  wire  _GEN_7863 = uncached ? _GEN_2379 : _GEN_6312; // @[ICache.scala 169:30]
  wire  _GEN_7864 = uncached ? _GEN_2891 : _GEN_6313; // @[ICache.scala 169:30]
  wire  _GEN_7865 = uncached ? _GEN_2380 : _GEN_6314; // @[ICache.scala 169:30]
  wire  _GEN_7866 = uncached ? _GEN_2892 : _GEN_6315; // @[ICache.scala 169:30]
  wire  _GEN_7867 = uncached ? _GEN_2381 : _GEN_6316; // @[ICache.scala 169:30]
  wire  _GEN_7868 = uncached ? _GEN_2893 : _GEN_6317; // @[ICache.scala 169:30]
  wire  _GEN_7869 = uncached ? _GEN_2382 : _GEN_6318; // @[ICache.scala 169:30]
  wire  _GEN_7870 = uncached ? _GEN_2894 : _GEN_6319; // @[ICache.scala 169:30]
  wire  _GEN_7871 = uncached ? _GEN_2383 : _GEN_6320; // @[ICache.scala 169:30]
  wire  _GEN_7872 = uncached ? _GEN_2895 : _GEN_6321; // @[ICache.scala 169:30]
  wire  _GEN_7873 = uncached ? _GEN_2384 : _GEN_6322; // @[ICache.scala 169:30]
  wire  _GEN_7874 = uncached ? _GEN_2896 : _GEN_6323; // @[ICache.scala 169:30]
  wire  _GEN_7875 = uncached ? _GEN_2385 : _GEN_6324; // @[ICache.scala 169:30]
  wire  _GEN_7876 = uncached ? _GEN_2897 : _GEN_6325; // @[ICache.scala 169:30]
  wire  _GEN_7877 = uncached ? _GEN_2386 : _GEN_6326; // @[ICache.scala 169:30]
  wire  _GEN_7878 = uncached ? _GEN_2898 : _GEN_6327; // @[ICache.scala 169:30]
  wire  _GEN_7879 = uncached ? _GEN_2387 : _GEN_6328; // @[ICache.scala 169:30]
  wire  _GEN_7880 = uncached ? _GEN_2899 : _GEN_6329; // @[ICache.scala 169:30]
  wire  _GEN_7881 = uncached ? _GEN_2388 : _GEN_6330; // @[ICache.scala 169:30]
  wire  _GEN_7882 = uncached ? _GEN_2900 : _GEN_6331; // @[ICache.scala 169:30]
  wire  _GEN_7883 = uncached ? _GEN_2389 : _GEN_6332; // @[ICache.scala 169:30]
  wire  _GEN_7884 = uncached ? _GEN_2901 : _GEN_6333; // @[ICache.scala 169:30]
  wire  _GEN_7885 = uncached ? _GEN_2390 : _GEN_6334; // @[ICache.scala 169:30]
  wire  _GEN_7886 = uncached ? _GEN_2902 : _GEN_6335; // @[ICache.scala 169:30]
  wire  _GEN_7887 = uncached ? _GEN_2391 : _GEN_6336; // @[ICache.scala 169:30]
  wire  _GEN_7888 = uncached ? _GEN_2903 : _GEN_6337; // @[ICache.scala 169:30]
  wire  _GEN_7889 = uncached ? _GEN_2392 : _GEN_6338; // @[ICache.scala 169:30]
  wire  _GEN_7890 = uncached ? _GEN_2904 : _GEN_6339; // @[ICache.scala 169:30]
  wire  _GEN_7891 = uncached ? _GEN_2393 : _GEN_6340; // @[ICache.scala 169:30]
  wire  _GEN_7892 = uncached ? _GEN_2905 : _GEN_6341; // @[ICache.scala 169:30]
  wire  _GEN_7893 = uncached ? _GEN_2394 : _GEN_6342; // @[ICache.scala 169:30]
  wire  _GEN_7894 = uncached ? _GEN_2906 : _GEN_6343; // @[ICache.scala 169:30]
  wire  _GEN_7895 = uncached ? _GEN_2395 : _GEN_6344; // @[ICache.scala 169:30]
  wire  _GEN_7896 = uncached ? _GEN_2907 : _GEN_6345; // @[ICache.scala 169:30]
  wire  _GEN_7897 = uncached ? _GEN_2396 : _GEN_6346; // @[ICache.scala 169:30]
  wire  _GEN_7898 = uncached ? _GEN_2908 : _GEN_6347; // @[ICache.scala 169:30]
  wire  _GEN_7899 = uncached ? _GEN_2397 : _GEN_6348; // @[ICache.scala 169:30]
  wire  _GEN_7900 = uncached ? _GEN_2909 : _GEN_6349; // @[ICache.scala 169:30]
  wire  _GEN_7901 = uncached ? _GEN_2398 : _GEN_6350; // @[ICache.scala 169:30]
  wire  _GEN_7902 = uncached ? _GEN_2910 : _GEN_6351; // @[ICache.scala 169:30]
  wire  _GEN_7903 = uncached ? _GEN_2399 : _GEN_6352; // @[ICache.scala 169:30]
  wire  _GEN_7904 = uncached ? _GEN_2911 : _GEN_6353; // @[ICache.scala 169:30]
  wire  _GEN_7905 = uncached ? _GEN_2400 : _GEN_6354; // @[ICache.scala 169:30]
  wire  _GEN_7906 = uncached ? _GEN_2912 : _GEN_6355; // @[ICache.scala 169:30]
  wire  _GEN_7907 = uncached ? _GEN_2401 : _GEN_6356; // @[ICache.scala 169:30]
  wire  _GEN_7908 = uncached ? _GEN_2913 : _GEN_6357; // @[ICache.scala 169:30]
  wire  _GEN_7909 = uncached ? _GEN_2402 : _GEN_6358; // @[ICache.scala 169:30]
  wire  _GEN_7910 = uncached ? _GEN_2914 : _GEN_6359; // @[ICache.scala 169:30]
  wire  _GEN_7911 = uncached ? _GEN_2403 : _GEN_6360; // @[ICache.scala 169:30]
  wire  _GEN_7912 = uncached ? _GEN_2915 : _GEN_6361; // @[ICache.scala 169:30]
  wire  _GEN_7913 = uncached ? _GEN_2404 : _GEN_6362; // @[ICache.scala 169:30]
  wire  _GEN_7914 = uncached ? _GEN_2916 : _GEN_6363; // @[ICache.scala 169:30]
  wire  _GEN_7915 = uncached ? _GEN_2405 : _GEN_6364; // @[ICache.scala 169:30]
  wire  _GEN_7916 = uncached ? _GEN_2917 : _GEN_6365; // @[ICache.scala 169:30]
  wire  _GEN_7917 = uncached ? _GEN_2406 : _GEN_6366; // @[ICache.scala 169:30]
  wire  _GEN_7918 = uncached ? _GEN_2918 : _GEN_6367; // @[ICache.scala 169:30]
  wire  _GEN_7919 = uncached ? _GEN_2407 : _GEN_6368; // @[ICache.scala 169:30]
  wire  _GEN_7920 = uncached ? _GEN_2919 : _GEN_6369; // @[ICache.scala 169:30]
  wire  _GEN_7921 = uncached ? _GEN_2408 : _GEN_6370; // @[ICache.scala 169:30]
  wire  _GEN_7922 = uncached ? _GEN_2920 : _GEN_6371; // @[ICache.scala 169:30]
  wire  _GEN_7923 = uncached ? _GEN_2409 : _GEN_6372; // @[ICache.scala 169:30]
  wire  _GEN_7924 = uncached ? _GEN_2921 : _GEN_6373; // @[ICache.scala 169:30]
  wire  _GEN_7925 = uncached ? _GEN_2410 : _GEN_6374; // @[ICache.scala 169:30]
  wire  _GEN_7926 = uncached ? _GEN_2922 : _GEN_6375; // @[ICache.scala 169:30]
  wire  _GEN_7927 = uncached ? _GEN_2411 : _GEN_6376; // @[ICache.scala 169:30]
  wire  _GEN_7928 = uncached ? _GEN_2923 : _GEN_6377; // @[ICache.scala 169:30]
  wire  _GEN_7929 = uncached ? _GEN_2412 : _GEN_6378; // @[ICache.scala 169:30]
  wire  _GEN_7930 = uncached ? _GEN_2924 : _GEN_6379; // @[ICache.scala 169:30]
  wire  _GEN_7931 = uncached ? _GEN_2413 : _GEN_6380; // @[ICache.scala 169:30]
  wire  _GEN_7932 = uncached ? _GEN_2925 : _GEN_6381; // @[ICache.scala 169:30]
  wire  _GEN_7933 = uncached ? _GEN_2414 : _GEN_6382; // @[ICache.scala 169:30]
  wire  _GEN_7934 = uncached ? _GEN_2926 : _GEN_6383; // @[ICache.scala 169:30]
  wire  _GEN_7935 = uncached ? _GEN_2415 : _GEN_6384; // @[ICache.scala 169:30]
  wire  _GEN_7936 = uncached ? _GEN_2927 : _GEN_6385; // @[ICache.scala 169:30]
  wire  _GEN_7937 = uncached ? _GEN_2416 : _GEN_6386; // @[ICache.scala 169:30]
  wire  _GEN_7938 = uncached ? _GEN_2928 : _GEN_6387; // @[ICache.scala 169:30]
  wire  _GEN_7939 = uncached ? _GEN_2417 : _GEN_6388; // @[ICache.scala 169:30]
  wire  _GEN_7940 = uncached ? _GEN_2929 : _GEN_6389; // @[ICache.scala 169:30]
  wire  _GEN_7941 = uncached ? _GEN_2418 : _GEN_6390; // @[ICache.scala 169:30]
  wire  _GEN_7942 = uncached ? _GEN_2930 : _GEN_6391; // @[ICache.scala 169:30]
  wire  _GEN_7943 = uncached ? _GEN_2419 : _GEN_6392; // @[ICache.scala 169:30]
  wire  _GEN_7944 = uncached ? _GEN_2931 : _GEN_6393; // @[ICache.scala 169:30]
  wire  _GEN_7945 = uncached ? _GEN_2420 : _GEN_6394; // @[ICache.scala 169:30]
  wire  _GEN_7946 = uncached ? _GEN_2932 : _GEN_6395; // @[ICache.scala 169:30]
  wire  _GEN_7947 = uncached ? _GEN_2421 : _GEN_6396; // @[ICache.scala 169:30]
  wire  _GEN_7948 = uncached ? _GEN_2933 : _GEN_6397; // @[ICache.scala 169:30]
  wire  _GEN_7949 = uncached ? _GEN_2422 : _GEN_6398; // @[ICache.scala 169:30]
  wire  _GEN_7950 = uncached ? _GEN_2934 : _GEN_6399; // @[ICache.scala 169:30]
  wire  _GEN_7951 = uncached ? _GEN_2423 : _GEN_6400; // @[ICache.scala 169:30]
  wire  _GEN_7952 = uncached ? _GEN_2935 : _GEN_6401; // @[ICache.scala 169:30]
  wire  _GEN_7953 = uncached ? _GEN_2424 : _GEN_6402; // @[ICache.scala 169:30]
  wire  _GEN_7954 = uncached ? _GEN_2936 : _GEN_6403; // @[ICache.scala 169:30]
  wire  _GEN_7955 = uncached ? _GEN_2425 : _GEN_6404; // @[ICache.scala 169:30]
  wire  _GEN_7956 = uncached ? _GEN_2937 : _GEN_6405; // @[ICache.scala 169:30]
  wire  _GEN_7957 = uncached ? _GEN_2426 : _GEN_6406; // @[ICache.scala 169:30]
  wire  _GEN_7958 = uncached ? _GEN_2938 : _GEN_6407; // @[ICache.scala 169:30]
  wire  _GEN_7959 = uncached ? _GEN_2427 : _GEN_6408; // @[ICache.scala 169:30]
  wire  _GEN_7960 = uncached ? _GEN_2939 : _GEN_6409; // @[ICache.scala 169:30]
  wire  _GEN_7961 = uncached ? _GEN_2428 : _GEN_6410; // @[ICache.scala 169:30]
  wire  _GEN_7962 = uncached ? _GEN_2940 : _GEN_6411; // @[ICache.scala 169:30]
  wire  _GEN_7963 = uncached ? _GEN_2429 : _GEN_6412; // @[ICache.scala 169:30]
  wire  _GEN_7964 = uncached ? _GEN_2941 : _GEN_6413; // @[ICache.scala 169:30]
  wire  _GEN_7965 = uncached ? _GEN_2430 : _GEN_6414; // @[ICache.scala 169:30]
  wire  _GEN_7966 = uncached ? _GEN_2942 : _GEN_6415; // @[ICache.scala 169:30]
  wire  _GEN_7967 = uncached ? _GEN_2431 : _GEN_6416; // @[ICache.scala 169:30]
  wire  _GEN_7968 = uncached ? _GEN_2943 : _GEN_6417; // @[ICache.scala 169:30]
  wire  _GEN_7969 = uncached ? _GEN_2432 : _GEN_6418; // @[ICache.scala 169:30]
  wire  _GEN_7970 = uncached ? _GEN_2944 : _GEN_6419; // @[ICache.scala 169:30]
  wire  _GEN_7971 = uncached ? _GEN_2433 : _GEN_6420; // @[ICache.scala 169:30]
  wire  _GEN_7972 = uncached ? _GEN_2945 : _GEN_6421; // @[ICache.scala 169:30]
  wire  _GEN_7973 = uncached ? _GEN_2434 : _GEN_6422; // @[ICache.scala 169:30]
  wire  _GEN_7974 = uncached ? _GEN_2946 : _GEN_6423; // @[ICache.scala 169:30]
  wire  _GEN_7975 = uncached ? _GEN_2435 : _GEN_6424; // @[ICache.scala 169:30]
  wire  _GEN_7976 = uncached ? _GEN_2947 : _GEN_6425; // @[ICache.scala 169:30]
  wire  _GEN_7977 = uncached ? _GEN_2436 : _GEN_6426; // @[ICache.scala 169:30]
  wire  _GEN_7978 = uncached ? _GEN_2948 : _GEN_6427; // @[ICache.scala 169:30]
  wire  _GEN_7979 = uncached ? _GEN_2437 : _GEN_6428; // @[ICache.scala 169:30]
  wire  _GEN_7980 = uncached ? _GEN_2949 : _GEN_6429; // @[ICache.scala 169:30]
  wire  _GEN_7981 = uncached ? _GEN_2438 : _GEN_6430; // @[ICache.scala 169:30]
  wire  _GEN_7982 = uncached ? _GEN_2950 : _GEN_6431; // @[ICache.scala 169:30]
  wire  _GEN_7983 = uncached ? _GEN_2439 : _GEN_6432; // @[ICache.scala 169:30]
  wire  _GEN_7984 = uncached ? _GEN_2951 : _GEN_6433; // @[ICache.scala 169:30]
  wire  _GEN_7985 = uncached ? _GEN_2440 : _GEN_6434; // @[ICache.scala 169:30]
  wire  _GEN_7986 = uncached ? _GEN_2952 : _GEN_6435; // @[ICache.scala 169:30]
  wire  _GEN_7987 = uncached ? _GEN_2441 : _GEN_6436; // @[ICache.scala 169:30]
  wire  _GEN_7988 = uncached ? _GEN_2953 : _GEN_6437; // @[ICache.scala 169:30]
  wire  _GEN_7989 = uncached ? _GEN_2442 : _GEN_6438; // @[ICache.scala 169:30]
  wire  _GEN_7990 = uncached ? _GEN_2954 : _GEN_6439; // @[ICache.scala 169:30]
  wire  _GEN_7991 = uncached ? _GEN_2443 : _GEN_6440; // @[ICache.scala 169:30]
  wire  _GEN_7992 = uncached ? _GEN_2955 : _GEN_6441; // @[ICache.scala 169:30]
  wire  _GEN_7993 = uncached ? _GEN_2444 : _GEN_6442; // @[ICache.scala 169:30]
  wire  _GEN_7994 = uncached ? _GEN_2956 : _GEN_6443; // @[ICache.scala 169:30]
  wire  _GEN_7995 = uncached ? _GEN_2445 : _GEN_6444; // @[ICache.scala 169:30]
  wire  _GEN_7996 = uncached ? _GEN_2957 : _GEN_6445; // @[ICache.scala 169:30]
  wire  _GEN_7997 = uncached ? _GEN_2446 : _GEN_6446; // @[ICache.scala 169:30]
  wire  _GEN_7998 = uncached ? _GEN_2958 : _GEN_6447; // @[ICache.scala 169:30]
  wire  _GEN_7999 = uncached ? _GEN_2447 : _GEN_6448; // @[ICache.scala 169:30]
  wire  _GEN_8000 = uncached ? _GEN_2959 : _GEN_6449; // @[ICache.scala 169:30]
  wire  _GEN_8001 = uncached ? _GEN_2448 : _GEN_6450; // @[ICache.scala 169:30]
  wire  _GEN_8002 = uncached ? _GEN_2960 : _GEN_6451; // @[ICache.scala 169:30]
  wire  _GEN_8003 = uncached ? _GEN_2449 : _GEN_6452; // @[ICache.scala 169:30]
  wire  _GEN_8004 = uncached ? _GEN_2961 : _GEN_6453; // @[ICache.scala 169:30]
  wire  _GEN_8005 = uncached ? _GEN_2450 : _GEN_6454; // @[ICache.scala 169:30]
  wire  _GEN_8006 = uncached ? _GEN_2962 : _GEN_6455; // @[ICache.scala 169:30]
  wire  _GEN_8007 = uncached ? _GEN_2451 : _GEN_6456; // @[ICache.scala 169:30]
  wire  _GEN_8008 = uncached ? _GEN_2963 : _GEN_6457; // @[ICache.scala 169:30]
  wire  _GEN_8009 = uncached ? _GEN_2452 : _GEN_6458; // @[ICache.scala 169:30]
  wire  _GEN_8010 = uncached ? _GEN_2964 : _GEN_6459; // @[ICache.scala 169:30]
  wire  _GEN_8011 = uncached ? _GEN_2453 : _GEN_6460; // @[ICache.scala 169:30]
  wire  _GEN_8012 = uncached ? _GEN_2965 : _GEN_6461; // @[ICache.scala 169:30]
  wire  _GEN_8013 = uncached ? _GEN_2454 : _GEN_6462; // @[ICache.scala 169:30]
  wire  _GEN_8014 = uncached ? _GEN_2966 : _GEN_6463; // @[ICache.scala 169:30]
  wire  _GEN_8015 = uncached ? _GEN_2455 : _GEN_6464; // @[ICache.scala 169:30]
  wire  _GEN_8016 = uncached ? _GEN_2967 : _GEN_6465; // @[ICache.scala 169:30]
  wire  _GEN_8017 = uncached ? _GEN_2456 : _GEN_6466; // @[ICache.scala 169:30]
  wire  _GEN_8018 = uncached ? _GEN_2968 : _GEN_6467; // @[ICache.scala 169:30]
  wire  _GEN_8019 = uncached ? _GEN_2457 : _GEN_6468; // @[ICache.scala 169:30]
  wire  _GEN_8020 = uncached ? _GEN_2969 : _GEN_6469; // @[ICache.scala 169:30]
  wire  _GEN_8021 = uncached ? _GEN_2458 : _GEN_6470; // @[ICache.scala 169:30]
  wire  _GEN_8022 = uncached ? _GEN_2970 : _GEN_6471; // @[ICache.scala 169:30]
  wire  _GEN_8023 = uncached ? _GEN_2459 : _GEN_6472; // @[ICache.scala 169:30]
  wire  _GEN_8024 = uncached ? _GEN_2971 : _GEN_6473; // @[ICache.scala 169:30]
  wire  _GEN_8025 = uncached ? _GEN_2460 : _GEN_6474; // @[ICache.scala 169:30]
  wire  _GEN_8026 = uncached ? _GEN_2972 : _GEN_6475; // @[ICache.scala 169:30]
  wire  _GEN_8027 = uncached ? _GEN_2461 : _GEN_6476; // @[ICache.scala 169:30]
  wire  _GEN_8028 = uncached ? _GEN_2973 : _GEN_6477; // @[ICache.scala 169:30]
  wire  _GEN_8029 = uncached ? _GEN_2462 : _GEN_6478; // @[ICache.scala 169:30]
  wire  _GEN_8030 = uncached ? _GEN_2974 : _GEN_6479; // @[ICache.scala 169:30]
  wire  _GEN_8031 = uncached ? _GEN_2463 : _GEN_6480; // @[ICache.scala 169:30]
  wire  _GEN_8032 = uncached ? _GEN_2975 : _GEN_6481; // @[ICache.scala 169:30]
  wire  _GEN_8033 = uncached ? _GEN_2464 : _GEN_6482; // @[ICache.scala 169:30]
  wire  _GEN_8034 = uncached ? _GEN_2976 : _GEN_6483; // @[ICache.scala 169:30]
  wire  _GEN_8035 = uncached ? _GEN_2465 : _GEN_6484; // @[ICache.scala 169:30]
  wire  _GEN_8036 = uncached ? _GEN_2977 : _GEN_6485; // @[ICache.scala 169:30]
  wire  _GEN_8037 = uncached ? _GEN_2466 : _GEN_6486; // @[ICache.scala 169:30]
  wire  _GEN_8038 = uncached ? _GEN_2978 : _GEN_6487; // @[ICache.scala 169:30]
  wire  _GEN_8039 = uncached ? _GEN_2467 : _GEN_6488; // @[ICache.scala 169:30]
  wire  _GEN_8040 = uncached ? _GEN_2979 : _GEN_6489; // @[ICache.scala 169:30]
  wire  _GEN_8041 = uncached ? _GEN_2468 : _GEN_6490; // @[ICache.scala 169:30]
  wire  _GEN_8042 = uncached ? _GEN_2980 : _GEN_6491; // @[ICache.scala 169:30]
  wire  _GEN_8043 = uncached ? _GEN_2469 : _GEN_6492; // @[ICache.scala 169:30]
  wire  _GEN_8044 = uncached ? _GEN_2981 : _GEN_6493; // @[ICache.scala 169:30]
  wire  _GEN_8045 = uncached ? _GEN_2470 : _GEN_6494; // @[ICache.scala 169:30]
  wire  _GEN_8046 = uncached ? _GEN_2982 : _GEN_6495; // @[ICache.scala 169:30]
  wire  _GEN_8047 = uncached ? _GEN_2471 : _GEN_6496; // @[ICache.scala 169:30]
  wire  _GEN_8048 = uncached ? _GEN_2983 : _GEN_6497; // @[ICache.scala 169:30]
  wire  _GEN_8049 = uncached ? _GEN_2472 : _GEN_6498; // @[ICache.scala 169:30]
  wire  _GEN_8050 = uncached ? _GEN_2984 : _GEN_6499; // @[ICache.scala 169:30]
  wire  _GEN_8051 = uncached ? _GEN_2473 : _GEN_6500; // @[ICache.scala 169:30]
  wire  _GEN_8052 = uncached ? _GEN_2985 : _GEN_6501; // @[ICache.scala 169:30]
  wire  _GEN_8053 = uncached ? _GEN_2474 : _GEN_6502; // @[ICache.scala 169:30]
  wire  _GEN_8054 = uncached ? _GEN_2986 : _GEN_6503; // @[ICache.scala 169:30]
  wire  _GEN_8055 = uncached ? _GEN_2475 : _GEN_6504; // @[ICache.scala 169:30]
  wire  _GEN_8056 = uncached ? _GEN_2987 : _GEN_6505; // @[ICache.scala 169:30]
  wire  _GEN_8057 = uncached ? _GEN_2476 : _GEN_6506; // @[ICache.scala 169:30]
  wire  _GEN_8058 = uncached ? _GEN_2988 : _GEN_6507; // @[ICache.scala 169:30]
  wire  _GEN_8059 = uncached ? _GEN_2477 : _GEN_6508; // @[ICache.scala 169:30]
  wire  _GEN_8060 = uncached ? _GEN_2989 : _GEN_6509; // @[ICache.scala 169:30]
  wire  _GEN_8061 = uncached ? _GEN_2478 : _GEN_6510; // @[ICache.scala 169:30]
  wire  _GEN_8062 = uncached ? _GEN_2990 : _GEN_6511; // @[ICache.scala 169:30]
  wire  _GEN_8063 = uncached ? _GEN_2479 : _GEN_6512; // @[ICache.scala 169:30]
  wire  _GEN_8064 = uncached ? _GEN_2991 : _GEN_6513; // @[ICache.scala 169:30]
  wire  _GEN_8065 = uncached ? _GEN_2480 : _GEN_6514; // @[ICache.scala 169:30]
  wire  _GEN_8066 = uncached ? _GEN_2992 : _GEN_6515; // @[ICache.scala 169:30]
  wire  _GEN_8067 = uncached ? _GEN_2481 : _GEN_6516; // @[ICache.scala 169:30]
  wire  _GEN_8068 = uncached ? _GEN_2993 : _GEN_6517; // @[ICache.scala 169:30]
  wire  _GEN_8069 = uncached ? _GEN_2482 : _GEN_6518; // @[ICache.scala 169:30]
  wire  _GEN_8070 = uncached ? _GEN_2994 : _GEN_6519; // @[ICache.scala 169:30]
  wire  _GEN_8071 = uncached ? _GEN_2483 : _GEN_6520; // @[ICache.scala 169:30]
  wire  _GEN_8072 = uncached ? _GEN_2995 : _GEN_6521; // @[ICache.scala 169:30]
  wire  _GEN_8073 = uncached ? _GEN_2484 : _GEN_6522; // @[ICache.scala 169:30]
  wire  _GEN_8074 = uncached ? _GEN_2996 : _GEN_6523; // @[ICache.scala 169:30]
  wire  _GEN_8075 = uncached ? _GEN_2485 : _GEN_6524; // @[ICache.scala 169:30]
  wire  _GEN_8076 = uncached ? _GEN_2997 : _GEN_6525; // @[ICache.scala 169:30]
  wire  _GEN_8077 = uncached ? _GEN_2486 : _GEN_6526; // @[ICache.scala 169:30]
  wire  _GEN_8078 = uncached ? _GEN_2998 : _GEN_6527; // @[ICache.scala 169:30]
  wire  _GEN_8079 = uncached ? _GEN_2487 : _GEN_6528; // @[ICache.scala 169:30]
  wire  _GEN_8080 = uncached ? _GEN_2999 : _GEN_6529; // @[ICache.scala 169:30]
  wire  _GEN_8081 = uncached ? _GEN_2488 : _GEN_6530; // @[ICache.scala 169:30]
  wire  _GEN_8082 = uncached ? _GEN_3000 : _GEN_6531; // @[ICache.scala 169:30]
  wire  _GEN_8083 = uncached ? _GEN_2489 : _GEN_6532; // @[ICache.scala 169:30]
  wire  _GEN_8084 = uncached ? _GEN_3001 : _GEN_6533; // @[ICache.scala 169:30]
  wire  _GEN_8085 = uncached ? _GEN_2490 : _GEN_6534; // @[ICache.scala 169:30]
  wire  _GEN_8086 = uncached ? _GEN_3002 : _GEN_6535; // @[ICache.scala 169:30]
  wire  _GEN_8087 = uncached ? _GEN_2491 : _GEN_6536; // @[ICache.scala 169:30]
  wire  _GEN_8088 = uncached ? _GEN_3003 : _GEN_6537; // @[ICache.scala 169:30]
  wire  _GEN_8089 = uncached ? _GEN_2492 : _GEN_6538; // @[ICache.scala 169:30]
  wire  _GEN_8090 = uncached ? _GEN_3004 : _GEN_6539; // @[ICache.scala 169:30]
  wire  _GEN_8091 = uncached ? _GEN_2493 : _GEN_6540; // @[ICache.scala 169:30]
  wire  _GEN_8092 = uncached ? _GEN_3005 : _GEN_6541; // @[ICache.scala 169:30]
  wire  _GEN_8093 = uncached ? _GEN_2494 : _GEN_6542; // @[ICache.scala 169:30]
  wire  _GEN_8094 = uncached ? _GEN_3006 : _GEN_6543; // @[ICache.scala 169:30]
  wire  _GEN_8095 = uncached ? _GEN_2495 : _GEN_6544; // @[ICache.scala 169:30]
  wire  _GEN_8096 = uncached ? _GEN_3007 : _GEN_6545; // @[ICache.scala 169:30]
  wire  _GEN_8097 = uncached ? _GEN_2496 : _GEN_6546; // @[ICache.scala 169:30]
  wire  _GEN_8098 = uncached ? _GEN_3008 : _GEN_6547; // @[ICache.scala 169:30]
  wire  _GEN_8099 = uncached ? _GEN_2497 : _GEN_6548; // @[ICache.scala 169:30]
  wire  _GEN_8100 = uncached ? _GEN_3009 : _GEN_6549; // @[ICache.scala 169:30]
  wire  _GEN_8101 = uncached ? _GEN_2498 : _GEN_6550; // @[ICache.scala 169:30]
  wire  _GEN_8102 = uncached ? _GEN_3010 : _GEN_6551; // @[ICache.scala 169:30]
  wire  _GEN_8103 = uncached ? _GEN_2499 : _GEN_6552; // @[ICache.scala 169:30]
  wire  _GEN_8104 = uncached ? _GEN_3011 : _GEN_6553; // @[ICache.scala 169:30]
  wire  _GEN_8105 = uncached ? _GEN_2500 : _GEN_6554; // @[ICache.scala 169:30]
  wire  _GEN_8106 = uncached ? _GEN_3012 : _GEN_6555; // @[ICache.scala 169:30]
  wire  _GEN_8107 = uncached ? _GEN_2501 : _GEN_6556; // @[ICache.scala 169:30]
  wire  _GEN_8108 = uncached ? _GEN_3013 : _GEN_6557; // @[ICache.scala 169:30]
  wire  _GEN_8109 = uncached ? _GEN_2502 : _GEN_6558; // @[ICache.scala 169:30]
  wire  _GEN_8110 = uncached ? _GEN_3014 : _GEN_6559; // @[ICache.scala 169:30]
  wire  _GEN_8111 = uncached ? _GEN_2503 : _GEN_6560; // @[ICache.scala 169:30]
  wire  _GEN_8112 = uncached ? _GEN_3015 : _GEN_6561; // @[ICache.scala 169:30]
  wire  _GEN_8113 = uncached ? _GEN_2504 : _GEN_6562; // @[ICache.scala 169:30]
  wire  _GEN_8114 = uncached ? _GEN_3016 : _GEN_6563; // @[ICache.scala 169:30]
  wire  _GEN_8115 = uncached ? _GEN_2505 : _GEN_6564; // @[ICache.scala 169:30]
  wire  _GEN_8116 = uncached ? _GEN_3017 : _GEN_6565; // @[ICache.scala 169:30]
  wire  _GEN_8117 = uncached ? _GEN_2506 : _GEN_6566; // @[ICache.scala 169:30]
  wire  _GEN_8118 = uncached ? _GEN_3018 : _GEN_6567; // @[ICache.scala 169:30]
  wire  _GEN_8119 = uncached ? _GEN_2507 : _GEN_6568; // @[ICache.scala 169:30]
  wire  _GEN_8120 = uncached ? _GEN_3019 : _GEN_6569; // @[ICache.scala 169:30]
  wire  _GEN_8121 = uncached ? _GEN_2508 : _GEN_6570; // @[ICache.scala 169:30]
  wire  _GEN_8122 = uncached ? _GEN_3020 : _GEN_6571; // @[ICache.scala 169:30]
  wire  _GEN_8123 = uncached ? _GEN_2509 : _GEN_6572; // @[ICache.scala 169:30]
  wire  _GEN_8124 = uncached ? _GEN_3021 : _GEN_6573; // @[ICache.scala 169:30]
  wire  _GEN_8125 = uncached ? _GEN_2510 : _GEN_6574; // @[ICache.scala 169:30]
  wire  _GEN_8126 = uncached ? _GEN_3022 : _GEN_6575; // @[ICache.scala 169:30]
  wire  _GEN_8127 = uncached ? _GEN_2511 : _GEN_6576; // @[ICache.scala 169:30]
  wire  _GEN_8128 = uncached ? _GEN_3023 : _GEN_6577; // @[ICache.scala 169:30]
  wire  _GEN_8129 = uncached ? _GEN_2512 : _GEN_6578; // @[ICache.scala 169:30]
  wire  _GEN_8130 = uncached ? _GEN_3024 : _GEN_6579; // @[ICache.scala 169:30]
  wire  _GEN_8131 = uncached ? _GEN_2513 : _GEN_6580; // @[ICache.scala 169:30]
  wire  _GEN_8132 = uncached ? _GEN_3025 : _GEN_6581; // @[ICache.scala 169:30]
  wire  _GEN_8133 = uncached ? _GEN_2514 : _GEN_6582; // @[ICache.scala 169:30]
  wire  _GEN_8134 = uncached ? _GEN_3026 : _GEN_6583; // @[ICache.scala 169:30]
  wire  _GEN_8135 = uncached ? _GEN_2515 : _GEN_6584; // @[ICache.scala 169:30]
  wire  _GEN_8136 = uncached ? _GEN_3027 : _GEN_6585; // @[ICache.scala 169:30]
  wire  _GEN_8137 = uncached ? _GEN_2516 : _GEN_6586; // @[ICache.scala 169:30]
  wire  _GEN_8138 = uncached ? _GEN_3028 : _GEN_6587; // @[ICache.scala 169:30]
  wire  _GEN_8139 = uncached ? _GEN_2517 : _GEN_6588; // @[ICache.scala 169:30]
  wire  _GEN_8140 = uncached ? _GEN_3029 : _GEN_6589; // @[ICache.scala 169:30]
  wire  _GEN_8141 = uncached ? _GEN_2518 : _GEN_6590; // @[ICache.scala 169:30]
  wire  _GEN_8142 = uncached ? _GEN_3030 : _GEN_6591; // @[ICache.scala 169:30]
  wire  _GEN_8143 = uncached ? _GEN_2519 : _GEN_6592; // @[ICache.scala 169:30]
  wire  _GEN_8144 = uncached ? _GEN_3031 : _GEN_6593; // @[ICache.scala 169:30]
  wire  _GEN_8145 = uncached ? _GEN_2520 : _GEN_6594; // @[ICache.scala 169:30]
  wire  _GEN_8146 = uncached ? _GEN_3032 : _GEN_6595; // @[ICache.scala 169:30]
  wire  _GEN_8147 = uncached ? _GEN_2521 : _GEN_6596; // @[ICache.scala 169:30]
  wire  _GEN_8148 = uncached ? _GEN_3033 : _GEN_6597; // @[ICache.scala 169:30]
  wire  _GEN_8149 = uncached ? _GEN_2522 : _GEN_6598; // @[ICache.scala 169:30]
  wire  _GEN_8150 = uncached ? _GEN_3034 : _GEN_6599; // @[ICache.scala 169:30]
  wire  _GEN_8151 = uncached ? _GEN_2523 : _GEN_6600; // @[ICache.scala 169:30]
  wire  _GEN_8152 = uncached ? _GEN_3035 : _GEN_6601; // @[ICache.scala 169:30]
  wire  _GEN_8153 = uncached ? _GEN_2524 : _GEN_6602; // @[ICache.scala 169:30]
  wire  _GEN_8154 = uncached ? _GEN_3036 : _GEN_6603; // @[ICache.scala 169:30]
  wire  _GEN_8155 = uncached ? _GEN_2525 : _GEN_6604; // @[ICache.scala 169:30]
  wire  _GEN_8156 = uncached ? _GEN_3037 : _GEN_6605; // @[ICache.scala 169:30]
  wire  _GEN_8157 = uncached ? _GEN_2526 : _GEN_6606; // @[ICache.scala 169:30]
  wire  _GEN_8158 = uncached ? _GEN_3038 : _GEN_6607; // @[ICache.scala 169:30]
  wire  _GEN_8159 = uncached ? _GEN_2527 : _GEN_6608; // @[ICache.scala 169:30]
  wire  _GEN_8160 = uncached ? _GEN_3039 : _GEN_6609; // @[ICache.scala 169:30]
  wire  _GEN_8161 = uncached ? _GEN_2528 : _GEN_6610; // @[ICache.scala 169:30]
  wire  _GEN_8162 = uncached ? _GEN_3040 : _GEN_6611; // @[ICache.scala 169:30]
  wire  _GEN_8163 = uncached ? _GEN_2529 : _GEN_6612; // @[ICache.scala 169:30]
  wire  _GEN_8164 = uncached ? _GEN_3041 : _GEN_6613; // @[ICache.scala 169:30]
  wire  _GEN_8165 = uncached ? _GEN_2530 : _GEN_6614; // @[ICache.scala 169:30]
  wire  _GEN_8166 = uncached ? _GEN_3042 : _GEN_6615; // @[ICache.scala 169:30]
  wire  _GEN_8167 = uncached ? _GEN_2531 : _GEN_6616; // @[ICache.scala 169:30]
  wire  _GEN_8168 = uncached ? _GEN_3043 : _GEN_6617; // @[ICache.scala 169:30]
  wire  _GEN_8169 = uncached ? _GEN_2532 : _GEN_6618; // @[ICache.scala 169:30]
  wire  _GEN_8170 = uncached ? _GEN_3044 : _GEN_6619; // @[ICache.scala 169:30]
  wire  _GEN_8171 = uncached ? _GEN_2533 : _GEN_6620; // @[ICache.scala 169:30]
  wire  _GEN_8172 = uncached ? _GEN_3045 : _GEN_6621; // @[ICache.scala 169:30]
  wire  _GEN_8173 = uncached ? _GEN_2534 : _GEN_6622; // @[ICache.scala 169:30]
  wire  _GEN_8174 = uncached ? _GEN_3046 : _GEN_6623; // @[ICache.scala 169:30]
  wire  _GEN_8175 = uncached ? _GEN_2535 : _GEN_6624; // @[ICache.scala 169:30]
  wire  _GEN_8176 = uncached ? _GEN_3047 : _GEN_6625; // @[ICache.scala 169:30]
  wire  _GEN_8177 = uncached ? _GEN_2536 : _GEN_6626; // @[ICache.scala 169:30]
  wire  _GEN_8178 = uncached ? _GEN_3048 : _GEN_6627; // @[ICache.scala 169:30]
  wire  _GEN_8179 = uncached ? _GEN_2537 : _GEN_6628; // @[ICache.scala 169:30]
  wire  _GEN_8180 = uncached ? _GEN_3049 : _GEN_6629; // @[ICache.scala 169:30]
  wire  _GEN_8181 = uncached ? _GEN_2538 : _GEN_6630; // @[ICache.scala 169:30]
  wire  _GEN_8182 = uncached ? _GEN_3050 : _GEN_6631; // @[ICache.scala 169:30]
  wire  _GEN_8183 = uncached ? _GEN_2539 : _GEN_6632; // @[ICache.scala 169:30]
  wire  _GEN_8184 = uncached ? _GEN_3051 : _GEN_6633; // @[ICache.scala 169:30]
  wire  _GEN_8185 = uncached ? _GEN_2540 : _GEN_6634; // @[ICache.scala 169:30]
  wire  _GEN_8186 = uncached ? _GEN_3052 : _GEN_6635; // @[ICache.scala 169:30]
  wire  _GEN_8187 = uncached ? _GEN_2541 : _GEN_6636; // @[ICache.scala 169:30]
  wire  _GEN_8188 = uncached ? _GEN_3053 : _GEN_6637; // @[ICache.scala 169:30]
  wire  _GEN_8189 = uncached ? _GEN_2542 : _GEN_6638; // @[ICache.scala 169:30]
  wire  _GEN_8190 = uncached ? _GEN_3054 : _GEN_6639; // @[ICache.scala 169:30]
  wire  _GEN_8191 = uncached ? _GEN_2543 : _GEN_6640; // @[ICache.scala 169:30]
  wire  _GEN_8192 = uncached ? _GEN_3055 : _GEN_6641; // @[ICache.scala 169:30]
  wire  _GEN_8193 = uncached ? _GEN_2544 : _GEN_6642; // @[ICache.scala 169:30]
  wire  _GEN_8194 = uncached ? _GEN_3056 : _GEN_6643; // @[ICache.scala 169:30]
  wire  _GEN_8195 = uncached ? _GEN_2545 : _GEN_6644; // @[ICache.scala 169:30]
  wire  _GEN_8196 = uncached ? _GEN_3057 : _GEN_6645; // @[ICache.scala 169:30]
  wire  _GEN_8197 = uncached ? _GEN_2546 : _GEN_6646; // @[ICache.scala 169:30]
  wire  _GEN_8198 = uncached ? _GEN_3058 : _GEN_6647; // @[ICache.scala 169:30]
  wire  _GEN_8199 = uncached ? _GEN_2547 : _GEN_6648; // @[ICache.scala 169:30]
  wire  _GEN_8200 = uncached ? _GEN_3059 : _GEN_6649; // @[ICache.scala 169:30]
  wire  _GEN_8201 = uncached ? _GEN_2548 : _GEN_6650; // @[ICache.scala 169:30]
  wire  _GEN_8202 = uncached ? _GEN_3060 : _GEN_6651; // @[ICache.scala 169:30]
  wire  _GEN_8203 = uncached ? _GEN_2549 : _GEN_6652; // @[ICache.scala 169:30]
  wire  _GEN_8204 = uncached ? _GEN_3061 : _GEN_6653; // @[ICache.scala 169:30]
  wire  _GEN_8205 = uncached ? _GEN_2550 : _GEN_6654; // @[ICache.scala 169:30]
  wire  _GEN_8206 = uncached ? _GEN_3062 : _GEN_6655; // @[ICache.scala 169:30]
  wire  _GEN_8207 = uncached ? _GEN_2551 : _GEN_6656; // @[ICache.scala 169:30]
  wire  _GEN_8208 = uncached ? _GEN_3063 : _GEN_6657; // @[ICache.scala 169:30]
  wire  _GEN_8209 = uncached ? _GEN_2552 : _GEN_6658; // @[ICache.scala 169:30]
  wire  _GEN_8210 = uncached ? _GEN_3064 : _GEN_6659; // @[ICache.scala 169:30]
  wire  _GEN_8211 = uncached ? _GEN_2553 : _GEN_6660; // @[ICache.scala 169:30]
  wire  _GEN_8212 = uncached ? _GEN_3065 : _GEN_6661; // @[ICache.scala 169:30]
  wire  _GEN_8213 = uncached ? _GEN_2554 : _GEN_6662; // @[ICache.scala 169:30]
  wire  _GEN_8214 = uncached ? _GEN_3066 : _GEN_6663; // @[ICache.scala 169:30]
  wire  _GEN_8215 = uncached ? _GEN_2555 : _GEN_6664; // @[ICache.scala 169:30]
  wire  _GEN_8216 = uncached ? _GEN_3067 : _GEN_6665; // @[ICache.scala 169:30]
  wire  _GEN_8217 = uncached ? _GEN_2556 : _GEN_6666; // @[ICache.scala 169:30]
  wire  _GEN_8218 = uncached ? _GEN_3068 : _GEN_6667; // @[ICache.scala 169:30]
  wire  _GEN_8219 = uncached ? _GEN_2557 : _GEN_6668; // @[ICache.scala 169:30]
  wire  _GEN_8220 = uncached ? _GEN_3069 : _GEN_6669; // @[ICache.scala 169:30]
  wire  _GEN_8221 = uncached ? _GEN_2558 : _GEN_6670; // @[ICache.scala 169:30]
  wire  _GEN_8222 = uncached ? _GEN_3070 : _GEN_6671; // @[ICache.scala 169:30]
  wire  _GEN_8223 = uncached ? _GEN_2559 : _GEN_6672; // @[ICache.scala 169:30]
  wire  _GEN_8224 = uncached ? _GEN_3071 : _GEN_6673; // @[ICache.scala 169:30]
  wire  _GEN_8225 = uncached ? _GEN_2560 : _GEN_6674; // @[ICache.scala 169:30]
  wire  _GEN_8226 = uncached ? _GEN_3072 : _GEN_6675; // @[ICache.scala 169:30]
  wire  _GEN_8227 = uncached ? _GEN_2561 : _GEN_6676; // @[ICache.scala 169:30]
  wire  _GEN_8228 = uncached ? _GEN_3073 : _GEN_6677; // @[ICache.scala 169:30]
  wire  _GEN_8229 = uncached ? _GEN_2562 : _GEN_6678; // @[ICache.scala 169:30]
  wire  _GEN_8230 = uncached ? _GEN_3074 : _GEN_6679; // @[ICache.scala 169:30]
  wire  _GEN_8231 = uncached ? _GEN_2563 : _GEN_6680; // @[ICache.scala 169:30]
  wire  _GEN_8232 = uncached ? _GEN_3075 : _GEN_6681; // @[ICache.scala 169:30]
  wire  _GEN_8233 = uncached ? _GEN_2564 : _GEN_6682; // @[ICache.scala 169:30]
  wire  _GEN_8234 = uncached ? _GEN_3076 : _GEN_6683; // @[ICache.scala 169:30]
  wire [4:0] _GEN_8235 = uncached ? axi_cnt : _GEN_6684; // @[ICache.scala 109:24 169:30]
  wire  _GEN_8236 = uncached ? meta_0_lru : _GEN_6685; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8237 = uncached ? meta_1_lru : _GEN_6686; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8238 = uncached ? meta_2_lru : _GEN_6687; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8239 = uncached ? meta_3_lru : _GEN_6688; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8240 = uncached ? meta_4_lru : _GEN_6689; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8241 = uncached ? meta_5_lru : _GEN_6690; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8242 = uncached ? meta_6_lru : _GEN_6691; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8243 = uncached ? meta_7_lru : _GEN_6692; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8244 = uncached ? meta_8_lru : _GEN_6693; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8245 = uncached ? meta_9_lru : _GEN_6694; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8246 = uncached ? meta_10_lru : _GEN_6695; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8247 = uncached ? meta_11_lru : _GEN_6696; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8248 = uncached ? meta_12_lru : _GEN_6697; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8249 = uncached ? meta_13_lru : _GEN_6698; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8250 = uncached ? meta_14_lru : _GEN_6699; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8251 = uncached ? meta_15_lru : _GEN_6700; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8252 = uncached ? meta_16_lru : _GEN_6701; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8253 = uncached ? meta_17_lru : _GEN_6702; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8254 = uncached ? meta_18_lru : _GEN_6703; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8255 = uncached ? meta_19_lru : _GEN_6704; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8256 = uncached ? meta_20_lru : _GEN_6705; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8257 = uncached ? meta_21_lru : _GEN_6706; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8258 = uncached ? meta_22_lru : _GEN_6707; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8259 = uncached ? meta_23_lru : _GEN_6708; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8260 = uncached ? meta_24_lru : _GEN_6709; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8261 = uncached ? meta_25_lru : _GEN_6710; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8262 = uncached ? meta_26_lru : _GEN_6711; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8263 = uncached ? meta_27_lru : _GEN_6712; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8264 = uncached ? meta_28_lru : _GEN_6713; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8265 = uncached ? meta_29_lru : _GEN_6714; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8266 = uncached ? meta_30_lru : _GEN_6715; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8267 = uncached ? meta_31_lru : _GEN_6716; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8268 = uncached ? meta_32_lru : _GEN_6717; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8269 = uncached ? meta_33_lru : _GEN_6718; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8270 = uncached ? meta_34_lru : _GEN_6719; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8271 = uncached ? meta_35_lru : _GEN_6720; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8272 = uncached ? meta_36_lru : _GEN_6721; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8273 = uncached ? meta_37_lru : _GEN_6722; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8274 = uncached ? meta_38_lru : _GEN_6723; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8275 = uncached ? meta_39_lru : _GEN_6724; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8276 = uncached ? meta_40_lru : _GEN_6725; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8277 = uncached ? meta_41_lru : _GEN_6726; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8278 = uncached ? meta_42_lru : _GEN_6727; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8279 = uncached ? meta_43_lru : _GEN_6728; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8280 = uncached ? meta_44_lru : _GEN_6729; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8281 = uncached ? meta_45_lru : _GEN_6730; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8282 = uncached ? meta_46_lru : _GEN_6731; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8283 = uncached ? meta_47_lru : _GEN_6732; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8284 = uncached ? meta_48_lru : _GEN_6733; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8285 = uncached ? meta_49_lru : _GEN_6734; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8286 = uncached ? meta_50_lru : _GEN_6735; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8287 = uncached ? meta_51_lru : _GEN_6736; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8288 = uncached ? meta_52_lru : _GEN_6737; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8289 = uncached ? meta_53_lru : _GEN_6738; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8290 = uncached ? meta_54_lru : _GEN_6739; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8291 = uncached ? meta_55_lru : _GEN_6740; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8292 = uncached ? meta_56_lru : _GEN_6741; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8293 = uncached ? meta_57_lru : _GEN_6742; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8294 = uncached ? meta_58_lru : _GEN_6743; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8295 = uncached ? meta_59_lru : _GEN_6744; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8296 = uncached ? meta_60_lru : _GEN_6745; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8297 = uncached ? meta_61_lru : _GEN_6746; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8298 = uncached ? meta_62_lru : _GEN_6747; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8299 = uncached ? meta_63_lru : _GEN_6748; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8300 = uncached ? meta_64_lru : _GEN_6749; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8301 = uncached ? meta_65_lru : _GEN_6750; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8302 = uncached ? meta_66_lru : _GEN_6751; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8303 = uncached ? meta_67_lru : _GEN_6752; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8304 = uncached ? meta_68_lru : _GEN_6753; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8305 = uncached ? meta_69_lru : _GEN_6754; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8306 = uncached ? meta_70_lru : _GEN_6755; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8307 = uncached ? meta_71_lru : _GEN_6756; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8308 = uncached ? meta_72_lru : _GEN_6757; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8309 = uncached ? meta_73_lru : _GEN_6758; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8310 = uncached ? meta_74_lru : _GEN_6759; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8311 = uncached ? meta_75_lru : _GEN_6760; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8312 = uncached ? meta_76_lru : _GEN_6761; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8313 = uncached ? meta_77_lru : _GEN_6762; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8314 = uncached ? meta_78_lru : _GEN_6763; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8315 = uncached ? meta_79_lru : _GEN_6764; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8316 = uncached ? meta_80_lru : _GEN_6765; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8317 = uncached ? meta_81_lru : _GEN_6766; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8318 = uncached ? meta_82_lru : _GEN_6767; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8319 = uncached ? meta_83_lru : _GEN_6768; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8320 = uncached ? meta_84_lru : _GEN_6769; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8321 = uncached ? meta_85_lru : _GEN_6770; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8322 = uncached ? meta_86_lru : _GEN_6771; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8323 = uncached ? meta_87_lru : _GEN_6772; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8324 = uncached ? meta_88_lru : _GEN_6773; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8325 = uncached ? meta_89_lru : _GEN_6774; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8326 = uncached ? meta_90_lru : _GEN_6775; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8327 = uncached ? meta_91_lru : _GEN_6776; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8328 = uncached ? meta_92_lru : _GEN_6777; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8329 = uncached ? meta_93_lru : _GEN_6778; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8330 = uncached ? meta_94_lru : _GEN_6779; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8331 = uncached ? meta_95_lru : _GEN_6780; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8332 = uncached ? meta_96_lru : _GEN_6781; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8333 = uncached ? meta_97_lru : _GEN_6782; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8334 = uncached ? meta_98_lru : _GEN_6783; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8335 = uncached ? meta_99_lru : _GEN_6784; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8336 = uncached ? meta_100_lru : _GEN_6785; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8337 = uncached ? meta_101_lru : _GEN_6786; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8338 = uncached ? meta_102_lru : _GEN_6787; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8339 = uncached ? meta_103_lru : _GEN_6788; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8340 = uncached ? meta_104_lru : _GEN_6789; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8341 = uncached ? meta_105_lru : _GEN_6790; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8342 = uncached ? meta_106_lru : _GEN_6791; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8343 = uncached ? meta_107_lru : _GEN_6792; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8344 = uncached ? meta_108_lru : _GEN_6793; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8345 = uncached ? meta_109_lru : _GEN_6794; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8346 = uncached ? meta_110_lru : _GEN_6795; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8347 = uncached ? meta_111_lru : _GEN_6796; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8348 = uncached ? meta_112_lru : _GEN_6797; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8349 = uncached ? meta_113_lru : _GEN_6798; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8350 = uncached ? meta_114_lru : _GEN_6799; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8351 = uncached ? meta_115_lru : _GEN_6800; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8352 = uncached ? meta_116_lru : _GEN_6801; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8353 = uncached ? meta_117_lru : _GEN_6802; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8354 = uncached ? meta_118_lru : _GEN_6803; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8355 = uncached ? meta_119_lru : _GEN_6804; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8356 = uncached ? meta_120_lru : _GEN_6805; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8357 = uncached ? meta_121_lru : _GEN_6806; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8358 = uncached ? meta_122_lru : _GEN_6807; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8359 = uncached ? meta_123_lru : _GEN_6808; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8360 = uncached ? meta_124_lru : _GEN_6809; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8361 = uncached ? meta_125_lru : _GEN_6810; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8362 = uncached ? meta_126_lru : _GEN_6811; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8363 = uncached ? meta_127_lru : _GEN_6812; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8364 = uncached ? meta_128_lru : _GEN_6813; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8365 = uncached ? meta_129_lru : _GEN_6814; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8366 = uncached ? meta_130_lru : _GEN_6815; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8367 = uncached ? meta_131_lru : _GEN_6816; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8368 = uncached ? meta_132_lru : _GEN_6817; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8369 = uncached ? meta_133_lru : _GEN_6818; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8370 = uncached ? meta_134_lru : _GEN_6819; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8371 = uncached ? meta_135_lru : _GEN_6820; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8372 = uncached ? meta_136_lru : _GEN_6821; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8373 = uncached ? meta_137_lru : _GEN_6822; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8374 = uncached ? meta_138_lru : _GEN_6823; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8375 = uncached ? meta_139_lru : _GEN_6824; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8376 = uncached ? meta_140_lru : _GEN_6825; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8377 = uncached ? meta_141_lru : _GEN_6826; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8378 = uncached ? meta_142_lru : _GEN_6827; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8379 = uncached ? meta_143_lru : _GEN_6828; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8380 = uncached ? meta_144_lru : _GEN_6829; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8381 = uncached ? meta_145_lru : _GEN_6830; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8382 = uncached ? meta_146_lru : _GEN_6831; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8383 = uncached ? meta_147_lru : _GEN_6832; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8384 = uncached ? meta_148_lru : _GEN_6833; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8385 = uncached ? meta_149_lru : _GEN_6834; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8386 = uncached ? meta_150_lru : _GEN_6835; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8387 = uncached ? meta_151_lru : _GEN_6836; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8388 = uncached ? meta_152_lru : _GEN_6837; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8389 = uncached ? meta_153_lru : _GEN_6838; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8390 = uncached ? meta_154_lru : _GEN_6839; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8391 = uncached ? meta_155_lru : _GEN_6840; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8392 = uncached ? meta_156_lru : _GEN_6841; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8393 = uncached ? meta_157_lru : _GEN_6842; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8394 = uncached ? meta_158_lru : _GEN_6843; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8395 = uncached ? meta_159_lru : _GEN_6844; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8396 = uncached ? meta_160_lru : _GEN_6845; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8397 = uncached ? meta_161_lru : _GEN_6846; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8398 = uncached ? meta_162_lru : _GEN_6847; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8399 = uncached ? meta_163_lru : _GEN_6848; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8400 = uncached ? meta_164_lru : _GEN_6849; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8401 = uncached ? meta_165_lru : _GEN_6850; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8402 = uncached ? meta_166_lru : _GEN_6851; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8403 = uncached ? meta_167_lru : _GEN_6852; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8404 = uncached ? meta_168_lru : _GEN_6853; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8405 = uncached ? meta_169_lru : _GEN_6854; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8406 = uncached ? meta_170_lru : _GEN_6855; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8407 = uncached ? meta_171_lru : _GEN_6856; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8408 = uncached ? meta_172_lru : _GEN_6857; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8409 = uncached ? meta_173_lru : _GEN_6858; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8410 = uncached ? meta_174_lru : _GEN_6859; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8411 = uncached ? meta_175_lru : _GEN_6860; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8412 = uncached ? meta_176_lru : _GEN_6861; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8413 = uncached ? meta_177_lru : _GEN_6862; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8414 = uncached ? meta_178_lru : _GEN_6863; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8415 = uncached ? meta_179_lru : _GEN_6864; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8416 = uncached ? meta_180_lru : _GEN_6865; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8417 = uncached ? meta_181_lru : _GEN_6866; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8418 = uncached ? meta_182_lru : _GEN_6867; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8419 = uncached ? meta_183_lru : _GEN_6868; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8420 = uncached ? meta_184_lru : _GEN_6869; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8421 = uncached ? meta_185_lru : _GEN_6870; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8422 = uncached ? meta_186_lru : _GEN_6871; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8423 = uncached ? meta_187_lru : _GEN_6872; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8424 = uncached ? meta_188_lru : _GEN_6873; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8425 = uncached ? meta_189_lru : _GEN_6874; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8426 = uncached ? meta_190_lru : _GEN_6875; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8427 = uncached ? meta_191_lru : _GEN_6876; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8428 = uncached ? meta_192_lru : _GEN_6877; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8429 = uncached ? meta_193_lru : _GEN_6878; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8430 = uncached ? meta_194_lru : _GEN_6879; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8431 = uncached ? meta_195_lru : _GEN_6880; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8432 = uncached ? meta_196_lru : _GEN_6881; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8433 = uncached ? meta_197_lru : _GEN_6882; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8434 = uncached ? meta_198_lru : _GEN_6883; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8435 = uncached ? meta_199_lru : _GEN_6884; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8436 = uncached ? meta_200_lru : _GEN_6885; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8437 = uncached ? meta_201_lru : _GEN_6886; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8438 = uncached ? meta_202_lru : _GEN_6887; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8439 = uncached ? meta_203_lru : _GEN_6888; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8440 = uncached ? meta_204_lru : _GEN_6889; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8441 = uncached ? meta_205_lru : _GEN_6890; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8442 = uncached ? meta_206_lru : _GEN_6891; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8443 = uncached ? meta_207_lru : _GEN_6892; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8444 = uncached ? meta_208_lru : _GEN_6893; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8445 = uncached ? meta_209_lru : _GEN_6894; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8446 = uncached ? meta_210_lru : _GEN_6895; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8447 = uncached ? meta_211_lru : _GEN_6896; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8448 = uncached ? meta_212_lru : _GEN_6897; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8449 = uncached ? meta_213_lru : _GEN_6898; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8450 = uncached ? meta_214_lru : _GEN_6899; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8451 = uncached ? meta_215_lru : _GEN_6900; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8452 = uncached ? meta_216_lru : _GEN_6901; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8453 = uncached ? meta_217_lru : _GEN_6902; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8454 = uncached ? meta_218_lru : _GEN_6903; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8455 = uncached ? meta_219_lru : _GEN_6904; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8456 = uncached ? meta_220_lru : _GEN_6905; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8457 = uncached ? meta_221_lru : _GEN_6906; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8458 = uncached ? meta_222_lru : _GEN_6907; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8459 = uncached ? meta_223_lru : _GEN_6908; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8460 = uncached ? meta_224_lru : _GEN_6909; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8461 = uncached ? meta_225_lru : _GEN_6910; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8462 = uncached ? meta_226_lru : _GEN_6911; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8463 = uncached ? meta_227_lru : _GEN_6912; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8464 = uncached ? meta_228_lru : _GEN_6913; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8465 = uncached ? meta_229_lru : _GEN_6914; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8466 = uncached ? meta_230_lru : _GEN_6915; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8467 = uncached ? meta_231_lru : _GEN_6916; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8468 = uncached ? meta_232_lru : _GEN_6917; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8469 = uncached ? meta_233_lru : _GEN_6918; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8470 = uncached ? meta_234_lru : _GEN_6919; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8471 = uncached ? meta_235_lru : _GEN_6920; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8472 = uncached ? meta_236_lru : _GEN_6921; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8473 = uncached ? meta_237_lru : _GEN_6922; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8474 = uncached ? meta_238_lru : _GEN_6923; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8475 = uncached ? meta_239_lru : _GEN_6924; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8476 = uncached ? meta_240_lru : _GEN_6925; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8477 = uncached ? meta_241_lru : _GEN_6926; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8478 = uncached ? meta_242_lru : _GEN_6927; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8479 = uncached ? meta_243_lru : _GEN_6928; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8480 = uncached ? meta_244_lru : _GEN_6929; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8481 = uncached ? meta_245_lru : _GEN_6930; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8482 = uncached ? meta_246_lru : _GEN_6931; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8483 = uncached ? meta_247_lru : _GEN_6932; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8484 = uncached ? meta_248_lru : _GEN_6933; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8485 = uncached ? meta_249_lru : _GEN_6934; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8486 = uncached ? meta_250_lru : _GEN_6935; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8487 = uncached ? meta_251_lru : _GEN_6936; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8488 = uncached ? meta_252_lru : _GEN_6937; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8489 = uncached ? meta_253_lru : _GEN_6938; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8490 = uncached ? meta_254_lru : _GEN_6939; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8491 = uncached ? meta_255_lru : _GEN_6940; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8492 = uncached ? meta_256_lru : _GEN_6941; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8493 = uncached ? meta_257_lru : _GEN_6942; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8494 = uncached ? meta_258_lru : _GEN_6943; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8495 = uncached ? meta_259_lru : _GEN_6944; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8496 = uncached ? meta_260_lru : _GEN_6945; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8497 = uncached ? meta_261_lru : _GEN_6946; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8498 = uncached ? meta_262_lru : _GEN_6947; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8499 = uncached ? meta_263_lru : _GEN_6948; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8500 = uncached ? meta_264_lru : _GEN_6949; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8501 = uncached ? meta_265_lru : _GEN_6950; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8502 = uncached ? meta_266_lru : _GEN_6951; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8503 = uncached ? meta_267_lru : _GEN_6952; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8504 = uncached ? meta_268_lru : _GEN_6953; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8505 = uncached ? meta_269_lru : _GEN_6954; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8506 = uncached ? meta_270_lru : _GEN_6955; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8507 = uncached ? meta_271_lru : _GEN_6956; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8508 = uncached ? meta_272_lru : _GEN_6957; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8509 = uncached ? meta_273_lru : _GEN_6958; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8510 = uncached ? meta_274_lru : _GEN_6959; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8511 = uncached ? meta_275_lru : _GEN_6960; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8512 = uncached ? meta_276_lru : _GEN_6961; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8513 = uncached ? meta_277_lru : _GEN_6962; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8514 = uncached ? meta_278_lru : _GEN_6963; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8515 = uncached ? meta_279_lru : _GEN_6964; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8516 = uncached ? meta_280_lru : _GEN_6965; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8517 = uncached ? meta_281_lru : _GEN_6966; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8518 = uncached ? meta_282_lru : _GEN_6967; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8519 = uncached ? meta_283_lru : _GEN_6968; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8520 = uncached ? meta_284_lru : _GEN_6969; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8521 = uncached ? meta_285_lru : _GEN_6970; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8522 = uncached ? meta_286_lru : _GEN_6971; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8523 = uncached ? meta_287_lru : _GEN_6972; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8524 = uncached ? meta_288_lru : _GEN_6973; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8525 = uncached ? meta_289_lru : _GEN_6974; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8526 = uncached ? meta_290_lru : _GEN_6975; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8527 = uncached ? meta_291_lru : _GEN_6976; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8528 = uncached ? meta_292_lru : _GEN_6977; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8529 = uncached ? meta_293_lru : _GEN_6978; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8530 = uncached ? meta_294_lru : _GEN_6979; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8531 = uncached ? meta_295_lru : _GEN_6980; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8532 = uncached ? meta_296_lru : _GEN_6981; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8533 = uncached ? meta_297_lru : _GEN_6982; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8534 = uncached ? meta_298_lru : _GEN_6983; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8535 = uncached ? meta_299_lru : _GEN_6984; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8536 = uncached ? meta_300_lru : _GEN_6985; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8537 = uncached ? meta_301_lru : _GEN_6986; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8538 = uncached ? meta_302_lru : _GEN_6987; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8539 = uncached ? meta_303_lru : _GEN_6988; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8540 = uncached ? meta_304_lru : _GEN_6989; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8541 = uncached ? meta_305_lru : _GEN_6990; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8542 = uncached ? meta_306_lru : _GEN_6991; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8543 = uncached ? meta_307_lru : _GEN_6992; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8544 = uncached ? meta_308_lru : _GEN_6993; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8545 = uncached ? meta_309_lru : _GEN_6994; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8546 = uncached ? meta_310_lru : _GEN_6995; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8547 = uncached ? meta_311_lru : _GEN_6996; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8548 = uncached ? meta_312_lru : _GEN_6997; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8549 = uncached ? meta_313_lru : _GEN_6998; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8550 = uncached ? meta_314_lru : _GEN_6999; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8551 = uncached ? meta_315_lru : _GEN_7000; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8552 = uncached ? meta_316_lru : _GEN_7001; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8553 = uncached ? meta_317_lru : _GEN_7002; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8554 = uncached ? meta_318_lru : _GEN_7003; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8555 = uncached ? meta_319_lru : _GEN_7004; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8556 = uncached ? meta_320_lru : _GEN_7005; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8557 = uncached ? meta_321_lru : _GEN_7006; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8558 = uncached ? meta_322_lru : _GEN_7007; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8559 = uncached ? meta_323_lru : _GEN_7008; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8560 = uncached ? meta_324_lru : _GEN_7009; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8561 = uncached ? meta_325_lru : _GEN_7010; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8562 = uncached ? meta_326_lru : _GEN_7011; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8563 = uncached ? meta_327_lru : _GEN_7012; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8564 = uncached ? meta_328_lru : _GEN_7013; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8565 = uncached ? meta_329_lru : _GEN_7014; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8566 = uncached ? meta_330_lru : _GEN_7015; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8567 = uncached ? meta_331_lru : _GEN_7016; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8568 = uncached ? meta_332_lru : _GEN_7017; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8569 = uncached ? meta_333_lru : _GEN_7018; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8570 = uncached ? meta_334_lru : _GEN_7019; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8571 = uncached ? meta_335_lru : _GEN_7020; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8572 = uncached ? meta_336_lru : _GEN_7021; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8573 = uncached ? meta_337_lru : _GEN_7022; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8574 = uncached ? meta_338_lru : _GEN_7023; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8575 = uncached ? meta_339_lru : _GEN_7024; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8576 = uncached ? meta_340_lru : _GEN_7025; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8577 = uncached ? meta_341_lru : _GEN_7026; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8578 = uncached ? meta_342_lru : _GEN_7027; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8579 = uncached ? meta_343_lru : _GEN_7028; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8580 = uncached ? meta_344_lru : _GEN_7029; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8581 = uncached ? meta_345_lru : _GEN_7030; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8582 = uncached ? meta_346_lru : _GEN_7031; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8583 = uncached ? meta_347_lru : _GEN_7032; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8584 = uncached ? meta_348_lru : _GEN_7033; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8585 = uncached ? meta_349_lru : _GEN_7034; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8586 = uncached ? meta_350_lru : _GEN_7035; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8587 = uncached ? meta_351_lru : _GEN_7036; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8588 = uncached ? meta_352_lru : _GEN_7037; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8589 = uncached ? meta_353_lru : _GEN_7038; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8590 = uncached ? meta_354_lru : _GEN_7039; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8591 = uncached ? meta_355_lru : _GEN_7040; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8592 = uncached ? meta_356_lru : _GEN_7041; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8593 = uncached ? meta_357_lru : _GEN_7042; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8594 = uncached ? meta_358_lru : _GEN_7043; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8595 = uncached ? meta_359_lru : _GEN_7044; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8596 = uncached ? meta_360_lru : _GEN_7045; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8597 = uncached ? meta_361_lru : _GEN_7046; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8598 = uncached ? meta_362_lru : _GEN_7047; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8599 = uncached ? meta_363_lru : _GEN_7048; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8600 = uncached ? meta_364_lru : _GEN_7049; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8601 = uncached ? meta_365_lru : _GEN_7050; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8602 = uncached ? meta_366_lru : _GEN_7051; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8603 = uncached ? meta_367_lru : _GEN_7052; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8604 = uncached ? meta_368_lru : _GEN_7053; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8605 = uncached ? meta_369_lru : _GEN_7054; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8606 = uncached ? meta_370_lru : _GEN_7055; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8607 = uncached ? meta_371_lru : _GEN_7056; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8608 = uncached ? meta_372_lru : _GEN_7057; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8609 = uncached ? meta_373_lru : _GEN_7058; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8610 = uncached ? meta_374_lru : _GEN_7059; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8611 = uncached ? meta_375_lru : _GEN_7060; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8612 = uncached ? meta_376_lru : _GEN_7061; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8613 = uncached ? meta_377_lru : _GEN_7062; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8614 = uncached ? meta_378_lru : _GEN_7063; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8615 = uncached ? meta_379_lru : _GEN_7064; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8616 = uncached ? meta_380_lru : _GEN_7065; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8617 = uncached ? meta_381_lru : _GEN_7066; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8618 = uncached ? meta_382_lru : _GEN_7067; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8619 = uncached ? meta_383_lru : _GEN_7068; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8620 = uncached ? meta_384_lru : _GEN_7069; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8621 = uncached ? meta_385_lru : _GEN_7070; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8622 = uncached ? meta_386_lru : _GEN_7071; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8623 = uncached ? meta_387_lru : _GEN_7072; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8624 = uncached ? meta_388_lru : _GEN_7073; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8625 = uncached ? meta_389_lru : _GEN_7074; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8626 = uncached ? meta_390_lru : _GEN_7075; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8627 = uncached ? meta_391_lru : _GEN_7076; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8628 = uncached ? meta_392_lru : _GEN_7077; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8629 = uncached ? meta_393_lru : _GEN_7078; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8630 = uncached ? meta_394_lru : _GEN_7079; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8631 = uncached ? meta_395_lru : _GEN_7080; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8632 = uncached ? meta_396_lru : _GEN_7081; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8633 = uncached ? meta_397_lru : _GEN_7082; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8634 = uncached ? meta_398_lru : _GEN_7083; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8635 = uncached ? meta_399_lru : _GEN_7084; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8636 = uncached ? meta_400_lru : _GEN_7085; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8637 = uncached ? meta_401_lru : _GEN_7086; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8638 = uncached ? meta_402_lru : _GEN_7087; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8639 = uncached ? meta_403_lru : _GEN_7088; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8640 = uncached ? meta_404_lru : _GEN_7089; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8641 = uncached ? meta_405_lru : _GEN_7090; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8642 = uncached ? meta_406_lru : _GEN_7091; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8643 = uncached ? meta_407_lru : _GEN_7092; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8644 = uncached ? meta_408_lru : _GEN_7093; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8645 = uncached ? meta_409_lru : _GEN_7094; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8646 = uncached ? meta_410_lru : _GEN_7095; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8647 = uncached ? meta_411_lru : _GEN_7096; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8648 = uncached ? meta_412_lru : _GEN_7097; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8649 = uncached ? meta_413_lru : _GEN_7098; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8650 = uncached ? meta_414_lru : _GEN_7099; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8651 = uncached ? meta_415_lru : _GEN_7100; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8652 = uncached ? meta_416_lru : _GEN_7101; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8653 = uncached ? meta_417_lru : _GEN_7102; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8654 = uncached ? meta_418_lru : _GEN_7103; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8655 = uncached ? meta_419_lru : _GEN_7104; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8656 = uncached ? meta_420_lru : _GEN_7105; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8657 = uncached ? meta_421_lru : _GEN_7106; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8658 = uncached ? meta_422_lru : _GEN_7107; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8659 = uncached ? meta_423_lru : _GEN_7108; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8660 = uncached ? meta_424_lru : _GEN_7109; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8661 = uncached ? meta_425_lru : _GEN_7110; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8662 = uncached ? meta_426_lru : _GEN_7111; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8663 = uncached ? meta_427_lru : _GEN_7112; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8664 = uncached ? meta_428_lru : _GEN_7113; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8665 = uncached ? meta_429_lru : _GEN_7114; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8666 = uncached ? meta_430_lru : _GEN_7115; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8667 = uncached ? meta_431_lru : _GEN_7116; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8668 = uncached ? meta_432_lru : _GEN_7117; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8669 = uncached ? meta_433_lru : _GEN_7118; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8670 = uncached ? meta_434_lru : _GEN_7119; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8671 = uncached ? meta_435_lru : _GEN_7120; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8672 = uncached ? meta_436_lru : _GEN_7121; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8673 = uncached ? meta_437_lru : _GEN_7122; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8674 = uncached ? meta_438_lru : _GEN_7123; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8675 = uncached ? meta_439_lru : _GEN_7124; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8676 = uncached ? meta_440_lru : _GEN_7125; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8677 = uncached ? meta_441_lru : _GEN_7126; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8678 = uncached ? meta_442_lru : _GEN_7127; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8679 = uncached ? meta_443_lru : _GEN_7128; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8680 = uncached ? meta_444_lru : _GEN_7129; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8681 = uncached ? meta_445_lru : _GEN_7130; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8682 = uncached ? meta_446_lru : _GEN_7131; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8683 = uncached ? meta_447_lru : _GEN_7132; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8684 = uncached ? meta_448_lru : _GEN_7133; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8685 = uncached ? meta_449_lru : _GEN_7134; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8686 = uncached ? meta_450_lru : _GEN_7135; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8687 = uncached ? meta_451_lru : _GEN_7136; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8688 = uncached ? meta_452_lru : _GEN_7137; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8689 = uncached ? meta_453_lru : _GEN_7138; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8690 = uncached ? meta_454_lru : _GEN_7139; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8691 = uncached ? meta_455_lru : _GEN_7140; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8692 = uncached ? meta_456_lru : _GEN_7141; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8693 = uncached ? meta_457_lru : _GEN_7142; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8694 = uncached ? meta_458_lru : _GEN_7143; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8695 = uncached ? meta_459_lru : _GEN_7144; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8696 = uncached ? meta_460_lru : _GEN_7145; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8697 = uncached ? meta_461_lru : _GEN_7146; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8698 = uncached ? meta_462_lru : _GEN_7147; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8699 = uncached ? meta_463_lru : _GEN_7148; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8700 = uncached ? meta_464_lru : _GEN_7149; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8701 = uncached ? meta_465_lru : _GEN_7150; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8702 = uncached ? meta_466_lru : _GEN_7151; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8703 = uncached ? meta_467_lru : _GEN_7152; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8704 = uncached ? meta_468_lru : _GEN_7153; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8705 = uncached ? meta_469_lru : _GEN_7154; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8706 = uncached ? meta_470_lru : _GEN_7155; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8707 = uncached ? meta_471_lru : _GEN_7156; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8708 = uncached ? meta_472_lru : _GEN_7157; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8709 = uncached ? meta_473_lru : _GEN_7158; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8710 = uncached ? meta_474_lru : _GEN_7159; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8711 = uncached ? meta_475_lru : _GEN_7160; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8712 = uncached ? meta_476_lru : _GEN_7161; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8713 = uncached ? meta_477_lru : _GEN_7162; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8714 = uncached ? meta_478_lru : _GEN_7163; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8715 = uncached ? meta_479_lru : _GEN_7164; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8716 = uncached ? meta_480_lru : _GEN_7165; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8717 = uncached ? meta_481_lru : _GEN_7166; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8718 = uncached ? meta_482_lru : _GEN_7167; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8719 = uncached ? meta_483_lru : _GEN_7168; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8720 = uncached ? meta_484_lru : _GEN_7169; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8721 = uncached ? meta_485_lru : _GEN_7170; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8722 = uncached ? meta_486_lru : _GEN_7171; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8723 = uncached ? meta_487_lru : _GEN_7172; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8724 = uncached ? meta_488_lru : _GEN_7173; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8725 = uncached ? meta_489_lru : _GEN_7174; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8726 = uncached ? meta_490_lru : _GEN_7175; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8727 = uncached ? meta_491_lru : _GEN_7176; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8728 = uncached ? meta_492_lru : _GEN_7177; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8729 = uncached ? meta_493_lru : _GEN_7178; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8730 = uncached ? meta_494_lru : _GEN_7179; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8731 = uncached ? meta_495_lru : _GEN_7180; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8732 = uncached ? meta_496_lru : _GEN_7181; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8733 = uncached ? meta_497_lru : _GEN_7182; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8734 = uncached ? meta_498_lru : _GEN_7183; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8735 = uncached ? meta_499_lru : _GEN_7184; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8736 = uncached ? meta_500_lru : _GEN_7185; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8737 = uncached ? meta_501_lru : _GEN_7186; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8738 = uncached ? meta_502_lru : _GEN_7187; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8739 = uncached ? meta_503_lru : _GEN_7188; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8740 = uncached ? meta_504_lru : _GEN_7189; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8741 = uncached ? meta_505_lru : _GEN_7190; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8742 = uncached ? meta_506_lru : _GEN_7191; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8743 = uncached ? meta_507_lru : _GEN_7192; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8744 = uncached ? meta_508_lru : _GEN_7193; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8745 = uncached ? meta_509_lru : _GEN_7194; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8746 = uncached ? meta_510_lru : _GEN_7195; // @[ICache.scala 169:30 34:21]
  wire  _GEN_8747 = uncached ? meta_511_lru : _GEN_7196; // @[ICache.scala 169:30 34:21]
  wire [63:0] _GEN_8748 = uncached ? {{32'd0}, saved_1_inst} : _GEN_7197; // @[ICache.scala 169:30 91:22]
  wire  _GEN_8749 = uncached ? saved_0_valid : _GEN_7198; // @[ICache.scala 169:30 91:22]
  wire  _GEN_8750 = uncached ? saved_1_valid : _GEN_7199; // @[ICache.scala 169:30 91:22]
  wire [19:0] _GEN_8762 = ~translation_ok ? {{3'd0}, tag_ram_wdata} : _GEN_7210; // @[ICache.scala 166:31 68:30]
  wire [63:0] _GEN_10300 = ~translation_ok ? {{32'd0}, saved_1_inst} : _GEN_8748; // @[ICache.scala 166:31 91:22]
  wire [19:0] _GEN_10314 = io_cpu_req ? _GEN_8762 : {{3'd0}, tag_ram_wdata}; // @[ICache.scala 165:24 68:30]
  wire [63:0] _GEN_11852 = io_cpu_req ? _GEN_10300 : {{32'd0}, saved_1_inst}; // @[ICache.scala 165:24 91:22]
  wire  _T_16 = ~inst_vpn[12]; // @[ICache.scala 201:71]
  wire  _T_17 = _T_16 & io_cpu_tlb2_entry_V0; // @[ICache.scala 203:11]
  wire  _T_19 = io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_V1 | _T_17); // @[ICache.scala 201:27]
  wire [19:0] _tlb_ppn_T_1 = inst_vpn[12] ? io_cpu_tlb2_entry_PFN1 : io_cpu_tlb2_entry_PFN0; // @[ICache.scala 207:28]
  wire  _tlb_uncached_T_1 = inst_vpn[12] ? io_cpu_tlb2_entry_C1 : io_cpu_tlb2_entry_C0; // @[ICache.scala 208:28]
  wire [18:0] _GEN_11856 = _T_19 ? io_cpu_tlb2_vpn : {{2'd0}, tlb_vpn}; // @[ICache.scala 204:9 206:22 40:20]
  wire [19:0] _GEN_11857 = _T_19 ? _tlb_ppn_T_1 : {{3'd0}, tlb_ppn}; // @[ICache.scala 204:9 207:22 40:20]
  wire  _GEN_11859 = _T_19 | _GEN_1028; // @[ICache.scala 204:9 209:22]
  wire  _GEN_11863 = io_axi_ar_ready ? 1'h0 : arvalid; // @[ICache.scala 219:31 220:19 142:24]
  wire  _GEN_11864 = io_axi_ar_ready | rready; // @[ICache.scala 219:31 221:19 147:23]
  wire  _T_21 = io_axi_r_ready & io_axi_r_valid; // @[Decoupled.scala 52:35]
  wire [2:0] _GEN_11865 = _T_21 ? 3'h4 : state; // @[ICache.scala 223:33 224:24 48:81]
  wire [31:0] _GEN_11866 = _T_21 ? io_axi_r_bits_data : saved_0_inst; // @[ICache.scala 223:33 225:24 91:22]
  wire  _GEN_11867 = _T_21 | saved_0_valid; // @[ICache.scala 223:33 226:24 91:22]
  wire  _GEN_11868 = _T_21 ? 1'h0 : rready; // @[ICache.scala 147:23 223:33 227:24]
  wire  _GEN_11869 = io_axi_ar_valid ? _GEN_11863 : arvalid; // @[ICache.scala 142:24 218:29]
  wire  _GEN_11870 = io_axi_ar_valid ? _GEN_11864 : _GEN_11868; // @[ICache.scala 218:29]
  wire [2:0] _GEN_11871 = io_axi_ar_valid ? state : _GEN_11865; // @[ICache.scala 218:29 48:81]
  wire [31:0] _GEN_11872 = io_axi_ar_valid ? saved_0_inst : _GEN_11866; // @[ICache.scala 218:29 91:22]
  wire  _GEN_11873 = io_axi_ar_valid ? saved_0_valid : _GEN_11867; // @[ICache.scala 218:29 91:22]
  wire [4:0] _axi_cnt_T_1 = axi_cnt + 5'h1; // @[ICache.scala 239:57]
  wire [7:0] _GEN_11875 = _GEN_3588 ? data_wen_1 : data_wen_0; // @[ICache.scala 240:{49,49}]
  wire [7:0] _data_wen_T = ~_GEN_11875; // @[ICache.scala 240:49]
  wire [7:0] _GEN_11876 = ~_GEN_3588 ? _data_wen_T : data_wen_0; // @[ICache.scala 240:{46,46} 66:30]
  wire [7:0] _GEN_11877 = _GEN_3588 ? _data_wen_T : data_wen_1; // @[ICache.scala 240:{46,46} 66:30]
  wire [7:0] _GEN_11878 = ~_GEN_3588 ? 8'h0 : data_wen_0; // @[ICache.scala 243:{46,46} 66:30]
  wire [7:0] _GEN_11879 = _GEN_3588 ? 8'h0 : data_wen_1; // @[ICache.scala 243:{46,46} 66:30]
  wire  _GEN_11880 = ~_GEN_3588 ? 1'h0 : tag_wen_0; // @[ICache.scala 244:{46,46} 67:30]
  wire  _GEN_11881 = _GEN_3588 ? 1'h0 : tag_wen_1; // @[ICache.scala 244:{46,46} 67:30]
  wire [4:0] _GEN_11882 = ~io_axi_r_bits_last ? _axi_cnt_T_1 : axi_cnt; // @[ICache.scala 109:24 238:37 239:46]
  wire [7:0] _GEN_11883 = ~io_axi_r_bits_last ? _GEN_11876 : _GEN_11878; // @[ICache.scala 238:37]
  wire [7:0] _GEN_11884 = ~io_axi_r_bits_last ? _GEN_11877 : _GEN_11879; // @[ICache.scala 238:37]
  wire  _GEN_11885 = ~io_axi_r_bits_last & rready; // @[ICache.scala 147:23 238:37 242:46]
  wire  _GEN_11886 = ~io_axi_r_bits_last ? tag_wen_0 : _GEN_11880; // @[ICache.scala 238:37 67:30]
  wire  _GEN_11887 = ~io_axi_r_bits_last ? tag_wen_1 : _GEN_11881; // @[ICache.scala 238:37 67:30]
  wire [2:0] _GEN_11888 = ~io_axi_r_ready ? 3'h0 : state; // @[ICache.scala 246:37 247:17 48:81]
  wire [4:0] _GEN_11889 = _T_21 ? _GEN_11882 : axi_cnt; // @[ICache.scala 109:24 237:29]
  wire [7:0] _GEN_11890 = _T_21 ? _GEN_11883 : data_wen_0; // @[ICache.scala 237:29 66:30]
  wire [7:0] _GEN_11891 = _T_21 ? _GEN_11884 : data_wen_1; // @[ICache.scala 237:29 66:30]
  wire  _GEN_11892 = _T_21 ? _GEN_11885 : rready; // @[ICache.scala 147:23 237:29]
  wire  _GEN_11893 = _T_21 ? _GEN_11886 : tag_wen_0; // @[ICache.scala 237:29 67:30]
  wire  _GEN_11894 = _T_21 ? _GEN_11887 : tag_wen_1; // @[ICache.scala 237:29 67:30]
  wire [2:0] _GEN_11895 = _T_21 ? state : _GEN_11888; // @[ICache.scala 237:29 48:81]
  wire  _GEN_11896 = io_axi_ar_valid ? _GEN_11864 : _GEN_11892; // @[ICache.scala 231:29]
  wire [4:0] _GEN_11897 = io_axi_ar_valid ? axi_cnt : _GEN_11889; // @[ICache.scala 109:24 231:29]
  wire [7:0] _GEN_11898 = io_axi_ar_valid ? data_wen_0 : _GEN_11890; // @[ICache.scala 231:29 66:30]
  wire [7:0] _GEN_11899 = io_axi_ar_valid ? data_wen_1 : _GEN_11891; // @[ICache.scala 231:29 66:30]
  wire  _GEN_11900 = io_axi_ar_valid ? tag_wen_0 : _GEN_11893; // @[ICache.scala 231:29 67:30]
  wire  _GEN_11901 = io_axi_ar_valid ? tag_wen_1 : _GEN_11894; // @[ICache.scala 231:29 67:30]
  wire [2:0] _GEN_11902 = io_axi_ar_valid ? state : _GEN_11895; // @[ICache.scala 231:29 48:81]
  wire [2:0] _GEN_11903 = _T_2 & _T ? 3'h0 : state; // @[ICache.scala 252:55 253:24 48:81]
  wire  _GEN_11904 = _T_2 & _T ? 1'h0 : tlb1_invalid; // @[ICache.scala 151:21 252:55 254:24]
  wire  _GEN_11906 = _T_2 & _T ? 1'h0 : saved_0_valid; // @[ICache.scala 252:55 256:24 91:22]
  wire  _GEN_11907 = _T_2 & _T ? 1'h0 : saved_1_valid; // @[ICache.scala 252:55 257:24 91:22]
  wire [2:0] _GEN_11908 = 3'h4 == state ? _GEN_11903 : state; // @[ICache.scala 163:17 48:81]
  wire  _GEN_11909 = 3'h4 == state ? _GEN_11904 : tlb1_invalid; // @[ICache.scala 163:17 151:21]
  wire  _GEN_11911 = 3'h4 == state ? _GEN_11906 : saved_0_valid; // @[ICache.scala 163:17 91:22]
  wire  _GEN_11912 = 3'h4 == state ? _GEN_11907 : saved_1_valid; // @[ICache.scala 163:17 91:22]
  wire  _GEN_11913 = 3'h3 == state ? _GEN_11869 : arvalid; // @[ICache.scala 163:17 142:24]
  wire  _GEN_11914 = 3'h3 == state ? _GEN_11896 : rready; // @[ICache.scala 163:17 147:23]
  wire [4:0] _GEN_11915 = 3'h3 == state ? _GEN_11897 : axi_cnt; // @[ICache.scala 163:17 109:24]
  wire [7:0] _GEN_11916 = 3'h3 == state ? _GEN_11898 : data_wen_0; // @[ICache.scala 163:17 66:30]
  wire [7:0] _GEN_11917 = 3'h3 == state ? _GEN_11899 : data_wen_1; // @[ICache.scala 163:17 66:30]
  wire  _GEN_11918 = 3'h3 == state ? _GEN_11900 : tag_wen_0; // @[ICache.scala 163:17 67:30]
  wire  _GEN_11919 = 3'h3 == state ? _GEN_11901 : tag_wen_1; // @[ICache.scala 163:17 67:30]
  wire [2:0] _GEN_11920 = 3'h3 == state ? _GEN_11902 : _GEN_11908; // @[ICache.scala 163:17]
  wire  _GEN_11921 = 3'h3 == state ? tlb1_invalid : _GEN_11909; // @[ICache.scala 163:17 151:21]
  wire  _GEN_11923 = 3'h3 == state ? saved_0_valid : _GEN_11911; // @[ICache.scala 163:17 91:22]
  wire  _GEN_11924 = 3'h3 == state ? saved_1_valid : _GEN_11912; // @[ICache.scala 163:17 91:22]
  wire [18:0] _GEN_11939 = 3'h1 == state ? _GEN_11856 : {{2'd0}, tlb_vpn}; // @[ICache.scala 163:17 40:20]
  wire [19:0] _GEN_11940 = 3'h1 == state ? _GEN_11857 : {{3'd0}, tlb_ppn}; // @[ICache.scala 163:17 40:20]
  wire [19:0] _GEN_11966 = 3'h0 == state ? _GEN_10314 : {{3'd0}, tag_ram_wdata}; // @[ICache.scala 163:17 68:30]
  wire [63:0] _GEN_13504 = 3'h0 == state ? _GEN_11852 : {{32'd0}, saved_1_inst}; // @[ICache.scala 163:17 91:22]
  wire [18:0] _GEN_13507 = 3'h0 == state ? {{2'd0}, tlb_vpn} : _GEN_11939; // @[ICache.scala 163:17 40:20]
  wire [19:0] _GEN_13508 = 3'h0 == state ? {{3'd0}, tlb_ppn} : _GEN_11940; // @[ICache.scala 163:17 40:20]
  wire [18:0] _GEN_19663 = reset ? 19'h0 : _GEN_13507; // @[ICache.scala 40:{20,20}]
  wire [19:0] _GEN_19664 = reset ? 20'h0 : _GEN_13508; // @[ICache.scala 40:{20,20}]
  wire [19:0] _GEN_19665 = reset ? 20'h0 : _GEN_11966; // @[ICache.scala 68:{30,30}]
  wire [63:0] _GEN_19666 = reset ? 64'h0 : _GEN_13504; // @[ICache.scala 91:{22,22}]
  Bank bank_ram ( // @[ICache.scala 112:24]
    .clock(bank_ram_clock),
    .reset(bank_ram_reset),
    .io_way_0_r_addr(bank_ram_io_way_0_r_addr),
    .io_way_0_r_data(bank_ram_io_way_0_r_data),
    .io_way_0_w_addr(bank_ram_io_way_0_w_addr),
    .io_way_0_w_en(bank_ram_io_way_0_w_en),
    .io_way_0_w_data(bank_ram_io_way_0_w_data),
    .io_way_1_r_addr(bank_ram_io_way_1_r_addr),
    .io_way_1_r_data(bank_ram_io_way_1_r_data),
    .io_way_1_w_addr(bank_ram_io_way_1_w_addr),
    .io_way_1_w_en(bank_ram_io_way_1_w_en),
    .io_way_1_w_data(bank_ram_io_way_1_w_data)
  );
  Tag tag_ram ( // @[ICache.scala 125:23]
    .clock(tag_ram_clock),
    .reset(tag_ram_reset),
    .io_way_0_r_addr(tag_ram_io_way_0_r_addr),
    .io_way_0_r_data(tag_ram_io_way_0_r_data),
    .io_way_0_w_addr(tag_ram_io_way_0_w_addr),
    .io_way_0_w_en(tag_ram_io_way_0_w_en),
    .io_way_0_w_data(tag_ram_io_way_0_w_data),
    .io_way_1_r_addr(tag_ram_io_way_1_r_addr),
    .io_way_1_r_data(tag_ram_io_way_1_r_data),
    .io_way_1_w_addr(tag_ram_io_way_1_w_addr),
    .io_way_1_w_en(tag_ram_io_way_1_w_en),
    .io_way_1_w_data(tag_ram_io_way_1_w_data)
  );
  assign io_cpu_inst_0 = _io_cpu_icache_stall_T ? cache_inst_0 : saved_0_inst; // @[ICache.scala 106:30]
  assign io_cpu_inst_1 = _io_cpu_icache_stall_T ? _GEN_3[63:32] : saved_1_inst; // @[ICache.scala 107:30]
  assign io_cpu_inst_valid_0 = _io_cpu_inst_valid_0_T_1 & io_cpu_req; // @[ICache.scala 104:83]
  assign io_cpu_inst_valid_1 = _io_cpu_inst_valid_1_T_1 & io_cpu_req; // @[ICache.scala 105:83]
  assign io_cpu_icache_stall = _io_cpu_icache_stall_T ? _io_cpu_icache_stall_T_2 : _bram_addr_choose_next_T_1; // @[ICache.scala 98:29]
  assign io_cpu_tlb1_refill = 1'h0; // @[ICache.scala 155:8]
  assign io_cpu_tlb1_invalid = tlb1_invalid; // @[ICache.scala 155:8]
  assign io_cpu_tlb2_vpn = 19'h0; // @[ICache.scala 162:19]
  assign io_axi_ar_valid = arvalid; // @[ICache.scala 144:11]
  assign io_axi_ar_bits_addr = ar_addr; // @[ICache.scala 143:6]
  assign io_axi_ar_bits_len = ar_len; // @[ICache.scala 143:6]
  assign io_axi_ar_bits_size = ar_size; // @[ICache.scala 143:6]
  assign io_axi_r_ready = rready; // @[ICache.scala 149:10]
  assign bank_ram_clock = clock;
  assign bank_ram_reset = reset;
  assign bank_ram_io_way_0_r_addr = _GEN_1[11:3]; // @[ICache.scala 61:58]
  assign bank_ram_io_way_0_w_addr = {replace_line_addr,axi_cnt[3:1]}; // @[Cat.scala 33:92]
  assign bank_ram_io_way_0_w_en = data_wen_0; // @[ICache.scala 115:31]
  assign bank_ram_io_way_0_w_data = axi_cnt[0] ? _bank_ram_io_way_0_w_data_T_1 : _bank_ram_io_way_0_w_data_T_2; // @[ICache.scala 117:37]
  assign bank_ram_io_way_1_r_addr = _GEN_1[11:3]; // @[ICache.scala 61:58]
  assign bank_ram_io_way_1_w_addr = {replace_line_addr,axi_cnt[3:1]}; // @[Cat.scala 33:92]
  assign bank_ram_io_way_1_w_en = data_wen_1; // @[ICache.scala 115:31]
  assign bank_ram_io_way_1_w_data = axi_cnt[0] ? _bank_ram_io_way_0_w_data_T_1 : _bank_ram_io_way_0_w_data_T_2; // @[ICache.scala 117:37]
  assign tag_ram_clock = clock;
  assign tag_ram_reset = reset;
  assign tag_ram_io_way_0_r_addr = {{3'd0}, bram_line_addr}; // @[ICache.scala 127:30]
  assign tag_ram_io_way_0_w_addr = {{3'd0}, replace_line_addr}; // @[ICache.scala 129:30]
  assign tag_ram_io_way_0_w_en = tag_wen_0; // @[ICache.scala 128:30]
  assign tag_ram_io_way_0_w_data = tag_ram_wdata; // @[ICache.scala 130:30]
  assign tag_ram_io_way_1_r_addr = {{3'd0}, bram_line_addr}; // @[ICache.scala 127:30]
  assign tag_ram_io_way_1_w_addr = {{3'd0}, replace_line_addr}; // @[ICache.scala 129:30]
  assign tag_ram_io_way_1_w_en = tag_wen_1; // @[ICache.scala 128:30]
  assign tag_ram_io_way_1_w_data = tag_ram_wdata; // @[ICache.scala 130:30]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 34:21]
      meta_0_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_0_valid_0 <= _GEN_2053;
        end else begin
          meta_0_valid_0 <= _GEN_7211;
        end
      end else begin
        meta_0_valid_0 <= _GEN_2053;
      end
    end else begin
      meta_0_valid_0 <= _GEN_2053;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_0_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_0_valid_1 <= _GEN_2565;
        end else begin
          meta_0_valid_1 <= _GEN_7212;
        end
      end else begin
        meta_0_valid_1 <= _GEN_2565;
      end
    end else begin
      meta_0_valid_1 <= _GEN_2565;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_0_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_0_lru <= _GEN_8236;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_1_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_1_valid_0 <= _GEN_2054;
        end else begin
          meta_1_valid_0 <= _GEN_7213;
        end
      end else begin
        meta_1_valid_0 <= _GEN_2054;
      end
    end else begin
      meta_1_valid_0 <= _GEN_2054;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_1_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_1_valid_1 <= _GEN_2566;
        end else begin
          meta_1_valid_1 <= _GEN_7214;
        end
      end else begin
        meta_1_valid_1 <= _GEN_2566;
      end
    end else begin
      meta_1_valid_1 <= _GEN_2566;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_1_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_1_lru <= _GEN_8237;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_2_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_2_valid_0 <= _GEN_2055;
        end else begin
          meta_2_valid_0 <= _GEN_7215;
        end
      end else begin
        meta_2_valid_0 <= _GEN_2055;
      end
    end else begin
      meta_2_valid_0 <= _GEN_2055;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_2_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_2_valid_1 <= _GEN_2567;
        end else begin
          meta_2_valid_1 <= _GEN_7216;
        end
      end else begin
        meta_2_valid_1 <= _GEN_2567;
      end
    end else begin
      meta_2_valid_1 <= _GEN_2567;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_2_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_2_lru <= _GEN_8238;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_3_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_3_valid_0 <= _GEN_2056;
        end else begin
          meta_3_valid_0 <= _GEN_7217;
        end
      end else begin
        meta_3_valid_0 <= _GEN_2056;
      end
    end else begin
      meta_3_valid_0 <= _GEN_2056;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_3_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_3_valid_1 <= _GEN_2568;
        end else begin
          meta_3_valid_1 <= _GEN_7218;
        end
      end else begin
        meta_3_valid_1 <= _GEN_2568;
      end
    end else begin
      meta_3_valid_1 <= _GEN_2568;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_3_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_3_lru <= _GEN_8239;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_4_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_4_valid_0 <= _GEN_2057;
        end else begin
          meta_4_valid_0 <= _GEN_7219;
        end
      end else begin
        meta_4_valid_0 <= _GEN_2057;
      end
    end else begin
      meta_4_valid_0 <= _GEN_2057;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_4_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_4_valid_1 <= _GEN_2569;
        end else begin
          meta_4_valid_1 <= _GEN_7220;
        end
      end else begin
        meta_4_valid_1 <= _GEN_2569;
      end
    end else begin
      meta_4_valid_1 <= _GEN_2569;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_4_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_4_lru <= _GEN_8240;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_5_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_5_valid_0 <= _GEN_2058;
        end else begin
          meta_5_valid_0 <= _GEN_7221;
        end
      end else begin
        meta_5_valid_0 <= _GEN_2058;
      end
    end else begin
      meta_5_valid_0 <= _GEN_2058;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_5_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_5_valid_1 <= _GEN_2570;
        end else begin
          meta_5_valid_1 <= _GEN_7222;
        end
      end else begin
        meta_5_valid_1 <= _GEN_2570;
      end
    end else begin
      meta_5_valid_1 <= _GEN_2570;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_5_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_5_lru <= _GEN_8241;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_6_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_6_valid_0 <= _GEN_2059;
        end else begin
          meta_6_valid_0 <= _GEN_7223;
        end
      end else begin
        meta_6_valid_0 <= _GEN_2059;
      end
    end else begin
      meta_6_valid_0 <= _GEN_2059;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_6_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_6_valid_1 <= _GEN_2571;
        end else begin
          meta_6_valid_1 <= _GEN_7224;
        end
      end else begin
        meta_6_valid_1 <= _GEN_2571;
      end
    end else begin
      meta_6_valid_1 <= _GEN_2571;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_6_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_6_lru <= _GEN_8242;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_7_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_7_valid_0 <= _GEN_2060;
        end else begin
          meta_7_valid_0 <= _GEN_7225;
        end
      end else begin
        meta_7_valid_0 <= _GEN_2060;
      end
    end else begin
      meta_7_valid_0 <= _GEN_2060;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_7_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_7_valid_1 <= _GEN_2572;
        end else begin
          meta_7_valid_1 <= _GEN_7226;
        end
      end else begin
        meta_7_valid_1 <= _GEN_2572;
      end
    end else begin
      meta_7_valid_1 <= _GEN_2572;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_7_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_7_lru <= _GEN_8243;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_8_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_8_valid_0 <= _GEN_2061;
        end else begin
          meta_8_valid_0 <= _GEN_7227;
        end
      end else begin
        meta_8_valid_0 <= _GEN_2061;
      end
    end else begin
      meta_8_valid_0 <= _GEN_2061;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_8_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_8_valid_1 <= _GEN_2573;
        end else begin
          meta_8_valid_1 <= _GEN_7228;
        end
      end else begin
        meta_8_valid_1 <= _GEN_2573;
      end
    end else begin
      meta_8_valid_1 <= _GEN_2573;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_8_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_8_lru <= _GEN_8244;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_9_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_9_valid_0 <= _GEN_2062;
        end else begin
          meta_9_valid_0 <= _GEN_7229;
        end
      end else begin
        meta_9_valid_0 <= _GEN_2062;
      end
    end else begin
      meta_9_valid_0 <= _GEN_2062;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_9_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_9_valid_1 <= _GEN_2574;
        end else begin
          meta_9_valid_1 <= _GEN_7230;
        end
      end else begin
        meta_9_valid_1 <= _GEN_2574;
      end
    end else begin
      meta_9_valid_1 <= _GEN_2574;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_9_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_9_lru <= _GEN_8245;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_10_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_10_valid_0 <= _GEN_2063;
        end else begin
          meta_10_valid_0 <= _GEN_7231;
        end
      end else begin
        meta_10_valid_0 <= _GEN_2063;
      end
    end else begin
      meta_10_valid_0 <= _GEN_2063;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_10_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_10_valid_1 <= _GEN_2575;
        end else begin
          meta_10_valid_1 <= _GEN_7232;
        end
      end else begin
        meta_10_valid_1 <= _GEN_2575;
      end
    end else begin
      meta_10_valid_1 <= _GEN_2575;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_10_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_10_lru <= _GEN_8246;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_11_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_11_valid_0 <= _GEN_2064;
        end else begin
          meta_11_valid_0 <= _GEN_7233;
        end
      end else begin
        meta_11_valid_0 <= _GEN_2064;
      end
    end else begin
      meta_11_valid_0 <= _GEN_2064;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_11_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_11_valid_1 <= _GEN_2576;
        end else begin
          meta_11_valid_1 <= _GEN_7234;
        end
      end else begin
        meta_11_valid_1 <= _GEN_2576;
      end
    end else begin
      meta_11_valid_1 <= _GEN_2576;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_11_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_11_lru <= _GEN_8247;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_12_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_12_valid_0 <= _GEN_2065;
        end else begin
          meta_12_valid_0 <= _GEN_7235;
        end
      end else begin
        meta_12_valid_0 <= _GEN_2065;
      end
    end else begin
      meta_12_valid_0 <= _GEN_2065;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_12_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_12_valid_1 <= _GEN_2577;
        end else begin
          meta_12_valid_1 <= _GEN_7236;
        end
      end else begin
        meta_12_valid_1 <= _GEN_2577;
      end
    end else begin
      meta_12_valid_1 <= _GEN_2577;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_12_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_12_lru <= _GEN_8248;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_13_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_13_valid_0 <= _GEN_2066;
        end else begin
          meta_13_valid_0 <= _GEN_7237;
        end
      end else begin
        meta_13_valid_0 <= _GEN_2066;
      end
    end else begin
      meta_13_valid_0 <= _GEN_2066;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_13_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_13_valid_1 <= _GEN_2578;
        end else begin
          meta_13_valid_1 <= _GEN_7238;
        end
      end else begin
        meta_13_valid_1 <= _GEN_2578;
      end
    end else begin
      meta_13_valid_1 <= _GEN_2578;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_13_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_13_lru <= _GEN_8249;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_14_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_14_valid_0 <= _GEN_2067;
        end else begin
          meta_14_valid_0 <= _GEN_7239;
        end
      end else begin
        meta_14_valid_0 <= _GEN_2067;
      end
    end else begin
      meta_14_valid_0 <= _GEN_2067;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_14_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_14_valid_1 <= _GEN_2579;
        end else begin
          meta_14_valid_1 <= _GEN_7240;
        end
      end else begin
        meta_14_valid_1 <= _GEN_2579;
      end
    end else begin
      meta_14_valid_1 <= _GEN_2579;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_14_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_14_lru <= _GEN_8250;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_15_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_15_valid_0 <= _GEN_2068;
        end else begin
          meta_15_valid_0 <= _GEN_7241;
        end
      end else begin
        meta_15_valid_0 <= _GEN_2068;
      end
    end else begin
      meta_15_valid_0 <= _GEN_2068;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_15_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_15_valid_1 <= _GEN_2580;
        end else begin
          meta_15_valid_1 <= _GEN_7242;
        end
      end else begin
        meta_15_valid_1 <= _GEN_2580;
      end
    end else begin
      meta_15_valid_1 <= _GEN_2580;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_15_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_15_lru <= _GEN_8251;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_16_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_16_valid_0 <= _GEN_2069;
        end else begin
          meta_16_valid_0 <= _GEN_7243;
        end
      end else begin
        meta_16_valid_0 <= _GEN_2069;
      end
    end else begin
      meta_16_valid_0 <= _GEN_2069;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_16_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_16_valid_1 <= _GEN_2581;
        end else begin
          meta_16_valid_1 <= _GEN_7244;
        end
      end else begin
        meta_16_valid_1 <= _GEN_2581;
      end
    end else begin
      meta_16_valid_1 <= _GEN_2581;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_16_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_16_lru <= _GEN_8252;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_17_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_17_valid_0 <= _GEN_2070;
        end else begin
          meta_17_valid_0 <= _GEN_7245;
        end
      end else begin
        meta_17_valid_0 <= _GEN_2070;
      end
    end else begin
      meta_17_valid_0 <= _GEN_2070;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_17_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_17_valid_1 <= _GEN_2582;
        end else begin
          meta_17_valid_1 <= _GEN_7246;
        end
      end else begin
        meta_17_valid_1 <= _GEN_2582;
      end
    end else begin
      meta_17_valid_1 <= _GEN_2582;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_17_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_17_lru <= _GEN_8253;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_18_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_18_valid_0 <= _GEN_2071;
        end else begin
          meta_18_valid_0 <= _GEN_7247;
        end
      end else begin
        meta_18_valid_0 <= _GEN_2071;
      end
    end else begin
      meta_18_valid_0 <= _GEN_2071;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_18_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_18_valid_1 <= _GEN_2583;
        end else begin
          meta_18_valid_1 <= _GEN_7248;
        end
      end else begin
        meta_18_valid_1 <= _GEN_2583;
      end
    end else begin
      meta_18_valid_1 <= _GEN_2583;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_18_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_18_lru <= _GEN_8254;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_19_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_19_valid_0 <= _GEN_2072;
        end else begin
          meta_19_valid_0 <= _GEN_7249;
        end
      end else begin
        meta_19_valid_0 <= _GEN_2072;
      end
    end else begin
      meta_19_valid_0 <= _GEN_2072;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_19_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_19_valid_1 <= _GEN_2584;
        end else begin
          meta_19_valid_1 <= _GEN_7250;
        end
      end else begin
        meta_19_valid_1 <= _GEN_2584;
      end
    end else begin
      meta_19_valid_1 <= _GEN_2584;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_19_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_19_lru <= _GEN_8255;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_20_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_20_valid_0 <= _GEN_2073;
        end else begin
          meta_20_valid_0 <= _GEN_7251;
        end
      end else begin
        meta_20_valid_0 <= _GEN_2073;
      end
    end else begin
      meta_20_valid_0 <= _GEN_2073;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_20_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_20_valid_1 <= _GEN_2585;
        end else begin
          meta_20_valid_1 <= _GEN_7252;
        end
      end else begin
        meta_20_valid_1 <= _GEN_2585;
      end
    end else begin
      meta_20_valid_1 <= _GEN_2585;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_20_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_20_lru <= _GEN_8256;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_21_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_21_valid_0 <= _GEN_2074;
        end else begin
          meta_21_valid_0 <= _GEN_7253;
        end
      end else begin
        meta_21_valid_0 <= _GEN_2074;
      end
    end else begin
      meta_21_valid_0 <= _GEN_2074;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_21_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_21_valid_1 <= _GEN_2586;
        end else begin
          meta_21_valid_1 <= _GEN_7254;
        end
      end else begin
        meta_21_valid_1 <= _GEN_2586;
      end
    end else begin
      meta_21_valid_1 <= _GEN_2586;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_21_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_21_lru <= _GEN_8257;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_22_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_22_valid_0 <= _GEN_2075;
        end else begin
          meta_22_valid_0 <= _GEN_7255;
        end
      end else begin
        meta_22_valid_0 <= _GEN_2075;
      end
    end else begin
      meta_22_valid_0 <= _GEN_2075;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_22_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_22_valid_1 <= _GEN_2587;
        end else begin
          meta_22_valid_1 <= _GEN_7256;
        end
      end else begin
        meta_22_valid_1 <= _GEN_2587;
      end
    end else begin
      meta_22_valid_1 <= _GEN_2587;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_22_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_22_lru <= _GEN_8258;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_23_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_23_valid_0 <= _GEN_2076;
        end else begin
          meta_23_valid_0 <= _GEN_7257;
        end
      end else begin
        meta_23_valid_0 <= _GEN_2076;
      end
    end else begin
      meta_23_valid_0 <= _GEN_2076;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_23_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_23_valid_1 <= _GEN_2588;
        end else begin
          meta_23_valid_1 <= _GEN_7258;
        end
      end else begin
        meta_23_valid_1 <= _GEN_2588;
      end
    end else begin
      meta_23_valid_1 <= _GEN_2588;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_23_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_23_lru <= _GEN_8259;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_24_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_24_valid_0 <= _GEN_2077;
        end else begin
          meta_24_valid_0 <= _GEN_7259;
        end
      end else begin
        meta_24_valid_0 <= _GEN_2077;
      end
    end else begin
      meta_24_valid_0 <= _GEN_2077;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_24_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_24_valid_1 <= _GEN_2589;
        end else begin
          meta_24_valid_1 <= _GEN_7260;
        end
      end else begin
        meta_24_valid_1 <= _GEN_2589;
      end
    end else begin
      meta_24_valid_1 <= _GEN_2589;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_24_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_24_lru <= _GEN_8260;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_25_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_25_valid_0 <= _GEN_2078;
        end else begin
          meta_25_valid_0 <= _GEN_7261;
        end
      end else begin
        meta_25_valid_0 <= _GEN_2078;
      end
    end else begin
      meta_25_valid_0 <= _GEN_2078;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_25_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_25_valid_1 <= _GEN_2590;
        end else begin
          meta_25_valid_1 <= _GEN_7262;
        end
      end else begin
        meta_25_valid_1 <= _GEN_2590;
      end
    end else begin
      meta_25_valid_1 <= _GEN_2590;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_25_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_25_lru <= _GEN_8261;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_26_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_26_valid_0 <= _GEN_2079;
        end else begin
          meta_26_valid_0 <= _GEN_7263;
        end
      end else begin
        meta_26_valid_0 <= _GEN_2079;
      end
    end else begin
      meta_26_valid_0 <= _GEN_2079;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_26_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_26_valid_1 <= _GEN_2591;
        end else begin
          meta_26_valid_1 <= _GEN_7264;
        end
      end else begin
        meta_26_valid_1 <= _GEN_2591;
      end
    end else begin
      meta_26_valid_1 <= _GEN_2591;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_26_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_26_lru <= _GEN_8262;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_27_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_27_valid_0 <= _GEN_2080;
        end else begin
          meta_27_valid_0 <= _GEN_7265;
        end
      end else begin
        meta_27_valid_0 <= _GEN_2080;
      end
    end else begin
      meta_27_valid_0 <= _GEN_2080;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_27_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_27_valid_1 <= _GEN_2592;
        end else begin
          meta_27_valid_1 <= _GEN_7266;
        end
      end else begin
        meta_27_valid_1 <= _GEN_2592;
      end
    end else begin
      meta_27_valid_1 <= _GEN_2592;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_27_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_27_lru <= _GEN_8263;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_28_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_28_valid_0 <= _GEN_2081;
        end else begin
          meta_28_valid_0 <= _GEN_7267;
        end
      end else begin
        meta_28_valid_0 <= _GEN_2081;
      end
    end else begin
      meta_28_valid_0 <= _GEN_2081;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_28_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_28_valid_1 <= _GEN_2593;
        end else begin
          meta_28_valid_1 <= _GEN_7268;
        end
      end else begin
        meta_28_valid_1 <= _GEN_2593;
      end
    end else begin
      meta_28_valid_1 <= _GEN_2593;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_28_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_28_lru <= _GEN_8264;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_29_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_29_valid_0 <= _GEN_2082;
        end else begin
          meta_29_valid_0 <= _GEN_7269;
        end
      end else begin
        meta_29_valid_0 <= _GEN_2082;
      end
    end else begin
      meta_29_valid_0 <= _GEN_2082;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_29_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_29_valid_1 <= _GEN_2594;
        end else begin
          meta_29_valid_1 <= _GEN_7270;
        end
      end else begin
        meta_29_valid_1 <= _GEN_2594;
      end
    end else begin
      meta_29_valid_1 <= _GEN_2594;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_29_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_29_lru <= _GEN_8265;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_30_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_30_valid_0 <= _GEN_2083;
        end else begin
          meta_30_valid_0 <= _GEN_7271;
        end
      end else begin
        meta_30_valid_0 <= _GEN_2083;
      end
    end else begin
      meta_30_valid_0 <= _GEN_2083;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_30_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_30_valid_1 <= _GEN_2595;
        end else begin
          meta_30_valid_1 <= _GEN_7272;
        end
      end else begin
        meta_30_valid_1 <= _GEN_2595;
      end
    end else begin
      meta_30_valid_1 <= _GEN_2595;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_30_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_30_lru <= _GEN_8266;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_31_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_31_valid_0 <= _GEN_2084;
        end else begin
          meta_31_valid_0 <= _GEN_7273;
        end
      end else begin
        meta_31_valid_0 <= _GEN_2084;
      end
    end else begin
      meta_31_valid_0 <= _GEN_2084;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_31_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_31_valid_1 <= _GEN_2596;
        end else begin
          meta_31_valid_1 <= _GEN_7274;
        end
      end else begin
        meta_31_valid_1 <= _GEN_2596;
      end
    end else begin
      meta_31_valid_1 <= _GEN_2596;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_31_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_31_lru <= _GEN_8267;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_32_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_32_valid_0 <= _GEN_2085;
        end else begin
          meta_32_valid_0 <= _GEN_7275;
        end
      end else begin
        meta_32_valid_0 <= _GEN_2085;
      end
    end else begin
      meta_32_valid_0 <= _GEN_2085;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_32_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_32_valid_1 <= _GEN_2597;
        end else begin
          meta_32_valid_1 <= _GEN_7276;
        end
      end else begin
        meta_32_valid_1 <= _GEN_2597;
      end
    end else begin
      meta_32_valid_1 <= _GEN_2597;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_32_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_32_lru <= _GEN_8268;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_33_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_33_valid_0 <= _GEN_2086;
        end else begin
          meta_33_valid_0 <= _GEN_7277;
        end
      end else begin
        meta_33_valid_0 <= _GEN_2086;
      end
    end else begin
      meta_33_valid_0 <= _GEN_2086;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_33_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_33_valid_1 <= _GEN_2598;
        end else begin
          meta_33_valid_1 <= _GEN_7278;
        end
      end else begin
        meta_33_valid_1 <= _GEN_2598;
      end
    end else begin
      meta_33_valid_1 <= _GEN_2598;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_33_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_33_lru <= _GEN_8269;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_34_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_34_valid_0 <= _GEN_2087;
        end else begin
          meta_34_valid_0 <= _GEN_7279;
        end
      end else begin
        meta_34_valid_0 <= _GEN_2087;
      end
    end else begin
      meta_34_valid_0 <= _GEN_2087;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_34_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_34_valid_1 <= _GEN_2599;
        end else begin
          meta_34_valid_1 <= _GEN_7280;
        end
      end else begin
        meta_34_valid_1 <= _GEN_2599;
      end
    end else begin
      meta_34_valid_1 <= _GEN_2599;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_34_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_34_lru <= _GEN_8270;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_35_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_35_valid_0 <= _GEN_2088;
        end else begin
          meta_35_valid_0 <= _GEN_7281;
        end
      end else begin
        meta_35_valid_0 <= _GEN_2088;
      end
    end else begin
      meta_35_valid_0 <= _GEN_2088;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_35_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_35_valid_1 <= _GEN_2600;
        end else begin
          meta_35_valid_1 <= _GEN_7282;
        end
      end else begin
        meta_35_valid_1 <= _GEN_2600;
      end
    end else begin
      meta_35_valid_1 <= _GEN_2600;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_35_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_35_lru <= _GEN_8271;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_36_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_36_valid_0 <= _GEN_2089;
        end else begin
          meta_36_valid_0 <= _GEN_7283;
        end
      end else begin
        meta_36_valid_0 <= _GEN_2089;
      end
    end else begin
      meta_36_valid_0 <= _GEN_2089;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_36_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_36_valid_1 <= _GEN_2601;
        end else begin
          meta_36_valid_1 <= _GEN_7284;
        end
      end else begin
        meta_36_valid_1 <= _GEN_2601;
      end
    end else begin
      meta_36_valid_1 <= _GEN_2601;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_36_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_36_lru <= _GEN_8272;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_37_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_37_valid_0 <= _GEN_2090;
        end else begin
          meta_37_valid_0 <= _GEN_7285;
        end
      end else begin
        meta_37_valid_0 <= _GEN_2090;
      end
    end else begin
      meta_37_valid_0 <= _GEN_2090;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_37_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_37_valid_1 <= _GEN_2602;
        end else begin
          meta_37_valid_1 <= _GEN_7286;
        end
      end else begin
        meta_37_valid_1 <= _GEN_2602;
      end
    end else begin
      meta_37_valid_1 <= _GEN_2602;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_37_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_37_lru <= _GEN_8273;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_38_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_38_valid_0 <= _GEN_2091;
        end else begin
          meta_38_valid_0 <= _GEN_7287;
        end
      end else begin
        meta_38_valid_0 <= _GEN_2091;
      end
    end else begin
      meta_38_valid_0 <= _GEN_2091;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_38_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_38_valid_1 <= _GEN_2603;
        end else begin
          meta_38_valid_1 <= _GEN_7288;
        end
      end else begin
        meta_38_valid_1 <= _GEN_2603;
      end
    end else begin
      meta_38_valid_1 <= _GEN_2603;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_38_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_38_lru <= _GEN_8274;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_39_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_39_valid_0 <= _GEN_2092;
        end else begin
          meta_39_valid_0 <= _GEN_7289;
        end
      end else begin
        meta_39_valid_0 <= _GEN_2092;
      end
    end else begin
      meta_39_valid_0 <= _GEN_2092;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_39_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_39_valid_1 <= _GEN_2604;
        end else begin
          meta_39_valid_1 <= _GEN_7290;
        end
      end else begin
        meta_39_valid_1 <= _GEN_2604;
      end
    end else begin
      meta_39_valid_1 <= _GEN_2604;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_39_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_39_lru <= _GEN_8275;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_40_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_40_valid_0 <= _GEN_2093;
        end else begin
          meta_40_valid_0 <= _GEN_7291;
        end
      end else begin
        meta_40_valid_0 <= _GEN_2093;
      end
    end else begin
      meta_40_valid_0 <= _GEN_2093;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_40_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_40_valid_1 <= _GEN_2605;
        end else begin
          meta_40_valid_1 <= _GEN_7292;
        end
      end else begin
        meta_40_valid_1 <= _GEN_2605;
      end
    end else begin
      meta_40_valid_1 <= _GEN_2605;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_40_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_40_lru <= _GEN_8276;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_41_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_41_valid_0 <= _GEN_2094;
        end else begin
          meta_41_valid_0 <= _GEN_7293;
        end
      end else begin
        meta_41_valid_0 <= _GEN_2094;
      end
    end else begin
      meta_41_valid_0 <= _GEN_2094;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_41_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_41_valid_1 <= _GEN_2606;
        end else begin
          meta_41_valid_1 <= _GEN_7294;
        end
      end else begin
        meta_41_valid_1 <= _GEN_2606;
      end
    end else begin
      meta_41_valid_1 <= _GEN_2606;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_41_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_41_lru <= _GEN_8277;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_42_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_42_valid_0 <= _GEN_2095;
        end else begin
          meta_42_valid_0 <= _GEN_7295;
        end
      end else begin
        meta_42_valid_0 <= _GEN_2095;
      end
    end else begin
      meta_42_valid_0 <= _GEN_2095;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_42_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_42_valid_1 <= _GEN_2607;
        end else begin
          meta_42_valid_1 <= _GEN_7296;
        end
      end else begin
        meta_42_valid_1 <= _GEN_2607;
      end
    end else begin
      meta_42_valid_1 <= _GEN_2607;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_42_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_42_lru <= _GEN_8278;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_43_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_43_valid_0 <= _GEN_2096;
        end else begin
          meta_43_valid_0 <= _GEN_7297;
        end
      end else begin
        meta_43_valid_0 <= _GEN_2096;
      end
    end else begin
      meta_43_valid_0 <= _GEN_2096;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_43_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_43_valid_1 <= _GEN_2608;
        end else begin
          meta_43_valid_1 <= _GEN_7298;
        end
      end else begin
        meta_43_valid_1 <= _GEN_2608;
      end
    end else begin
      meta_43_valid_1 <= _GEN_2608;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_43_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_43_lru <= _GEN_8279;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_44_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_44_valid_0 <= _GEN_2097;
        end else begin
          meta_44_valid_0 <= _GEN_7299;
        end
      end else begin
        meta_44_valid_0 <= _GEN_2097;
      end
    end else begin
      meta_44_valid_0 <= _GEN_2097;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_44_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_44_valid_1 <= _GEN_2609;
        end else begin
          meta_44_valid_1 <= _GEN_7300;
        end
      end else begin
        meta_44_valid_1 <= _GEN_2609;
      end
    end else begin
      meta_44_valid_1 <= _GEN_2609;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_44_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_44_lru <= _GEN_8280;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_45_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_45_valid_0 <= _GEN_2098;
        end else begin
          meta_45_valid_0 <= _GEN_7301;
        end
      end else begin
        meta_45_valid_0 <= _GEN_2098;
      end
    end else begin
      meta_45_valid_0 <= _GEN_2098;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_45_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_45_valid_1 <= _GEN_2610;
        end else begin
          meta_45_valid_1 <= _GEN_7302;
        end
      end else begin
        meta_45_valid_1 <= _GEN_2610;
      end
    end else begin
      meta_45_valid_1 <= _GEN_2610;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_45_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_45_lru <= _GEN_8281;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_46_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_46_valid_0 <= _GEN_2099;
        end else begin
          meta_46_valid_0 <= _GEN_7303;
        end
      end else begin
        meta_46_valid_0 <= _GEN_2099;
      end
    end else begin
      meta_46_valid_0 <= _GEN_2099;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_46_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_46_valid_1 <= _GEN_2611;
        end else begin
          meta_46_valid_1 <= _GEN_7304;
        end
      end else begin
        meta_46_valid_1 <= _GEN_2611;
      end
    end else begin
      meta_46_valid_1 <= _GEN_2611;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_46_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_46_lru <= _GEN_8282;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_47_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_47_valid_0 <= _GEN_2100;
        end else begin
          meta_47_valid_0 <= _GEN_7305;
        end
      end else begin
        meta_47_valid_0 <= _GEN_2100;
      end
    end else begin
      meta_47_valid_0 <= _GEN_2100;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_47_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_47_valid_1 <= _GEN_2612;
        end else begin
          meta_47_valid_1 <= _GEN_7306;
        end
      end else begin
        meta_47_valid_1 <= _GEN_2612;
      end
    end else begin
      meta_47_valid_1 <= _GEN_2612;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_47_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_47_lru <= _GEN_8283;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_48_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_48_valid_0 <= _GEN_2101;
        end else begin
          meta_48_valid_0 <= _GEN_7307;
        end
      end else begin
        meta_48_valid_0 <= _GEN_2101;
      end
    end else begin
      meta_48_valid_0 <= _GEN_2101;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_48_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_48_valid_1 <= _GEN_2613;
        end else begin
          meta_48_valid_1 <= _GEN_7308;
        end
      end else begin
        meta_48_valid_1 <= _GEN_2613;
      end
    end else begin
      meta_48_valid_1 <= _GEN_2613;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_48_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_48_lru <= _GEN_8284;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_49_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_49_valid_0 <= _GEN_2102;
        end else begin
          meta_49_valid_0 <= _GEN_7309;
        end
      end else begin
        meta_49_valid_0 <= _GEN_2102;
      end
    end else begin
      meta_49_valid_0 <= _GEN_2102;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_49_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_49_valid_1 <= _GEN_2614;
        end else begin
          meta_49_valid_1 <= _GEN_7310;
        end
      end else begin
        meta_49_valid_1 <= _GEN_2614;
      end
    end else begin
      meta_49_valid_1 <= _GEN_2614;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_49_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_49_lru <= _GEN_8285;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_50_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_50_valid_0 <= _GEN_2103;
        end else begin
          meta_50_valid_0 <= _GEN_7311;
        end
      end else begin
        meta_50_valid_0 <= _GEN_2103;
      end
    end else begin
      meta_50_valid_0 <= _GEN_2103;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_50_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_50_valid_1 <= _GEN_2615;
        end else begin
          meta_50_valid_1 <= _GEN_7312;
        end
      end else begin
        meta_50_valid_1 <= _GEN_2615;
      end
    end else begin
      meta_50_valid_1 <= _GEN_2615;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_50_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_50_lru <= _GEN_8286;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_51_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_51_valid_0 <= _GEN_2104;
        end else begin
          meta_51_valid_0 <= _GEN_7313;
        end
      end else begin
        meta_51_valid_0 <= _GEN_2104;
      end
    end else begin
      meta_51_valid_0 <= _GEN_2104;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_51_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_51_valid_1 <= _GEN_2616;
        end else begin
          meta_51_valid_1 <= _GEN_7314;
        end
      end else begin
        meta_51_valid_1 <= _GEN_2616;
      end
    end else begin
      meta_51_valid_1 <= _GEN_2616;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_51_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_51_lru <= _GEN_8287;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_52_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_52_valid_0 <= _GEN_2105;
        end else begin
          meta_52_valid_0 <= _GEN_7315;
        end
      end else begin
        meta_52_valid_0 <= _GEN_2105;
      end
    end else begin
      meta_52_valid_0 <= _GEN_2105;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_52_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_52_valid_1 <= _GEN_2617;
        end else begin
          meta_52_valid_1 <= _GEN_7316;
        end
      end else begin
        meta_52_valid_1 <= _GEN_2617;
      end
    end else begin
      meta_52_valid_1 <= _GEN_2617;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_52_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_52_lru <= _GEN_8288;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_53_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_53_valid_0 <= _GEN_2106;
        end else begin
          meta_53_valid_0 <= _GEN_7317;
        end
      end else begin
        meta_53_valid_0 <= _GEN_2106;
      end
    end else begin
      meta_53_valid_0 <= _GEN_2106;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_53_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_53_valid_1 <= _GEN_2618;
        end else begin
          meta_53_valid_1 <= _GEN_7318;
        end
      end else begin
        meta_53_valid_1 <= _GEN_2618;
      end
    end else begin
      meta_53_valid_1 <= _GEN_2618;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_53_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_53_lru <= _GEN_8289;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_54_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_54_valid_0 <= _GEN_2107;
        end else begin
          meta_54_valid_0 <= _GEN_7319;
        end
      end else begin
        meta_54_valid_0 <= _GEN_2107;
      end
    end else begin
      meta_54_valid_0 <= _GEN_2107;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_54_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_54_valid_1 <= _GEN_2619;
        end else begin
          meta_54_valid_1 <= _GEN_7320;
        end
      end else begin
        meta_54_valid_1 <= _GEN_2619;
      end
    end else begin
      meta_54_valid_1 <= _GEN_2619;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_54_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_54_lru <= _GEN_8290;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_55_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_55_valid_0 <= _GEN_2108;
        end else begin
          meta_55_valid_0 <= _GEN_7321;
        end
      end else begin
        meta_55_valid_0 <= _GEN_2108;
      end
    end else begin
      meta_55_valid_0 <= _GEN_2108;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_55_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_55_valid_1 <= _GEN_2620;
        end else begin
          meta_55_valid_1 <= _GEN_7322;
        end
      end else begin
        meta_55_valid_1 <= _GEN_2620;
      end
    end else begin
      meta_55_valid_1 <= _GEN_2620;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_55_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_55_lru <= _GEN_8291;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_56_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_56_valid_0 <= _GEN_2109;
        end else begin
          meta_56_valid_0 <= _GEN_7323;
        end
      end else begin
        meta_56_valid_0 <= _GEN_2109;
      end
    end else begin
      meta_56_valid_0 <= _GEN_2109;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_56_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_56_valid_1 <= _GEN_2621;
        end else begin
          meta_56_valid_1 <= _GEN_7324;
        end
      end else begin
        meta_56_valid_1 <= _GEN_2621;
      end
    end else begin
      meta_56_valid_1 <= _GEN_2621;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_56_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_56_lru <= _GEN_8292;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_57_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_57_valid_0 <= _GEN_2110;
        end else begin
          meta_57_valid_0 <= _GEN_7325;
        end
      end else begin
        meta_57_valid_0 <= _GEN_2110;
      end
    end else begin
      meta_57_valid_0 <= _GEN_2110;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_57_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_57_valid_1 <= _GEN_2622;
        end else begin
          meta_57_valid_1 <= _GEN_7326;
        end
      end else begin
        meta_57_valid_1 <= _GEN_2622;
      end
    end else begin
      meta_57_valid_1 <= _GEN_2622;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_57_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_57_lru <= _GEN_8293;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_58_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_58_valid_0 <= _GEN_2111;
        end else begin
          meta_58_valid_0 <= _GEN_7327;
        end
      end else begin
        meta_58_valid_0 <= _GEN_2111;
      end
    end else begin
      meta_58_valid_0 <= _GEN_2111;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_58_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_58_valid_1 <= _GEN_2623;
        end else begin
          meta_58_valid_1 <= _GEN_7328;
        end
      end else begin
        meta_58_valid_1 <= _GEN_2623;
      end
    end else begin
      meta_58_valid_1 <= _GEN_2623;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_58_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_58_lru <= _GEN_8294;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_59_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_59_valid_0 <= _GEN_2112;
        end else begin
          meta_59_valid_0 <= _GEN_7329;
        end
      end else begin
        meta_59_valid_0 <= _GEN_2112;
      end
    end else begin
      meta_59_valid_0 <= _GEN_2112;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_59_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_59_valid_1 <= _GEN_2624;
        end else begin
          meta_59_valid_1 <= _GEN_7330;
        end
      end else begin
        meta_59_valid_1 <= _GEN_2624;
      end
    end else begin
      meta_59_valid_1 <= _GEN_2624;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_59_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_59_lru <= _GEN_8295;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_60_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_60_valid_0 <= _GEN_2113;
        end else begin
          meta_60_valid_0 <= _GEN_7331;
        end
      end else begin
        meta_60_valid_0 <= _GEN_2113;
      end
    end else begin
      meta_60_valid_0 <= _GEN_2113;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_60_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_60_valid_1 <= _GEN_2625;
        end else begin
          meta_60_valid_1 <= _GEN_7332;
        end
      end else begin
        meta_60_valid_1 <= _GEN_2625;
      end
    end else begin
      meta_60_valid_1 <= _GEN_2625;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_60_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_60_lru <= _GEN_8296;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_61_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_61_valid_0 <= _GEN_2114;
        end else begin
          meta_61_valid_0 <= _GEN_7333;
        end
      end else begin
        meta_61_valid_0 <= _GEN_2114;
      end
    end else begin
      meta_61_valid_0 <= _GEN_2114;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_61_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_61_valid_1 <= _GEN_2626;
        end else begin
          meta_61_valid_1 <= _GEN_7334;
        end
      end else begin
        meta_61_valid_1 <= _GEN_2626;
      end
    end else begin
      meta_61_valid_1 <= _GEN_2626;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_61_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_61_lru <= _GEN_8297;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_62_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_62_valid_0 <= _GEN_2115;
        end else begin
          meta_62_valid_0 <= _GEN_7335;
        end
      end else begin
        meta_62_valid_0 <= _GEN_2115;
      end
    end else begin
      meta_62_valid_0 <= _GEN_2115;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_62_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_62_valid_1 <= _GEN_2627;
        end else begin
          meta_62_valid_1 <= _GEN_7336;
        end
      end else begin
        meta_62_valid_1 <= _GEN_2627;
      end
    end else begin
      meta_62_valid_1 <= _GEN_2627;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_62_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_62_lru <= _GEN_8298;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_63_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_63_valid_0 <= _GEN_2116;
        end else begin
          meta_63_valid_0 <= _GEN_7337;
        end
      end else begin
        meta_63_valid_0 <= _GEN_2116;
      end
    end else begin
      meta_63_valid_0 <= _GEN_2116;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_63_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_63_valid_1 <= _GEN_2628;
        end else begin
          meta_63_valid_1 <= _GEN_7338;
        end
      end else begin
        meta_63_valid_1 <= _GEN_2628;
      end
    end else begin
      meta_63_valid_1 <= _GEN_2628;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_63_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_63_lru <= _GEN_8299;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_64_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_64_valid_0 <= _GEN_2117;
        end else begin
          meta_64_valid_0 <= _GEN_7339;
        end
      end else begin
        meta_64_valid_0 <= _GEN_2117;
      end
    end else begin
      meta_64_valid_0 <= _GEN_2117;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_64_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_64_valid_1 <= _GEN_2629;
        end else begin
          meta_64_valid_1 <= _GEN_7340;
        end
      end else begin
        meta_64_valid_1 <= _GEN_2629;
      end
    end else begin
      meta_64_valid_1 <= _GEN_2629;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_64_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_64_lru <= _GEN_8300;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_65_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_65_valid_0 <= _GEN_2118;
        end else begin
          meta_65_valid_0 <= _GEN_7341;
        end
      end else begin
        meta_65_valid_0 <= _GEN_2118;
      end
    end else begin
      meta_65_valid_0 <= _GEN_2118;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_65_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_65_valid_1 <= _GEN_2630;
        end else begin
          meta_65_valid_1 <= _GEN_7342;
        end
      end else begin
        meta_65_valid_1 <= _GEN_2630;
      end
    end else begin
      meta_65_valid_1 <= _GEN_2630;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_65_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_65_lru <= _GEN_8301;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_66_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_66_valid_0 <= _GEN_2119;
        end else begin
          meta_66_valid_0 <= _GEN_7343;
        end
      end else begin
        meta_66_valid_0 <= _GEN_2119;
      end
    end else begin
      meta_66_valid_0 <= _GEN_2119;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_66_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_66_valid_1 <= _GEN_2631;
        end else begin
          meta_66_valid_1 <= _GEN_7344;
        end
      end else begin
        meta_66_valid_1 <= _GEN_2631;
      end
    end else begin
      meta_66_valid_1 <= _GEN_2631;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_66_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_66_lru <= _GEN_8302;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_67_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_67_valid_0 <= _GEN_2120;
        end else begin
          meta_67_valid_0 <= _GEN_7345;
        end
      end else begin
        meta_67_valid_0 <= _GEN_2120;
      end
    end else begin
      meta_67_valid_0 <= _GEN_2120;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_67_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_67_valid_1 <= _GEN_2632;
        end else begin
          meta_67_valid_1 <= _GEN_7346;
        end
      end else begin
        meta_67_valid_1 <= _GEN_2632;
      end
    end else begin
      meta_67_valid_1 <= _GEN_2632;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_67_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_67_lru <= _GEN_8303;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_68_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_68_valid_0 <= _GEN_2121;
        end else begin
          meta_68_valid_0 <= _GEN_7347;
        end
      end else begin
        meta_68_valid_0 <= _GEN_2121;
      end
    end else begin
      meta_68_valid_0 <= _GEN_2121;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_68_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_68_valid_1 <= _GEN_2633;
        end else begin
          meta_68_valid_1 <= _GEN_7348;
        end
      end else begin
        meta_68_valid_1 <= _GEN_2633;
      end
    end else begin
      meta_68_valid_1 <= _GEN_2633;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_68_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_68_lru <= _GEN_8304;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_69_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_69_valid_0 <= _GEN_2122;
        end else begin
          meta_69_valid_0 <= _GEN_7349;
        end
      end else begin
        meta_69_valid_0 <= _GEN_2122;
      end
    end else begin
      meta_69_valid_0 <= _GEN_2122;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_69_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_69_valid_1 <= _GEN_2634;
        end else begin
          meta_69_valid_1 <= _GEN_7350;
        end
      end else begin
        meta_69_valid_1 <= _GEN_2634;
      end
    end else begin
      meta_69_valid_1 <= _GEN_2634;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_69_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_69_lru <= _GEN_8305;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_70_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_70_valid_0 <= _GEN_2123;
        end else begin
          meta_70_valid_0 <= _GEN_7351;
        end
      end else begin
        meta_70_valid_0 <= _GEN_2123;
      end
    end else begin
      meta_70_valid_0 <= _GEN_2123;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_70_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_70_valid_1 <= _GEN_2635;
        end else begin
          meta_70_valid_1 <= _GEN_7352;
        end
      end else begin
        meta_70_valid_1 <= _GEN_2635;
      end
    end else begin
      meta_70_valid_1 <= _GEN_2635;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_70_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_70_lru <= _GEN_8306;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_71_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_71_valid_0 <= _GEN_2124;
        end else begin
          meta_71_valid_0 <= _GEN_7353;
        end
      end else begin
        meta_71_valid_0 <= _GEN_2124;
      end
    end else begin
      meta_71_valid_0 <= _GEN_2124;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_71_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_71_valid_1 <= _GEN_2636;
        end else begin
          meta_71_valid_1 <= _GEN_7354;
        end
      end else begin
        meta_71_valid_1 <= _GEN_2636;
      end
    end else begin
      meta_71_valid_1 <= _GEN_2636;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_71_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_71_lru <= _GEN_8307;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_72_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_72_valid_0 <= _GEN_2125;
        end else begin
          meta_72_valid_0 <= _GEN_7355;
        end
      end else begin
        meta_72_valid_0 <= _GEN_2125;
      end
    end else begin
      meta_72_valid_0 <= _GEN_2125;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_72_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_72_valid_1 <= _GEN_2637;
        end else begin
          meta_72_valid_1 <= _GEN_7356;
        end
      end else begin
        meta_72_valid_1 <= _GEN_2637;
      end
    end else begin
      meta_72_valid_1 <= _GEN_2637;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_72_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_72_lru <= _GEN_8308;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_73_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_73_valid_0 <= _GEN_2126;
        end else begin
          meta_73_valid_0 <= _GEN_7357;
        end
      end else begin
        meta_73_valid_0 <= _GEN_2126;
      end
    end else begin
      meta_73_valid_0 <= _GEN_2126;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_73_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_73_valid_1 <= _GEN_2638;
        end else begin
          meta_73_valid_1 <= _GEN_7358;
        end
      end else begin
        meta_73_valid_1 <= _GEN_2638;
      end
    end else begin
      meta_73_valid_1 <= _GEN_2638;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_73_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_73_lru <= _GEN_8309;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_74_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_74_valid_0 <= _GEN_2127;
        end else begin
          meta_74_valid_0 <= _GEN_7359;
        end
      end else begin
        meta_74_valid_0 <= _GEN_2127;
      end
    end else begin
      meta_74_valid_0 <= _GEN_2127;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_74_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_74_valid_1 <= _GEN_2639;
        end else begin
          meta_74_valid_1 <= _GEN_7360;
        end
      end else begin
        meta_74_valid_1 <= _GEN_2639;
      end
    end else begin
      meta_74_valid_1 <= _GEN_2639;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_74_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_74_lru <= _GEN_8310;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_75_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_75_valid_0 <= _GEN_2128;
        end else begin
          meta_75_valid_0 <= _GEN_7361;
        end
      end else begin
        meta_75_valid_0 <= _GEN_2128;
      end
    end else begin
      meta_75_valid_0 <= _GEN_2128;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_75_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_75_valid_1 <= _GEN_2640;
        end else begin
          meta_75_valid_1 <= _GEN_7362;
        end
      end else begin
        meta_75_valid_1 <= _GEN_2640;
      end
    end else begin
      meta_75_valid_1 <= _GEN_2640;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_75_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_75_lru <= _GEN_8311;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_76_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_76_valid_0 <= _GEN_2129;
        end else begin
          meta_76_valid_0 <= _GEN_7363;
        end
      end else begin
        meta_76_valid_0 <= _GEN_2129;
      end
    end else begin
      meta_76_valid_0 <= _GEN_2129;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_76_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_76_valid_1 <= _GEN_2641;
        end else begin
          meta_76_valid_1 <= _GEN_7364;
        end
      end else begin
        meta_76_valid_1 <= _GEN_2641;
      end
    end else begin
      meta_76_valid_1 <= _GEN_2641;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_76_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_76_lru <= _GEN_8312;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_77_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_77_valid_0 <= _GEN_2130;
        end else begin
          meta_77_valid_0 <= _GEN_7365;
        end
      end else begin
        meta_77_valid_0 <= _GEN_2130;
      end
    end else begin
      meta_77_valid_0 <= _GEN_2130;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_77_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_77_valid_1 <= _GEN_2642;
        end else begin
          meta_77_valid_1 <= _GEN_7366;
        end
      end else begin
        meta_77_valid_1 <= _GEN_2642;
      end
    end else begin
      meta_77_valid_1 <= _GEN_2642;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_77_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_77_lru <= _GEN_8313;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_78_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_78_valid_0 <= _GEN_2131;
        end else begin
          meta_78_valid_0 <= _GEN_7367;
        end
      end else begin
        meta_78_valid_0 <= _GEN_2131;
      end
    end else begin
      meta_78_valid_0 <= _GEN_2131;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_78_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_78_valid_1 <= _GEN_2643;
        end else begin
          meta_78_valid_1 <= _GEN_7368;
        end
      end else begin
        meta_78_valid_1 <= _GEN_2643;
      end
    end else begin
      meta_78_valid_1 <= _GEN_2643;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_78_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_78_lru <= _GEN_8314;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_79_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_79_valid_0 <= _GEN_2132;
        end else begin
          meta_79_valid_0 <= _GEN_7369;
        end
      end else begin
        meta_79_valid_0 <= _GEN_2132;
      end
    end else begin
      meta_79_valid_0 <= _GEN_2132;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_79_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_79_valid_1 <= _GEN_2644;
        end else begin
          meta_79_valid_1 <= _GEN_7370;
        end
      end else begin
        meta_79_valid_1 <= _GEN_2644;
      end
    end else begin
      meta_79_valid_1 <= _GEN_2644;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_79_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_79_lru <= _GEN_8315;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_80_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_80_valid_0 <= _GEN_2133;
        end else begin
          meta_80_valid_0 <= _GEN_7371;
        end
      end else begin
        meta_80_valid_0 <= _GEN_2133;
      end
    end else begin
      meta_80_valid_0 <= _GEN_2133;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_80_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_80_valid_1 <= _GEN_2645;
        end else begin
          meta_80_valid_1 <= _GEN_7372;
        end
      end else begin
        meta_80_valid_1 <= _GEN_2645;
      end
    end else begin
      meta_80_valid_1 <= _GEN_2645;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_80_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_80_lru <= _GEN_8316;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_81_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_81_valid_0 <= _GEN_2134;
        end else begin
          meta_81_valid_0 <= _GEN_7373;
        end
      end else begin
        meta_81_valid_0 <= _GEN_2134;
      end
    end else begin
      meta_81_valid_0 <= _GEN_2134;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_81_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_81_valid_1 <= _GEN_2646;
        end else begin
          meta_81_valid_1 <= _GEN_7374;
        end
      end else begin
        meta_81_valid_1 <= _GEN_2646;
      end
    end else begin
      meta_81_valid_1 <= _GEN_2646;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_81_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_81_lru <= _GEN_8317;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_82_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_82_valid_0 <= _GEN_2135;
        end else begin
          meta_82_valid_0 <= _GEN_7375;
        end
      end else begin
        meta_82_valid_0 <= _GEN_2135;
      end
    end else begin
      meta_82_valid_0 <= _GEN_2135;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_82_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_82_valid_1 <= _GEN_2647;
        end else begin
          meta_82_valid_1 <= _GEN_7376;
        end
      end else begin
        meta_82_valid_1 <= _GEN_2647;
      end
    end else begin
      meta_82_valid_1 <= _GEN_2647;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_82_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_82_lru <= _GEN_8318;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_83_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_83_valid_0 <= _GEN_2136;
        end else begin
          meta_83_valid_0 <= _GEN_7377;
        end
      end else begin
        meta_83_valid_0 <= _GEN_2136;
      end
    end else begin
      meta_83_valid_0 <= _GEN_2136;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_83_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_83_valid_1 <= _GEN_2648;
        end else begin
          meta_83_valid_1 <= _GEN_7378;
        end
      end else begin
        meta_83_valid_1 <= _GEN_2648;
      end
    end else begin
      meta_83_valid_1 <= _GEN_2648;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_83_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_83_lru <= _GEN_8319;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_84_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_84_valid_0 <= _GEN_2137;
        end else begin
          meta_84_valid_0 <= _GEN_7379;
        end
      end else begin
        meta_84_valid_0 <= _GEN_2137;
      end
    end else begin
      meta_84_valid_0 <= _GEN_2137;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_84_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_84_valid_1 <= _GEN_2649;
        end else begin
          meta_84_valid_1 <= _GEN_7380;
        end
      end else begin
        meta_84_valid_1 <= _GEN_2649;
      end
    end else begin
      meta_84_valid_1 <= _GEN_2649;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_84_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_84_lru <= _GEN_8320;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_85_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_85_valid_0 <= _GEN_2138;
        end else begin
          meta_85_valid_0 <= _GEN_7381;
        end
      end else begin
        meta_85_valid_0 <= _GEN_2138;
      end
    end else begin
      meta_85_valid_0 <= _GEN_2138;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_85_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_85_valid_1 <= _GEN_2650;
        end else begin
          meta_85_valid_1 <= _GEN_7382;
        end
      end else begin
        meta_85_valid_1 <= _GEN_2650;
      end
    end else begin
      meta_85_valid_1 <= _GEN_2650;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_85_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_85_lru <= _GEN_8321;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_86_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_86_valid_0 <= _GEN_2139;
        end else begin
          meta_86_valid_0 <= _GEN_7383;
        end
      end else begin
        meta_86_valid_0 <= _GEN_2139;
      end
    end else begin
      meta_86_valid_0 <= _GEN_2139;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_86_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_86_valid_1 <= _GEN_2651;
        end else begin
          meta_86_valid_1 <= _GEN_7384;
        end
      end else begin
        meta_86_valid_1 <= _GEN_2651;
      end
    end else begin
      meta_86_valid_1 <= _GEN_2651;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_86_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_86_lru <= _GEN_8322;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_87_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_87_valid_0 <= _GEN_2140;
        end else begin
          meta_87_valid_0 <= _GEN_7385;
        end
      end else begin
        meta_87_valid_0 <= _GEN_2140;
      end
    end else begin
      meta_87_valid_0 <= _GEN_2140;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_87_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_87_valid_1 <= _GEN_2652;
        end else begin
          meta_87_valid_1 <= _GEN_7386;
        end
      end else begin
        meta_87_valid_1 <= _GEN_2652;
      end
    end else begin
      meta_87_valid_1 <= _GEN_2652;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_87_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_87_lru <= _GEN_8323;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_88_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_88_valid_0 <= _GEN_2141;
        end else begin
          meta_88_valid_0 <= _GEN_7387;
        end
      end else begin
        meta_88_valid_0 <= _GEN_2141;
      end
    end else begin
      meta_88_valid_0 <= _GEN_2141;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_88_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_88_valid_1 <= _GEN_2653;
        end else begin
          meta_88_valid_1 <= _GEN_7388;
        end
      end else begin
        meta_88_valid_1 <= _GEN_2653;
      end
    end else begin
      meta_88_valid_1 <= _GEN_2653;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_88_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_88_lru <= _GEN_8324;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_89_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_89_valid_0 <= _GEN_2142;
        end else begin
          meta_89_valid_0 <= _GEN_7389;
        end
      end else begin
        meta_89_valid_0 <= _GEN_2142;
      end
    end else begin
      meta_89_valid_0 <= _GEN_2142;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_89_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_89_valid_1 <= _GEN_2654;
        end else begin
          meta_89_valid_1 <= _GEN_7390;
        end
      end else begin
        meta_89_valid_1 <= _GEN_2654;
      end
    end else begin
      meta_89_valid_1 <= _GEN_2654;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_89_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_89_lru <= _GEN_8325;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_90_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_90_valid_0 <= _GEN_2143;
        end else begin
          meta_90_valid_0 <= _GEN_7391;
        end
      end else begin
        meta_90_valid_0 <= _GEN_2143;
      end
    end else begin
      meta_90_valid_0 <= _GEN_2143;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_90_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_90_valid_1 <= _GEN_2655;
        end else begin
          meta_90_valid_1 <= _GEN_7392;
        end
      end else begin
        meta_90_valid_1 <= _GEN_2655;
      end
    end else begin
      meta_90_valid_1 <= _GEN_2655;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_90_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_90_lru <= _GEN_8326;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_91_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_91_valid_0 <= _GEN_2144;
        end else begin
          meta_91_valid_0 <= _GEN_7393;
        end
      end else begin
        meta_91_valid_0 <= _GEN_2144;
      end
    end else begin
      meta_91_valid_0 <= _GEN_2144;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_91_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_91_valid_1 <= _GEN_2656;
        end else begin
          meta_91_valid_1 <= _GEN_7394;
        end
      end else begin
        meta_91_valid_1 <= _GEN_2656;
      end
    end else begin
      meta_91_valid_1 <= _GEN_2656;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_91_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_91_lru <= _GEN_8327;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_92_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_92_valid_0 <= _GEN_2145;
        end else begin
          meta_92_valid_0 <= _GEN_7395;
        end
      end else begin
        meta_92_valid_0 <= _GEN_2145;
      end
    end else begin
      meta_92_valid_0 <= _GEN_2145;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_92_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_92_valid_1 <= _GEN_2657;
        end else begin
          meta_92_valid_1 <= _GEN_7396;
        end
      end else begin
        meta_92_valid_1 <= _GEN_2657;
      end
    end else begin
      meta_92_valid_1 <= _GEN_2657;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_92_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_92_lru <= _GEN_8328;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_93_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_93_valid_0 <= _GEN_2146;
        end else begin
          meta_93_valid_0 <= _GEN_7397;
        end
      end else begin
        meta_93_valid_0 <= _GEN_2146;
      end
    end else begin
      meta_93_valid_0 <= _GEN_2146;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_93_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_93_valid_1 <= _GEN_2658;
        end else begin
          meta_93_valid_1 <= _GEN_7398;
        end
      end else begin
        meta_93_valid_1 <= _GEN_2658;
      end
    end else begin
      meta_93_valid_1 <= _GEN_2658;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_93_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_93_lru <= _GEN_8329;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_94_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_94_valid_0 <= _GEN_2147;
        end else begin
          meta_94_valid_0 <= _GEN_7399;
        end
      end else begin
        meta_94_valid_0 <= _GEN_2147;
      end
    end else begin
      meta_94_valid_0 <= _GEN_2147;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_94_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_94_valid_1 <= _GEN_2659;
        end else begin
          meta_94_valid_1 <= _GEN_7400;
        end
      end else begin
        meta_94_valid_1 <= _GEN_2659;
      end
    end else begin
      meta_94_valid_1 <= _GEN_2659;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_94_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_94_lru <= _GEN_8330;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_95_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_95_valid_0 <= _GEN_2148;
        end else begin
          meta_95_valid_0 <= _GEN_7401;
        end
      end else begin
        meta_95_valid_0 <= _GEN_2148;
      end
    end else begin
      meta_95_valid_0 <= _GEN_2148;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_95_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_95_valid_1 <= _GEN_2660;
        end else begin
          meta_95_valid_1 <= _GEN_7402;
        end
      end else begin
        meta_95_valid_1 <= _GEN_2660;
      end
    end else begin
      meta_95_valid_1 <= _GEN_2660;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_95_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_95_lru <= _GEN_8331;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_96_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_96_valid_0 <= _GEN_2149;
        end else begin
          meta_96_valid_0 <= _GEN_7403;
        end
      end else begin
        meta_96_valid_0 <= _GEN_2149;
      end
    end else begin
      meta_96_valid_0 <= _GEN_2149;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_96_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_96_valid_1 <= _GEN_2661;
        end else begin
          meta_96_valid_1 <= _GEN_7404;
        end
      end else begin
        meta_96_valid_1 <= _GEN_2661;
      end
    end else begin
      meta_96_valid_1 <= _GEN_2661;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_96_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_96_lru <= _GEN_8332;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_97_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_97_valid_0 <= _GEN_2150;
        end else begin
          meta_97_valid_0 <= _GEN_7405;
        end
      end else begin
        meta_97_valid_0 <= _GEN_2150;
      end
    end else begin
      meta_97_valid_0 <= _GEN_2150;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_97_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_97_valid_1 <= _GEN_2662;
        end else begin
          meta_97_valid_1 <= _GEN_7406;
        end
      end else begin
        meta_97_valid_1 <= _GEN_2662;
      end
    end else begin
      meta_97_valid_1 <= _GEN_2662;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_97_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_97_lru <= _GEN_8333;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_98_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_98_valid_0 <= _GEN_2151;
        end else begin
          meta_98_valid_0 <= _GEN_7407;
        end
      end else begin
        meta_98_valid_0 <= _GEN_2151;
      end
    end else begin
      meta_98_valid_0 <= _GEN_2151;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_98_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_98_valid_1 <= _GEN_2663;
        end else begin
          meta_98_valid_1 <= _GEN_7408;
        end
      end else begin
        meta_98_valid_1 <= _GEN_2663;
      end
    end else begin
      meta_98_valid_1 <= _GEN_2663;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_98_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_98_lru <= _GEN_8334;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_99_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_99_valid_0 <= _GEN_2152;
        end else begin
          meta_99_valid_0 <= _GEN_7409;
        end
      end else begin
        meta_99_valid_0 <= _GEN_2152;
      end
    end else begin
      meta_99_valid_0 <= _GEN_2152;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_99_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_99_valid_1 <= _GEN_2664;
        end else begin
          meta_99_valid_1 <= _GEN_7410;
        end
      end else begin
        meta_99_valid_1 <= _GEN_2664;
      end
    end else begin
      meta_99_valid_1 <= _GEN_2664;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_99_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_99_lru <= _GEN_8335;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_100_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_100_valid_0 <= _GEN_2153;
        end else begin
          meta_100_valid_0 <= _GEN_7411;
        end
      end else begin
        meta_100_valid_0 <= _GEN_2153;
      end
    end else begin
      meta_100_valid_0 <= _GEN_2153;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_100_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_100_valid_1 <= _GEN_2665;
        end else begin
          meta_100_valid_1 <= _GEN_7412;
        end
      end else begin
        meta_100_valid_1 <= _GEN_2665;
      end
    end else begin
      meta_100_valid_1 <= _GEN_2665;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_100_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_100_lru <= _GEN_8336;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_101_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_101_valid_0 <= _GEN_2154;
        end else begin
          meta_101_valid_0 <= _GEN_7413;
        end
      end else begin
        meta_101_valid_0 <= _GEN_2154;
      end
    end else begin
      meta_101_valid_0 <= _GEN_2154;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_101_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_101_valid_1 <= _GEN_2666;
        end else begin
          meta_101_valid_1 <= _GEN_7414;
        end
      end else begin
        meta_101_valid_1 <= _GEN_2666;
      end
    end else begin
      meta_101_valid_1 <= _GEN_2666;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_101_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_101_lru <= _GEN_8337;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_102_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_102_valid_0 <= _GEN_2155;
        end else begin
          meta_102_valid_0 <= _GEN_7415;
        end
      end else begin
        meta_102_valid_0 <= _GEN_2155;
      end
    end else begin
      meta_102_valid_0 <= _GEN_2155;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_102_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_102_valid_1 <= _GEN_2667;
        end else begin
          meta_102_valid_1 <= _GEN_7416;
        end
      end else begin
        meta_102_valid_1 <= _GEN_2667;
      end
    end else begin
      meta_102_valid_1 <= _GEN_2667;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_102_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_102_lru <= _GEN_8338;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_103_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_103_valid_0 <= _GEN_2156;
        end else begin
          meta_103_valid_0 <= _GEN_7417;
        end
      end else begin
        meta_103_valid_0 <= _GEN_2156;
      end
    end else begin
      meta_103_valid_0 <= _GEN_2156;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_103_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_103_valid_1 <= _GEN_2668;
        end else begin
          meta_103_valid_1 <= _GEN_7418;
        end
      end else begin
        meta_103_valid_1 <= _GEN_2668;
      end
    end else begin
      meta_103_valid_1 <= _GEN_2668;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_103_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_103_lru <= _GEN_8339;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_104_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_104_valid_0 <= _GEN_2157;
        end else begin
          meta_104_valid_0 <= _GEN_7419;
        end
      end else begin
        meta_104_valid_0 <= _GEN_2157;
      end
    end else begin
      meta_104_valid_0 <= _GEN_2157;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_104_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_104_valid_1 <= _GEN_2669;
        end else begin
          meta_104_valid_1 <= _GEN_7420;
        end
      end else begin
        meta_104_valid_1 <= _GEN_2669;
      end
    end else begin
      meta_104_valid_1 <= _GEN_2669;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_104_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_104_lru <= _GEN_8340;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_105_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_105_valid_0 <= _GEN_2158;
        end else begin
          meta_105_valid_0 <= _GEN_7421;
        end
      end else begin
        meta_105_valid_0 <= _GEN_2158;
      end
    end else begin
      meta_105_valid_0 <= _GEN_2158;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_105_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_105_valid_1 <= _GEN_2670;
        end else begin
          meta_105_valid_1 <= _GEN_7422;
        end
      end else begin
        meta_105_valid_1 <= _GEN_2670;
      end
    end else begin
      meta_105_valid_1 <= _GEN_2670;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_105_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_105_lru <= _GEN_8341;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_106_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_106_valid_0 <= _GEN_2159;
        end else begin
          meta_106_valid_0 <= _GEN_7423;
        end
      end else begin
        meta_106_valid_0 <= _GEN_2159;
      end
    end else begin
      meta_106_valid_0 <= _GEN_2159;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_106_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_106_valid_1 <= _GEN_2671;
        end else begin
          meta_106_valid_1 <= _GEN_7424;
        end
      end else begin
        meta_106_valid_1 <= _GEN_2671;
      end
    end else begin
      meta_106_valid_1 <= _GEN_2671;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_106_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_106_lru <= _GEN_8342;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_107_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_107_valid_0 <= _GEN_2160;
        end else begin
          meta_107_valid_0 <= _GEN_7425;
        end
      end else begin
        meta_107_valid_0 <= _GEN_2160;
      end
    end else begin
      meta_107_valid_0 <= _GEN_2160;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_107_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_107_valid_1 <= _GEN_2672;
        end else begin
          meta_107_valid_1 <= _GEN_7426;
        end
      end else begin
        meta_107_valid_1 <= _GEN_2672;
      end
    end else begin
      meta_107_valid_1 <= _GEN_2672;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_107_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_107_lru <= _GEN_8343;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_108_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_108_valid_0 <= _GEN_2161;
        end else begin
          meta_108_valid_0 <= _GEN_7427;
        end
      end else begin
        meta_108_valid_0 <= _GEN_2161;
      end
    end else begin
      meta_108_valid_0 <= _GEN_2161;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_108_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_108_valid_1 <= _GEN_2673;
        end else begin
          meta_108_valid_1 <= _GEN_7428;
        end
      end else begin
        meta_108_valid_1 <= _GEN_2673;
      end
    end else begin
      meta_108_valid_1 <= _GEN_2673;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_108_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_108_lru <= _GEN_8344;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_109_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_109_valid_0 <= _GEN_2162;
        end else begin
          meta_109_valid_0 <= _GEN_7429;
        end
      end else begin
        meta_109_valid_0 <= _GEN_2162;
      end
    end else begin
      meta_109_valid_0 <= _GEN_2162;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_109_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_109_valid_1 <= _GEN_2674;
        end else begin
          meta_109_valid_1 <= _GEN_7430;
        end
      end else begin
        meta_109_valid_1 <= _GEN_2674;
      end
    end else begin
      meta_109_valid_1 <= _GEN_2674;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_109_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_109_lru <= _GEN_8345;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_110_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_110_valid_0 <= _GEN_2163;
        end else begin
          meta_110_valid_0 <= _GEN_7431;
        end
      end else begin
        meta_110_valid_0 <= _GEN_2163;
      end
    end else begin
      meta_110_valid_0 <= _GEN_2163;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_110_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_110_valid_1 <= _GEN_2675;
        end else begin
          meta_110_valid_1 <= _GEN_7432;
        end
      end else begin
        meta_110_valid_1 <= _GEN_2675;
      end
    end else begin
      meta_110_valid_1 <= _GEN_2675;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_110_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_110_lru <= _GEN_8346;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_111_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_111_valid_0 <= _GEN_2164;
        end else begin
          meta_111_valid_0 <= _GEN_7433;
        end
      end else begin
        meta_111_valid_0 <= _GEN_2164;
      end
    end else begin
      meta_111_valid_0 <= _GEN_2164;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_111_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_111_valid_1 <= _GEN_2676;
        end else begin
          meta_111_valid_1 <= _GEN_7434;
        end
      end else begin
        meta_111_valid_1 <= _GEN_2676;
      end
    end else begin
      meta_111_valid_1 <= _GEN_2676;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_111_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_111_lru <= _GEN_8347;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_112_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_112_valid_0 <= _GEN_2165;
        end else begin
          meta_112_valid_0 <= _GEN_7435;
        end
      end else begin
        meta_112_valid_0 <= _GEN_2165;
      end
    end else begin
      meta_112_valid_0 <= _GEN_2165;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_112_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_112_valid_1 <= _GEN_2677;
        end else begin
          meta_112_valid_1 <= _GEN_7436;
        end
      end else begin
        meta_112_valid_1 <= _GEN_2677;
      end
    end else begin
      meta_112_valid_1 <= _GEN_2677;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_112_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_112_lru <= _GEN_8348;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_113_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_113_valid_0 <= _GEN_2166;
        end else begin
          meta_113_valid_0 <= _GEN_7437;
        end
      end else begin
        meta_113_valid_0 <= _GEN_2166;
      end
    end else begin
      meta_113_valid_0 <= _GEN_2166;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_113_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_113_valid_1 <= _GEN_2678;
        end else begin
          meta_113_valid_1 <= _GEN_7438;
        end
      end else begin
        meta_113_valid_1 <= _GEN_2678;
      end
    end else begin
      meta_113_valid_1 <= _GEN_2678;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_113_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_113_lru <= _GEN_8349;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_114_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_114_valid_0 <= _GEN_2167;
        end else begin
          meta_114_valid_0 <= _GEN_7439;
        end
      end else begin
        meta_114_valid_0 <= _GEN_2167;
      end
    end else begin
      meta_114_valid_0 <= _GEN_2167;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_114_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_114_valid_1 <= _GEN_2679;
        end else begin
          meta_114_valid_1 <= _GEN_7440;
        end
      end else begin
        meta_114_valid_1 <= _GEN_2679;
      end
    end else begin
      meta_114_valid_1 <= _GEN_2679;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_114_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_114_lru <= _GEN_8350;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_115_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_115_valid_0 <= _GEN_2168;
        end else begin
          meta_115_valid_0 <= _GEN_7441;
        end
      end else begin
        meta_115_valid_0 <= _GEN_2168;
      end
    end else begin
      meta_115_valid_0 <= _GEN_2168;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_115_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_115_valid_1 <= _GEN_2680;
        end else begin
          meta_115_valid_1 <= _GEN_7442;
        end
      end else begin
        meta_115_valid_1 <= _GEN_2680;
      end
    end else begin
      meta_115_valid_1 <= _GEN_2680;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_115_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_115_lru <= _GEN_8351;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_116_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_116_valid_0 <= _GEN_2169;
        end else begin
          meta_116_valid_0 <= _GEN_7443;
        end
      end else begin
        meta_116_valid_0 <= _GEN_2169;
      end
    end else begin
      meta_116_valid_0 <= _GEN_2169;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_116_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_116_valid_1 <= _GEN_2681;
        end else begin
          meta_116_valid_1 <= _GEN_7444;
        end
      end else begin
        meta_116_valid_1 <= _GEN_2681;
      end
    end else begin
      meta_116_valid_1 <= _GEN_2681;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_116_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_116_lru <= _GEN_8352;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_117_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_117_valid_0 <= _GEN_2170;
        end else begin
          meta_117_valid_0 <= _GEN_7445;
        end
      end else begin
        meta_117_valid_0 <= _GEN_2170;
      end
    end else begin
      meta_117_valid_0 <= _GEN_2170;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_117_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_117_valid_1 <= _GEN_2682;
        end else begin
          meta_117_valid_1 <= _GEN_7446;
        end
      end else begin
        meta_117_valid_1 <= _GEN_2682;
      end
    end else begin
      meta_117_valid_1 <= _GEN_2682;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_117_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_117_lru <= _GEN_8353;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_118_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_118_valid_0 <= _GEN_2171;
        end else begin
          meta_118_valid_0 <= _GEN_7447;
        end
      end else begin
        meta_118_valid_0 <= _GEN_2171;
      end
    end else begin
      meta_118_valid_0 <= _GEN_2171;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_118_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_118_valid_1 <= _GEN_2683;
        end else begin
          meta_118_valid_1 <= _GEN_7448;
        end
      end else begin
        meta_118_valid_1 <= _GEN_2683;
      end
    end else begin
      meta_118_valid_1 <= _GEN_2683;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_118_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_118_lru <= _GEN_8354;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_119_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_119_valid_0 <= _GEN_2172;
        end else begin
          meta_119_valid_0 <= _GEN_7449;
        end
      end else begin
        meta_119_valid_0 <= _GEN_2172;
      end
    end else begin
      meta_119_valid_0 <= _GEN_2172;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_119_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_119_valid_1 <= _GEN_2684;
        end else begin
          meta_119_valid_1 <= _GEN_7450;
        end
      end else begin
        meta_119_valid_1 <= _GEN_2684;
      end
    end else begin
      meta_119_valid_1 <= _GEN_2684;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_119_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_119_lru <= _GEN_8355;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_120_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_120_valid_0 <= _GEN_2173;
        end else begin
          meta_120_valid_0 <= _GEN_7451;
        end
      end else begin
        meta_120_valid_0 <= _GEN_2173;
      end
    end else begin
      meta_120_valid_0 <= _GEN_2173;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_120_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_120_valid_1 <= _GEN_2685;
        end else begin
          meta_120_valid_1 <= _GEN_7452;
        end
      end else begin
        meta_120_valid_1 <= _GEN_2685;
      end
    end else begin
      meta_120_valid_1 <= _GEN_2685;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_120_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_120_lru <= _GEN_8356;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_121_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_121_valid_0 <= _GEN_2174;
        end else begin
          meta_121_valid_0 <= _GEN_7453;
        end
      end else begin
        meta_121_valid_0 <= _GEN_2174;
      end
    end else begin
      meta_121_valid_0 <= _GEN_2174;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_121_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_121_valid_1 <= _GEN_2686;
        end else begin
          meta_121_valid_1 <= _GEN_7454;
        end
      end else begin
        meta_121_valid_1 <= _GEN_2686;
      end
    end else begin
      meta_121_valid_1 <= _GEN_2686;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_121_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_121_lru <= _GEN_8357;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_122_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_122_valid_0 <= _GEN_2175;
        end else begin
          meta_122_valid_0 <= _GEN_7455;
        end
      end else begin
        meta_122_valid_0 <= _GEN_2175;
      end
    end else begin
      meta_122_valid_0 <= _GEN_2175;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_122_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_122_valid_1 <= _GEN_2687;
        end else begin
          meta_122_valid_1 <= _GEN_7456;
        end
      end else begin
        meta_122_valid_1 <= _GEN_2687;
      end
    end else begin
      meta_122_valid_1 <= _GEN_2687;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_122_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_122_lru <= _GEN_8358;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_123_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_123_valid_0 <= _GEN_2176;
        end else begin
          meta_123_valid_0 <= _GEN_7457;
        end
      end else begin
        meta_123_valid_0 <= _GEN_2176;
      end
    end else begin
      meta_123_valid_0 <= _GEN_2176;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_123_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_123_valid_1 <= _GEN_2688;
        end else begin
          meta_123_valid_1 <= _GEN_7458;
        end
      end else begin
        meta_123_valid_1 <= _GEN_2688;
      end
    end else begin
      meta_123_valid_1 <= _GEN_2688;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_123_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_123_lru <= _GEN_8359;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_124_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_124_valid_0 <= _GEN_2177;
        end else begin
          meta_124_valid_0 <= _GEN_7459;
        end
      end else begin
        meta_124_valid_0 <= _GEN_2177;
      end
    end else begin
      meta_124_valid_0 <= _GEN_2177;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_124_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_124_valid_1 <= _GEN_2689;
        end else begin
          meta_124_valid_1 <= _GEN_7460;
        end
      end else begin
        meta_124_valid_1 <= _GEN_2689;
      end
    end else begin
      meta_124_valid_1 <= _GEN_2689;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_124_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_124_lru <= _GEN_8360;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_125_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_125_valid_0 <= _GEN_2178;
        end else begin
          meta_125_valid_0 <= _GEN_7461;
        end
      end else begin
        meta_125_valid_0 <= _GEN_2178;
      end
    end else begin
      meta_125_valid_0 <= _GEN_2178;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_125_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_125_valid_1 <= _GEN_2690;
        end else begin
          meta_125_valid_1 <= _GEN_7462;
        end
      end else begin
        meta_125_valid_1 <= _GEN_2690;
      end
    end else begin
      meta_125_valid_1 <= _GEN_2690;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_125_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_125_lru <= _GEN_8361;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_126_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_126_valid_0 <= _GEN_2179;
        end else begin
          meta_126_valid_0 <= _GEN_7463;
        end
      end else begin
        meta_126_valid_0 <= _GEN_2179;
      end
    end else begin
      meta_126_valid_0 <= _GEN_2179;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_126_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_126_valid_1 <= _GEN_2691;
        end else begin
          meta_126_valid_1 <= _GEN_7464;
        end
      end else begin
        meta_126_valid_1 <= _GEN_2691;
      end
    end else begin
      meta_126_valid_1 <= _GEN_2691;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_126_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_126_lru <= _GEN_8362;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_127_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_127_valid_0 <= _GEN_2180;
        end else begin
          meta_127_valid_0 <= _GEN_7465;
        end
      end else begin
        meta_127_valid_0 <= _GEN_2180;
      end
    end else begin
      meta_127_valid_0 <= _GEN_2180;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_127_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_127_valid_1 <= _GEN_2692;
        end else begin
          meta_127_valid_1 <= _GEN_7466;
        end
      end else begin
        meta_127_valid_1 <= _GEN_2692;
      end
    end else begin
      meta_127_valid_1 <= _GEN_2692;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_127_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_127_lru <= _GEN_8363;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_128_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_128_valid_0 <= _GEN_2181;
        end else begin
          meta_128_valid_0 <= _GEN_7467;
        end
      end else begin
        meta_128_valid_0 <= _GEN_2181;
      end
    end else begin
      meta_128_valid_0 <= _GEN_2181;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_128_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_128_valid_1 <= _GEN_2693;
        end else begin
          meta_128_valid_1 <= _GEN_7468;
        end
      end else begin
        meta_128_valid_1 <= _GEN_2693;
      end
    end else begin
      meta_128_valid_1 <= _GEN_2693;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_128_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_128_lru <= _GEN_8364;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_129_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_129_valid_0 <= _GEN_2182;
        end else begin
          meta_129_valid_0 <= _GEN_7469;
        end
      end else begin
        meta_129_valid_0 <= _GEN_2182;
      end
    end else begin
      meta_129_valid_0 <= _GEN_2182;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_129_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_129_valid_1 <= _GEN_2694;
        end else begin
          meta_129_valid_1 <= _GEN_7470;
        end
      end else begin
        meta_129_valid_1 <= _GEN_2694;
      end
    end else begin
      meta_129_valid_1 <= _GEN_2694;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_129_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_129_lru <= _GEN_8365;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_130_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_130_valid_0 <= _GEN_2183;
        end else begin
          meta_130_valid_0 <= _GEN_7471;
        end
      end else begin
        meta_130_valid_0 <= _GEN_2183;
      end
    end else begin
      meta_130_valid_0 <= _GEN_2183;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_130_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_130_valid_1 <= _GEN_2695;
        end else begin
          meta_130_valid_1 <= _GEN_7472;
        end
      end else begin
        meta_130_valid_1 <= _GEN_2695;
      end
    end else begin
      meta_130_valid_1 <= _GEN_2695;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_130_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_130_lru <= _GEN_8366;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_131_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_131_valid_0 <= _GEN_2184;
        end else begin
          meta_131_valid_0 <= _GEN_7473;
        end
      end else begin
        meta_131_valid_0 <= _GEN_2184;
      end
    end else begin
      meta_131_valid_0 <= _GEN_2184;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_131_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_131_valid_1 <= _GEN_2696;
        end else begin
          meta_131_valid_1 <= _GEN_7474;
        end
      end else begin
        meta_131_valid_1 <= _GEN_2696;
      end
    end else begin
      meta_131_valid_1 <= _GEN_2696;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_131_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_131_lru <= _GEN_8367;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_132_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_132_valid_0 <= _GEN_2185;
        end else begin
          meta_132_valid_0 <= _GEN_7475;
        end
      end else begin
        meta_132_valid_0 <= _GEN_2185;
      end
    end else begin
      meta_132_valid_0 <= _GEN_2185;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_132_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_132_valid_1 <= _GEN_2697;
        end else begin
          meta_132_valid_1 <= _GEN_7476;
        end
      end else begin
        meta_132_valid_1 <= _GEN_2697;
      end
    end else begin
      meta_132_valid_1 <= _GEN_2697;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_132_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_132_lru <= _GEN_8368;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_133_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_133_valid_0 <= _GEN_2186;
        end else begin
          meta_133_valid_0 <= _GEN_7477;
        end
      end else begin
        meta_133_valid_0 <= _GEN_2186;
      end
    end else begin
      meta_133_valid_0 <= _GEN_2186;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_133_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_133_valid_1 <= _GEN_2698;
        end else begin
          meta_133_valid_1 <= _GEN_7478;
        end
      end else begin
        meta_133_valid_1 <= _GEN_2698;
      end
    end else begin
      meta_133_valid_1 <= _GEN_2698;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_133_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_133_lru <= _GEN_8369;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_134_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_134_valid_0 <= _GEN_2187;
        end else begin
          meta_134_valid_0 <= _GEN_7479;
        end
      end else begin
        meta_134_valid_0 <= _GEN_2187;
      end
    end else begin
      meta_134_valid_0 <= _GEN_2187;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_134_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_134_valid_1 <= _GEN_2699;
        end else begin
          meta_134_valid_1 <= _GEN_7480;
        end
      end else begin
        meta_134_valid_1 <= _GEN_2699;
      end
    end else begin
      meta_134_valid_1 <= _GEN_2699;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_134_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_134_lru <= _GEN_8370;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_135_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_135_valid_0 <= _GEN_2188;
        end else begin
          meta_135_valid_0 <= _GEN_7481;
        end
      end else begin
        meta_135_valid_0 <= _GEN_2188;
      end
    end else begin
      meta_135_valid_0 <= _GEN_2188;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_135_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_135_valid_1 <= _GEN_2700;
        end else begin
          meta_135_valid_1 <= _GEN_7482;
        end
      end else begin
        meta_135_valid_1 <= _GEN_2700;
      end
    end else begin
      meta_135_valid_1 <= _GEN_2700;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_135_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_135_lru <= _GEN_8371;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_136_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_136_valid_0 <= _GEN_2189;
        end else begin
          meta_136_valid_0 <= _GEN_7483;
        end
      end else begin
        meta_136_valid_0 <= _GEN_2189;
      end
    end else begin
      meta_136_valid_0 <= _GEN_2189;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_136_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_136_valid_1 <= _GEN_2701;
        end else begin
          meta_136_valid_1 <= _GEN_7484;
        end
      end else begin
        meta_136_valid_1 <= _GEN_2701;
      end
    end else begin
      meta_136_valid_1 <= _GEN_2701;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_136_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_136_lru <= _GEN_8372;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_137_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_137_valid_0 <= _GEN_2190;
        end else begin
          meta_137_valid_0 <= _GEN_7485;
        end
      end else begin
        meta_137_valid_0 <= _GEN_2190;
      end
    end else begin
      meta_137_valid_0 <= _GEN_2190;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_137_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_137_valid_1 <= _GEN_2702;
        end else begin
          meta_137_valid_1 <= _GEN_7486;
        end
      end else begin
        meta_137_valid_1 <= _GEN_2702;
      end
    end else begin
      meta_137_valid_1 <= _GEN_2702;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_137_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_137_lru <= _GEN_8373;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_138_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_138_valid_0 <= _GEN_2191;
        end else begin
          meta_138_valid_0 <= _GEN_7487;
        end
      end else begin
        meta_138_valid_0 <= _GEN_2191;
      end
    end else begin
      meta_138_valid_0 <= _GEN_2191;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_138_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_138_valid_1 <= _GEN_2703;
        end else begin
          meta_138_valid_1 <= _GEN_7488;
        end
      end else begin
        meta_138_valid_1 <= _GEN_2703;
      end
    end else begin
      meta_138_valid_1 <= _GEN_2703;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_138_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_138_lru <= _GEN_8374;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_139_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_139_valid_0 <= _GEN_2192;
        end else begin
          meta_139_valid_0 <= _GEN_7489;
        end
      end else begin
        meta_139_valid_0 <= _GEN_2192;
      end
    end else begin
      meta_139_valid_0 <= _GEN_2192;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_139_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_139_valid_1 <= _GEN_2704;
        end else begin
          meta_139_valid_1 <= _GEN_7490;
        end
      end else begin
        meta_139_valid_1 <= _GEN_2704;
      end
    end else begin
      meta_139_valid_1 <= _GEN_2704;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_139_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_139_lru <= _GEN_8375;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_140_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_140_valid_0 <= _GEN_2193;
        end else begin
          meta_140_valid_0 <= _GEN_7491;
        end
      end else begin
        meta_140_valid_0 <= _GEN_2193;
      end
    end else begin
      meta_140_valid_0 <= _GEN_2193;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_140_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_140_valid_1 <= _GEN_2705;
        end else begin
          meta_140_valid_1 <= _GEN_7492;
        end
      end else begin
        meta_140_valid_1 <= _GEN_2705;
      end
    end else begin
      meta_140_valid_1 <= _GEN_2705;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_140_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_140_lru <= _GEN_8376;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_141_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_141_valid_0 <= _GEN_2194;
        end else begin
          meta_141_valid_0 <= _GEN_7493;
        end
      end else begin
        meta_141_valid_0 <= _GEN_2194;
      end
    end else begin
      meta_141_valid_0 <= _GEN_2194;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_141_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_141_valid_1 <= _GEN_2706;
        end else begin
          meta_141_valid_1 <= _GEN_7494;
        end
      end else begin
        meta_141_valid_1 <= _GEN_2706;
      end
    end else begin
      meta_141_valid_1 <= _GEN_2706;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_141_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_141_lru <= _GEN_8377;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_142_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_142_valid_0 <= _GEN_2195;
        end else begin
          meta_142_valid_0 <= _GEN_7495;
        end
      end else begin
        meta_142_valid_0 <= _GEN_2195;
      end
    end else begin
      meta_142_valid_0 <= _GEN_2195;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_142_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_142_valid_1 <= _GEN_2707;
        end else begin
          meta_142_valid_1 <= _GEN_7496;
        end
      end else begin
        meta_142_valid_1 <= _GEN_2707;
      end
    end else begin
      meta_142_valid_1 <= _GEN_2707;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_142_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_142_lru <= _GEN_8378;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_143_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_143_valid_0 <= _GEN_2196;
        end else begin
          meta_143_valid_0 <= _GEN_7497;
        end
      end else begin
        meta_143_valid_0 <= _GEN_2196;
      end
    end else begin
      meta_143_valid_0 <= _GEN_2196;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_143_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_143_valid_1 <= _GEN_2708;
        end else begin
          meta_143_valid_1 <= _GEN_7498;
        end
      end else begin
        meta_143_valid_1 <= _GEN_2708;
      end
    end else begin
      meta_143_valid_1 <= _GEN_2708;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_143_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_143_lru <= _GEN_8379;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_144_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_144_valid_0 <= _GEN_2197;
        end else begin
          meta_144_valid_0 <= _GEN_7499;
        end
      end else begin
        meta_144_valid_0 <= _GEN_2197;
      end
    end else begin
      meta_144_valid_0 <= _GEN_2197;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_144_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_144_valid_1 <= _GEN_2709;
        end else begin
          meta_144_valid_1 <= _GEN_7500;
        end
      end else begin
        meta_144_valid_1 <= _GEN_2709;
      end
    end else begin
      meta_144_valid_1 <= _GEN_2709;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_144_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_144_lru <= _GEN_8380;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_145_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_145_valid_0 <= _GEN_2198;
        end else begin
          meta_145_valid_0 <= _GEN_7501;
        end
      end else begin
        meta_145_valid_0 <= _GEN_2198;
      end
    end else begin
      meta_145_valid_0 <= _GEN_2198;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_145_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_145_valid_1 <= _GEN_2710;
        end else begin
          meta_145_valid_1 <= _GEN_7502;
        end
      end else begin
        meta_145_valid_1 <= _GEN_2710;
      end
    end else begin
      meta_145_valid_1 <= _GEN_2710;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_145_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_145_lru <= _GEN_8381;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_146_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_146_valid_0 <= _GEN_2199;
        end else begin
          meta_146_valid_0 <= _GEN_7503;
        end
      end else begin
        meta_146_valid_0 <= _GEN_2199;
      end
    end else begin
      meta_146_valid_0 <= _GEN_2199;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_146_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_146_valid_1 <= _GEN_2711;
        end else begin
          meta_146_valid_1 <= _GEN_7504;
        end
      end else begin
        meta_146_valid_1 <= _GEN_2711;
      end
    end else begin
      meta_146_valid_1 <= _GEN_2711;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_146_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_146_lru <= _GEN_8382;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_147_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_147_valid_0 <= _GEN_2200;
        end else begin
          meta_147_valid_0 <= _GEN_7505;
        end
      end else begin
        meta_147_valid_0 <= _GEN_2200;
      end
    end else begin
      meta_147_valid_0 <= _GEN_2200;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_147_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_147_valid_1 <= _GEN_2712;
        end else begin
          meta_147_valid_1 <= _GEN_7506;
        end
      end else begin
        meta_147_valid_1 <= _GEN_2712;
      end
    end else begin
      meta_147_valid_1 <= _GEN_2712;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_147_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_147_lru <= _GEN_8383;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_148_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_148_valid_0 <= _GEN_2201;
        end else begin
          meta_148_valid_0 <= _GEN_7507;
        end
      end else begin
        meta_148_valid_0 <= _GEN_2201;
      end
    end else begin
      meta_148_valid_0 <= _GEN_2201;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_148_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_148_valid_1 <= _GEN_2713;
        end else begin
          meta_148_valid_1 <= _GEN_7508;
        end
      end else begin
        meta_148_valid_1 <= _GEN_2713;
      end
    end else begin
      meta_148_valid_1 <= _GEN_2713;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_148_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_148_lru <= _GEN_8384;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_149_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_149_valid_0 <= _GEN_2202;
        end else begin
          meta_149_valid_0 <= _GEN_7509;
        end
      end else begin
        meta_149_valid_0 <= _GEN_2202;
      end
    end else begin
      meta_149_valid_0 <= _GEN_2202;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_149_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_149_valid_1 <= _GEN_2714;
        end else begin
          meta_149_valid_1 <= _GEN_7510;
        end
      end else begin
        meta_149_valid_1 <= _GEN_2714;
      end
    end else begin
      meta_149_valid_1 <= _GEN_2714;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_149_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_149_lru <= _GEN_8385;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_150_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_150_valid_0 <= _GEN_2203;
        end else begin
          meta_150_valid_0 <= _GEN_7511;
        end
      end else begin
        meta_150_valid_0 <= _GEN_2203;
      end
    end else begin
      meta_150_valid_0 <= _GEN_2203;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_150_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_150_valid_1 <= _GEN_2715;
        end else begin
          meta_150_valid_1 <= _GEN_7512;
        end
      end else begin
        meta_150_valid_1 <= _GEN_2715;
      end
    end else begin
      meta_150_valid_1 <= _GEN_2715;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_150_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_150_lru <= _GEN_8386;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_151_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_151_valid_0 <= _GEN_2204;
        end else begin
          meta_151_valid_0 <= _GEN_7513;
        end
      end else begin
        meta_151_valid_0 <= _GEN_2204;
      end
    end else begin
      meta_151_valid_0 <= _GEN_2204;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_151_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_151_valid_1 <= _GEN_2716;
        end else begin
          meta_151_valid_1 <= _GEN_7514;
        end
      end else begin
        meta_151_valid_1 <= _GEN_2716;
      end
    end else begin
      meta_151_valid_1 <= _GEN_2716;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_151_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_151_lru <= _GEN_8387;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_152_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_152_valid_0 <= _GEN_2205;
        end else begin
          meta_152_valid_0 <= _GEN_7515;
        end
      end else begin
        meta_152_valid_0 <= _GEN_2205;
      end
    end else begin
      meta_152_valid_0 <= _GEN_2205;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_152_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_152_valid_1 <= _GEN_2717;
        end else begin
          meta_152_valid_1 <= _GEN_7516;
        end
      end else begin
        meta_152_valid_1 <= _GEN_2717;
      end
    end else begin
      meta_152_valid_1 <= _GEN_2717;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_152_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_152_lru <= _GEN_8388;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_153_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_153_valid_0 <= _GEN_2206;
        end else begin
          meta_153_valid_0 <= _GEN_7517;
        end
      end else begin
        meta_153_valid_0 <= _GEN_2206;
      end
    end else begin
      meta_153_valid_0 <= _GEN_2206;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_153_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_153_valid_1 <= _GEN_2718;
        end else begin
          meta_153_valid_1 <= _GEN_7518;
        end
      end else begin
        meta_153_valid_1 <= _GEN_2718;
      end
    end else begin
      meta_153_valid_1 <= _GEN_2718;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_153_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_153_lru <= _GEN_8389;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_154_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_154_valid_0 <= _GEN_2207;
        end else begin
          meta_154_valid_0 <= _GEN_7519;
        end
      end else begin
        meta_154_valid_0 <= _GEN_2207;
      end
    end else begin
      meta_154_valid_0 <= _GEN_2207;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_154_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_154_valid_1 <= _GEN_2719;
        end else begin
          meta_154_valid_1 <= _GEN_7520;
        end
      end else begin
        meta_154_valid_1 <= _GEN_2719;
      end
    end else begin
      meta_154_valid_1 <= _GEN_2719;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_154_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_154_lru <= _GEN_8390;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_155_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_155_valid_0 <= _GEN_2208;
        end else begin
          meta_155_valid_0 <= _GEN_7521;
        end
      end else begin
        meta_155_valid_0 <= _GEN_2208;
      end
    end else begin
      meta_155_valid_0 <= _GEN_2208;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_155_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_155_valid_1 <= _GEN_2720;
        end else begin
          meta_155_valid_1 <= _GEN_7522;
        end
      end else begin
        meta_155_valid_1 <= _GEN_2720;
      end
    end else begin
      meta_155_valid_1 <= _GEN_2720;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_155_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_155_lru <= _GEN_8391;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_156_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_156_valid_0 <= _GEN_2209;
        end else begin
          meta_156_valid_0 <= _GEN_7523;
        end
      end else begin
        meta_156_valid_0 <= _GEN_2209;
      end
    end else begin
      meta_156_valid_0 <= _GEN_2209;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_156_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_156_valid_1 <= _GEN_2721;
        end else begin
          meta_156_valid_1 <= _GEN_7524;
        end
      end else begin
        meta_156_valid_1 <= _GEN_2721;
      end
    end else begin
      meta_156_valid_1 <= _GEN_2721;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_156_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_156_lru <= _GEN_8392;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_157_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_157_valid_0 <= _GEN_2210;
        end else begin
          meta_157_valid_0 <= _GEN_7525;
        end
      end else begin
        meta_157_valid_0 <= _GEN_2210;
      end
    end else begin
      meta_157_valid_0 <= _GEN_2210;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_157_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_157_valid_1 <= _GEN_2722;
        end else begin
          meta_157_valid_1 <= _GEN_7526;
        end
      end else begin
        meta_157_valid_1 <= _GEN_2722;
      end
    end else begin
      meta_157_valid_1 <= _GEN_2722;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_157_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_157_lru <= _GEN_8393;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_158_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_158_valid_0 <= _GEN_2211;
        end else begin
          meta_158_valid_0 <= _GEN_7527;
        end
      end else begin
        meta_158_valid_0 <= _GEN_2211;
      end
    end else begin
      meta_158_valid_0 <= _GEN_2211;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_158_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_158_valid_1 <= _GEN_2723;
        end else begin
          meta_158_valid_1 <= _GEN_7528;
        end
      end else begin
        meta_158_valid_1 <= _GEN_2723;
      end
    end else begin
      meta_158_valid_1 <= _GEN_2723;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_158_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_158_lru <= _GEN_8394;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_159_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_159_valid_0 <= _GEN_2212;
        end else begin
          meta_159_valid_0 <= _GEN_7529;
        end
      end else begin
        meta_159_valid_0 <= _GEN_2212;
      end
    end else begin
      meta_159_valid_0 <= _GEN_2212;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_159_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_159_valid_1 <= _GEN_2724;
        end else begin
          meta_159_valid_1 <= _GEN_7530;
        end
      end else begin
        meta_159_valid_1 <= _GEN_2724;
      end
    end else begin
      meta_159_valid_1 <= _GEN_2724;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_159_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_159_lru <= _GEN_8395;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_160_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_160_valid_0 <= _GEN_2213;
        end else begin
          meta_160_valid_0 <= _GEN_7531;
        end
      end else begin
        meta_160_valid_0 <= _GEN_2213;
      end
    end else begin
      meta_160_valid_0 <= _GEN_2213;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_160_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_160_valid_1 <= _GEN_2725;
        end else begin
          meta_160_valid_1 <= _GEN_7532;
        end
      end else begin
        meta_160_valid_1 <= _GEN_2725;
      end
    end else begin
      meta_160_valid_1 <= _GEN_2725;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_160_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_160_lru <= _GEN_8396;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_161_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_161_valid_0 <= _GEN_2214;
        end else begin
          meta_161_valid_0 <= _GEN_7533;
        end
      end else begin
        meta_161_valid_0 <= _GEN_2214;
      end
    end else begin
      meta_161_valid_0 <= _GEN_2214;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_161_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_161_valid_1 <= _GEN_2726;
        end else begin
          meta_161_valid_1 <= _GEN_7534;
        end
      end else begin
        meta_161_valid_1 <= _GEN_2726;
      end
    end else begin
      meta_161_valid_1 <= _GEN_2726;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_161_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_161_lru <= _GEN_8397;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_162_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_162_valid_0 <= _GEN_2215;
        end else begin
          meta_162_valid_0 <= _GEN_7535;
        end
      end else begin
        meta_162_valid_0 <= _GEN_2215;
      end
    end else begin
      meta_162_valid_0 <= _GEN_2215;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_162_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_162_valid_1 <= _GEN_2727;
        end else begin
          meta_162_valid_1 <= _GEN_7536;
        end
      end else begin
        meta_162_valid_1 <= _GEN_2727;
      end
    end else begin
      meta_162_valid_1 <= _GEN_2727;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_162_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_162_lru <= _GEN_8398;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_163_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_163_valid_0 <= _GEN_2216;
        end else begin
          meta_163_valid_0 <= _GEN_7537;
        end
      end else begin
        meta_163_valid_0 <= _GEN_2216;
      end
    end else begin
      meta_163_valid_0 <= _GEN_2216;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_163_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_163_valid_1 <= _GEN_2728;
        end else begin
          meta_163_valid_1 <= _GEN_7538;
        end
      end else begin
        meta_163_valid_1 <= _GEN_2728;
      end
    end else begin
      meta_163_valid_1 <= _GEN_2728;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_163_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_163_lru <= _GEN_8399;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_164_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_164_valid_0 <= _GEN_2217;
        end else begin
          meta_164_valid_0 <= _GEN_7539;
        end
      end else begin
        meta_164_valid_0 <= _GEN_2217;
      end
    end else begin
      meta_164_valid_0 <= _GEN_2217;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_164_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_164_valid_1 <= _GEN_2729;
        end else begin
          meta_164_valid_1 <= _GEN_7540;
        end
      end else begin
        meta_164_valid_1 <= _GEN_2729;
      end
    end else begin
      meta_164_valid_1 <= _GEN_2729;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_164_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_164_lru <= _GEN_8400;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_165_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_165_valid_0 <= _GEN_2218;
        end else begin
          meta_165_valid_0 <= _GEN_7541;
        end
      end else begin
        meta_165_valid_0 <= _GEN_2218;
      end
    end else begin
      meta_165_valid_0 <= _GEN_2218;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_165_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_165_valid_1 <= _GEN_2730;
        end else begin
          meta_165_valid_1 <= _GEN_7542;
        end
      end else begin
        meta_165_valid_1 <= _GEN_2730;
      end
    end else begin
      meta_165_valid_1 <= _GEN_2730;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_165_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_165_lru <= _GEN_8401;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_166_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_166_valid_0 <= _GEN_2219;
        end else begin
          meta_166_valid_0 <= _GEN_7543;
        end
      end else begin
        meta_166_valid_0 <= _GEN_2219;
      end
    end else begin
      meta_166_valid_0 <= _GEN_2219;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_166_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_166_valid_1 <= _GEN_2731;
        end else begin
          meta_166_valid_1 <= _GEN_7544;
        end
      end else begin
        meta_166_valid_1 <= _GEN_2731;
      end
    end else begin
      meta_166_valid_1 <= _GEN_2731;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_166_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_166_lru <= _GEN_8402;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_167_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_167_valid_0 <= _GEN_2220;
        end else begin
          meta_167_valid_0 <= _GEN_7545;
        end
      end else begin
        meta_167_valid_0 <= _GEN_2220;
      end
    end else begin
      meta_167_valid_0 <= _GEN_2220;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_167_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_167_valid_1 <= _GEN_2732;
        end else begin
          meta_167_valid_1 <= _GEN_7546;
        end
      end else begin
        meta_167_valid_1 <= _GEN_2732;
      end
    end else begin
      meta_167_valid_1 <= _GEN_2732;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_167_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_167_lru <= _GEN_8403;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_168_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_168_valid_0 <= _GEN_2221;
        end else begin
          meta_168_valid_0 <= _GEN_7547;
        end
      end else begin
        meta_168_valid_0 <= _GEN_2221;
      end
    end else begin
      meta_168_valid_0 <= _GEN_2221;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_168_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_168_valid_1 <= _GEN_2733;
        end else begin
          meta_168_valid_1 <= _GEN_7548;
        end
      end else begin
        meta_168_valid_1 <= _GEN_2733;
      end
    end else begin
      meta_168_valid_1 <= _GEN_2733;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_168_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_168_lru <= _GEN_8404;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_169_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_169_valid_0 <= _GEN_2222;
        end else begin
          meta_169_valid_0 <= _GEN_7549;
        end
      end else begin
        meta_169_valid_0 <= _GEN_2222;
      end
    end else begin
      meta_169_valid_0 <= _GEN_2222;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_169_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_169_valid_1 <= _GEN_2734;
        end else begin
          meta_169_valid_1 <= _GEN_7550;
        end
      end else begin
        meta_169_valid_1 <= _GEN_2734;
      end
    end else begin
      meta_169_valid_1 <= _GEN_2734;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_169_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_169_lru <= _GEN_8405;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_170_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_170_valid_0 <= _GEN_2223;
        end else begin
          meta_170_valid_0 <= _GEN_7551;
        end
      end else begin
        meta_170_valid_0 <= _GEN_2223;
      end
    end else begin
      meta_170_valid_0 <= _GEN_2223;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_170_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_170_valid_1 <= _GEN_2735;
        end else begin
          meta_170_valid_1 <= _GEN_7552;
        end
      end else begin
        meta_170_valid_1 <= _GEN_2735;
      end
    end else begin
      meta_170_valid_1 <= _GEN_2735;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_170_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_170_lru <= _GEN_8406;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_171_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_171_valid_0 <= _GEN_2224;
        end else begin
          meta_171_valid_0 <= _GEN_7553;
        end
      end else begin
        meta_171_valid_0 <= _GEN_2224;
      end
    end else begin
      meta_171_valid_0 <= _GEN_2224;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_171_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_171_valid_1 <= _GEN_2736;
        end else begin
          meta_171_valid_1 <= _GEN_7554;
        end
      end else begin
        meta_171_valid_1 <= _GEN_2736;
      end
    end else begin
      meta_171_valid_1 <= _GEN_2736;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_171_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_171_lru <= _GEN_8407;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_172_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_172_valid_0 <= _GEN_2225;
        end else begin
          meta_172_valid_0 <= _GEN_7555;
        end
      end else begin
        meta_172_valid_0 <= _GEN_2225;
      end
    end else begin
      meta_172_valid_0 <= _GEN_2225;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_172_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_172_valid_1 <= _GEN_2737;
        end else begin
          meta_172_valid_1 <= _GEN_7556;
        end
      end else begin
        meta_172_valid_1 <= _GEN_2737;
      end
    end else begin
      meta_172_valid_1 <= _GEN_2737;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_172_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_172_lru <= _GEN_8408;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_173_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_173_valid_0 <= _GEN_2226;
        end else begin
          meta_173_valid_0 <= _GEN_7557;
        end
      end else begin
        meta_173_valid_0 <= _GEN_2226;
      end
    end else begin
      meta_173_valid_0 <= _GEN_2226;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_173_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_173_valid_1 <= _GEN_2738;
        end else begin
          meta_173_valid_1 <= _GEN_7558;
        end
      end else begin
        meta_173_valid_1 <= _GEN_2738;
      end
    end else begin
      meta_173_valid_1 <= _GEN_2738;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_173_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_173_lru <= _GEN_8409;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_174_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_174_valid_0 <= _GEN_2227;
        end else begin
          meta_174_valid_0 <= _GEN_7559;
        end
      end else begin
        meta_174_valid_0 <= _GEN_2227;
      end
    end else begin
      meta_174_valid_0 <= _GEN_2227;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_174_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_174_valid_1 <= _GEN_2739;
        end else begin
          meta_174_valid_1 <= _GEN_7560;
        end
      end else begin
        meta_174_valid_1 <= _GEN_2739;
      end
    end else begin
      meta_174_valid_1 <= _GEN_2739;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_174_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_174_lru <= _GEN_8410;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_175_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_175_valid_0 <= _GEN_2228;
        end else begin
          meta_175_valid_0 <= _GEN_7561;
        end
      end else begin
        meta_175_valid_0 <= _GEN_2228;
      end
    end else begin
      meta_175_valid_0 <= _GEN_2228;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_175_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_175_valid_1 <= _GEN_2740;
        end else begin
          meta_175_valid_1 <= _GEN_7562;
        end
      end else begin
        meta_175_valid_1 <= _GEN_2740;
      end
    end else begin
      meta_175_valid_1 <= _GEN_2740;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_175_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_175_lru <= _GEN_8411;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_176_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_176_valid_0 <= _GEN_2229;
        end else begin
          meta_176_valid_0 <= _GEN_7563;
        end
      end else begin
        meta_176_valid_0 <= _GEN_2229;
      end
    end else begin
      meta_176_valid_0 <= _GEN_2229;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_176_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_176_valid_1 <= _GEN_2741;
        end else begin
          meta_176_valid_1 <= _GEN_7564;
        end
      end else begin
        meta_176_valid_1 <= _GEN_2741;
      end
    end else begin
      meta_176_valid_1 <= _GEN_2741;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_176_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_176_lru <= _GEN_8412;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_177_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_177_valid_0 <= _GEN_2230;
        end else begin
          meta_177_valid_0 <= _GEN_7565;
        end
      end else begin
        meta_177_valid_0 <= _GEN_2230;
      end
    end else begin
      meta_177_valid_0 <= _GEN_2230;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_177_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_177_valid_1 <= _GEN_2742;
        end else begin
          meta_177_valid_1 <= _GEN_7566;
        end
      end else begin
        meta_177_valid_1 <= _GEN_2742;
      end
    end else begin
      meta_177_valid_1 <= _GEN_2742;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_177_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_177_lru <= _GEN_8413;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_178_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_178_valid_0 <= _GEN_2231;
        end else begin
          meta_178_valid_0 <= _GEN_7567;
        end
      end else begin
        meta_178_valid_0 <= _GEN_2231;
      end
    end else begin
      meta_178_valid_0 <= _GEN_2231;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_178_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_178_valid_1 <= _GEN_2743;
        end else begin
          meta_178_valid_1 <= _GEN_7568;
        end
      end else begin
        meta_178_valid_1 <= _GEN_2743;
      end
    end else begin
      meta_178_valid_1 <= _GEN_2743;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_178_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_178_lru <= _GEN_8414;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_179_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_179_valid_0 <= _GEN_2232;
        end else begin
          meta_179_valid_0 <= _GEN_7569;
        end
      end else begin
        meta_179_valid_0 <= _GEN_2232;
      end
    end else begin
      meta_179_valid_0 <= _GEN_2232;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_179_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_179_valid_1 <= _GEN_2744;
        end else begin
          meta_179_valid_1 <= _GEN_7570;
        end
      end else begin
        meta_179_valid_1 <= _GEN_2744;
      end
    end else begin
      meta_179_valid_1 <= _GEN_2744;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_179_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_179_lru <= _GEN_8415;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_180_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_180_valid_0 <= _GEN_2233;
        end else begin
          meta_180_valid_0 <= _GEN_7571;
        end
      end else begin
        meta_180_valid_0 <= _GEN_2233;
      end
    end else begin
      meta_180_valid_0 <= _GEN_2233;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_180_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_180_valid_1 <= _GEN_2745;
        end else begin
          meta_180_valid_1 <= _GEN_7572;
        end
      end else begin
        meta_180_valid_1 <= _GEN_2745;
      end
    end else begin
      meta_180_valid_1 <= _GEN_2745;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_180_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_180_lru <= _GEN_8416;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_181_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_181_valid_0 <= _GEN_2234;
        end else begin
          meta_181_valid_0 <= _GEN_7573;
        end
      end else begin
        meta_181_valid_0 <= _GEN_2234;
      end
    end else begin
      meta_181_valid_0 <= _GEN_2234;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_181_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_181_valid_1 <= _GEN_2746;
        end else begin
          meta_181_valid_1 <= _GEN_7574;
        end
      end else begin
        meta_181_valid_1 <= _GEN_2746;
      end
    end else begin
      meta_181_valid_1 <= _GEN_2746;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_181_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_181_lru <= _GEN_8417;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_182_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_182_valid_0 <= _GEN_2235;
        end else begin
          meta_182_valid_0 <= _GEN_7575;
        end
      end else begin
        meta_182_valid_0 <= _GEN_2235;
      end
    end else begin
      meta_182_valid_0 <= _GEN_2235;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_182_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_182_valid_1 <= _GEN_2747;
        end else begin
          meta_182_valid_1 <= _GEN_7576;
        end
      end else begin
        meta_182_valid_1 <= _GEN_2747;
      end
    end else begin
      meta_182_valid_1 <= _GEN_2747;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_182_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_182_lru <= _GEN_8418;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_183_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_183_valid_0 <= _GEN_2236;
        end else begin
          meta_183_valid_0 <= _GEN_7577;
        end
      end else begin
        meta_183_valid_0 <= _GEN_2236;
      end
    end else begin
      meta_183_valid_0 <= _GEN_2236;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_183_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_183_valid_1 <= _GEN_2748;
        end else begin
          meta_183_valid_1 <= _GEN_7578;
        end
      end else begin
        meta_183_valid_1 <= _GEN_2748;
      end
    end else begin
      meta_183_valid_1 <= _GEN_2748;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_183_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_183_lru <= _GEN_8419;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_184_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_184_valid_0 <= _GEN_2237;
        end else begin
          meta_184_valid_0 <= _GEN_7579;
        end
      end else begin
        meta_184_valid_0 <= _GEN_2237;
      end
    end else begin
      meta_184_valid_0 <= _GEN_2237;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_184_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_184_valid_1 <= _GEN_2749;
        end else begin
          meta_184_valid_1 <= _GEN_7580;
        end
      end else begin
        meta_184_valid_1 <= _GEN_2749;
      end
    end else begin
      meta_184_valid_1 <= _GEN_2749;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_184_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_184_lru <= _GEN_8420;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_185_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_185_valid_0 <= _GEN_2238;
        end else begin
          meta_185_valid_0 <= _GEN_7581;
        end
      end else begin
        meta_185_valid_0 <= _GEN_2238;
      end
    end else begin
      meta_185_valid_0 <= _GEN_2238;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_185_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_185_valid_1 <= _GEN_2750;
        end else begin
          meta_185_valid_1 <= _GEN_7582;
        end
      end else begin
        meta_185_valid_1 <= _GEN_2750;
      end
    end else begin
      meta_185_valid_1 <= _GEN_2750;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_185_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_185_lru <= _GEN_8421;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_186_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_186_valid_0 <= _GEN_2239;
        end else begin
          meta_186_valid_0 <= _GEN_7583;
        end
      end else begin
        meta_186_valid_0 <= _GEN_2239;
      end
    end else begin
      meta_186_valid_0 <= _GEN_2239;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_186_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_186_valid_1 <= _GEN_2751;
        end else begin
          meta_186_valid_1 <= _GEN_7584;
        end
      end else begin
        meta_186_valid_1 <= _GEN_2751;
      end
    end else begin
      meta_186_valid_1 <= _GEN_2751;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_186_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_186_lru <= _GEN_8422;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_187_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_187_valid_0 <= _GEN_2240;
        end else begin
          meta_187_valid_0 <= _GEN_7585;
        end
      end else begin
        meta_187_valid_0 <= _GEN_2240;
      end
    end else begin
      meta_187_valid_0 <= _GEN_2240;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_187_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_187_valid_1 <= _GEN_2752;
        end else begin
          meta_187_valid_1 <= _GEN_7586;
        end
      end else begin
        meta_187_valid_1 <= _GEN_2752;
      end
    end else begin
      meta_187_valid_1 <= _GEN_2752;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_187_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_187_lru <= _GEN_8423;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_188_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_188_valid_0 <= _GEN_2241;
        end else begin
          meta_188_valid_0 <= _GEN_7587;
        end
      end else begin
        meta_188_valid_0 <= _GEN_2241;
      end
    end else begin
      meta_188_valid_0 <= _GEN_2241;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_188_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_188_valid_1 <= _GEN_2753;
        end else begin
          meta_188_valid_1 <= _GEN_7588;
        end
      end else begin
        meta_188_valid_1 <= _GEN_2753;
      end
    end else begin
      meta_188_valid_1 <= _GEN_2753;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_188_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_188_lru <= _GEN_8424;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_189_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_189_valid_0 <= _GEN_2242;
        end else begin
          meta_189_valid_0 <= _GEN_7589;
        end
      end else begin
        meta_189_valid_0 <= _GEN_2242;
      end
    end else begin
      meta_189_valid_0 <= _GEN_2242;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_189_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_189_valid_1 <= _GEN_2754;
        end else begin
          meta_189_valid_1 <= _GEN_7590;
        end
      end else begin
        meta_189_valid_1 <= _GEN_2754;
      end
    end else begin
      meta_189_valid_1 <= _GEN_2754;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_189_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_189_lru <= _GEN_8425;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_190_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_190_valid_0 <= _GEN_2243;
        end else begin
          meta_190_valid_0 <= _GEN_7591;
        end
      end else begin
        meta_190_valid_0 <= _GEN_2243;
      end
    end else begin
      meta_190_valid_0 <= _GEN_2243;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_190_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_190_valid_1 <= _GEN_2755;
        end else begin
          meta_190_valid_1 <= _GEN_7592;
        end
      end else begin
        meta_190_valid_1 <= _GEN_2755;
      end
    end else begin
      meta_190_valid_1 <= _GEN_2755;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_190_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_190_lru <= _GEN_8426;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_191_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_191_valid_0 <= _GEN_2244;
        end else begin
          meta_191_valid_0 <= _GEN_7593;
        end
      end else begin
        meta_191_valid_0 <= _GEN_2244;
      end
    end else begin
      meta_191_valid_0 <= _GEN_2244;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_191_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_191_valid_1 <= _GEN_2756;
        end else begin
          meta_191_valid_1 <= _GEN_7594;
        end
      end else begin
        meta_191_valid_1 <= _GEN_2756;
      end
    end else begin
      meta_191_valid_1 <= _GEN_2756;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_191_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_191_lru <= _GEN_8427;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_192_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_192_valid_0 <= _GEN_2245;
        end else begin
          meta_192_valid_0 <= _GEN_7595;
        end
      end else begin
        meta_192_valid_0 <= _GEN_2245;
      end
    end else begin
      meta_192_valid_0 <= _GEN_2245;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_192_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_192_valid_1 <= _GEN_2757;
        end else begin
          meta_192_valid_1 <= _GEN_7596;
        end
      end else begin
        meta_192_valid_1 <= _GEN_2757;
      end
    end else begin
      meta_192_valid_1 <= _GEN_2757;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_192_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_192_lru <= _GEN_8428;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_193_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_193_valid_0 <= _GEN_2246;
        end else begin
          meta_193_valid_0 <= _GEN_7597;
        end
      end else begin
        meta_193_valid_0 <= _GEN_2246;
      end
    end else begin
      meta_193_valid_0 <= _GEN_2246;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_193_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_193_valid_1 <= _GEN_2758;
        end else begin
          meta_193_valid_1 <= _GEN_7598;
        end
      end else begin
        meta_193_valid_1 <= _GEN_2758;
      end
    end else begin
      meta_193_valid_1 <= _GEN_2758;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_193_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_193_lru <= _GEN_8429;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_194_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_194_valid_0 <= _GEN_2247;
        end else begin
          meta_194_valid_0 <= _GEN_7599;
        end
      end else begin
        meta_194_valid_0 <= _GEN_2247;
      end
    end else begin
      meta_194_valid_0 <= _GEN_2247;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_194_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_194_valid_1 <= _GEN_2759;
        end else begin
          meta_194_valid_1 <= _GEN_7600;
        end
      end else begin
        meta_194_valid_1 <= _GEN_2759;
      end
    end else begin
      meta_194_valid_1 <= _GEN_2759;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_194_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_194_lru <= _GEN_8430;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_195_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_195_valid_0 <= _GEN_2248;
        end else begin
          meta_195_valid_0 <= _GEN_7601;
        end
      end else begin
        meta_195_valid_0 <= _GEN_2248;
      end
    end else begin
      meta_195_valid_0 <= _GEN_2248;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_195_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_195_valid_1 <= _GEN_2760;
        end else begin
          meta_195_valid_1 <= _GEN_7602;
        end
      end else begin
        meta_195_valid_1 <= _GEN_2760;
      end
    end else begin
      meta_195_valid_1 <= _GEN_2760;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_195_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_195_lru <= _GEN_8431;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_196_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_196_valid_0 <= _GEN_2249;
        end else begin
          meta_196_valid_0 <= _GEN_7603;
        end
      end else begin
        meta_196_valid_0 <= _GEN_2249;
      end
    end else begin
      meta_196_valid_0 <= _GEN_2249;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_196_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_196_valid_1 <= _GEN_2761;
        end else begin
          meta_196_valid_1 <= _GEN_7604;
        end
      end else begin
        meta_196_valid_1 <= _GEN_2761;
      end
    end else begin
      meta_196_valid_1 <= _GEN_2761;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_196_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_196_lru <= _GEN_8432;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_197_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_197_valid_0 <= _GEN_2250;
        end else begin
          meta_197_valid_0 <= _GEN_7605;
        end
      end else begin
        meta_197_valid_0 <= _GEN_2250;
      end
    end else begin
      meta_197_valid_0 <= _GEN_2250;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_197_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_197_valid_1 <= _GEN_2762;
        end else begin
          meta_197_valid_1 <= _GEN_7606;
        end
      end else begin
        meta_197_valid_1 <= _GEN_2762;
      end
    end else begin
      meta_197_valid_1 <= _GEN_2762;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_197_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_197_lru <= _GEN_8433;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_198_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_198_valid_0 <= _GEN_2251;
        end else begin
          meta_198_valid_0 <= _GEN_7607;
        end
      end else begin
        meta_198_valid_0 <= _GEN_2251;
      end
    end else begin
      meta_198_valid_0 <= _GEN_2251;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_198_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_198_valid_1 <= _GEN_2763;
        end else begin
          meta_198_valid_1 <= _GEN_7608;
        end
      end else begin
        meta_198_valid_1 <= _GEN_2763;
      end
    end else begin
      meta_198_valid_1 <= _GEN_2763;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_198_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_198_lru <= _GEN_8434;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_199_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_199_valid_0 <= _GEN_2252;
        end else begin
          meta_199_valid_0 <= _GEN_7609;
        end
      end else begin
        meta_199_valid_0 <= _GEN_2252;
      end
    end else begin
      meta_199_valid_0 <= _GEN_2252;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_199_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_199_valid_1 <= _GEN_2764;
        end else begin
          meta_199_valid_1 <= _GEN_7610;
        end
      end else begin
        meta_199_valid_1 <= _GEN_2764;
      end
    end else begin
      meta_199_valid_1 <= _GEN_2764;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_199_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_199_lru <= _GEN_8435;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_200_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_200_valid_0 <= _GEN_2253;
        end else begin
          meta_200_valid_0 <= _GEN_7611;
        end
      end else begin
        meta_200_valid_0 <= _GEN_2253;
      end
    end else begin
      meta_200_valid_0 <= _GEN_2253;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_200_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_200_valid_1 <= _GEN_2765;
        end else begin
          meta_200_valid_1 <= _GEN_7612;
        end
      end else begin
        meta_200_valid_1 <= _GEN_2765;
      end
    end else begin
      meta_200_valid_1 <= _GEN_2765;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_200_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_200_lru <= _GEN_8436;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_201_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_201_valid_0 <= _GEN_2254;
        end else begin
          meta_201_valid_0 <= _GEN_7613;
        end
      end else begin
        meta_201_valid_0 <= _GEN_2254;
      end
    end else begin
      meta_201_valid_0 <= _GEN_2254;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_201_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_201_valid_1 <= _GEN_2766;
        end else begin
          meta_201_valid_1 <= _GEN_7614;
        end
      end else begin
        meta_201_valid_1 <= _GEN_2766;
      end
    end else begin
      meta_201_valid_1 <= _GEN_2766;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_201_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_201_lru <= _GEN_8437;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_202_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_202_valid_0 <= _GEN_2255;
        end else begin
          meta_202_valid_0 <= _GEN_7615;
        end
      end else begin
        meta_202_valid_0 <= _GEN_2255;
      end
    end else begin
      meta_202_valid_0 <= _GEN_2255;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_202_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_202_valid_1 <= _GEN_2767;
        end else begin
          meta_202_valid_1 <= _GEN_7616;
        end
      end else begin
        meta_202_valid_1 <= _GEN_2767;
      end
    end else begin
      meta_202_valid_1 <= _GEN_2767;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_202_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_202_lru <= _GEN_8438;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_203_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_203_valid_0 <= _GEN_2256;
        end else begin
          meta_203_valid_0 <= _GEN_7617;
        end
      end else begin
        meta_203_valid_0 <= _GEN_2256;
      end
    end else begin
      meta_203_valid_0 <= _GEN_2256;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_203_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_203_valid_1 <= _GEN_2768;
        end else begin
          meta_203_valid_1 <= _GEN_7618;
        end
      end else begin
        meta_203_valid_1 <= _GEN_2768;
      end
    end else begin
      meta_203_valid_1 <= _GEN_2768;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_203_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_203_lru <= _GEN_8439;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_204_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_204_valid_0 <= _GEN_2257;
        end else begin
          meta_204_valid_0 <= _GEN_7619;
        end
      end else begin
        meta_204_valid_0 <= _GEN_2257;
      end
    end else begin
      meta_204_valid_0 <= _GEN_2257;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_204_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_204_valid_1 <= _GEN_2769;
        end else begin
          meta_204_valid_1 <= _GEN_7620;
        end
      end else begin
        meta_204_valid_1 <= _GEN_2769;
      end
    end else begin
      meta_204_valid_1 <= _GEN_2769;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_204_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_204_lru <= _GEN_8440;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_205_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_205_valid_0 <= _GEN_2258;
        end else begin
          meta_205_valid_0 <= _GEN_7621;
        end
      end else begin
        meta_205_valid_0 <= _GEN_2258;
      end
    end else begin
      meta_205_valid_0 <= _GEN_2258;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_205_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_205_valid_1 <= _GEN_2770;
        end else begin
          meta_205_valid_1 <= _GEN_7622;
        end
      end else begin
        meta_205_valid_1 <= _GEN_2770;
      end
    end else begin
      meta_205_valid_1 <= _GEN_2770;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_205_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_205_lru <= _GEN_8441;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_206_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_206_valid_0 <= _GEN_2259;
        end else begin
          meta_206_valid_0 <= _GEN_7623;
        end
      end else begin
        meta_206_valid_0 <= _GEN_2259;
      end
    end else begin
      meta_206_valid_0 <= _GEN_2259;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_206_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_206_valid_1 <= _GEN_2771;
        end else begin
          meta_206_valid_1 <= _GEN_7624;
        end
      end else begin
        meta_206_valid_1 <= _GEN_2771;
      end
    end else begin
      meta_206_valid_1 <= _GEN_2771;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_206_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_206_lru <= _GEN_8442;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_207_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_207_valid_0 <= _GEN_2260;
        end else begin
          meta_207_valid_0 <= _GEN_7625;
        end
      end else begin
        meta_207_valid_0 <= _GEN_2260;
      end
    end else begin
      meta_207_valid_0 <= _GEN_2260;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_207_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_207_valid_1 <= _GEN_2772;
        end else begin
          meta_207_valid_1 <= _GEN_7626;
        end
      end else begin
        meta_207_valid_1 <= _GEN_2772;
      end
    end else begin
      meta_207_valid_1 <= _GEN_2772;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_207_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_207_lru <= _GEN_8443;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_208_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_208_valid_0 <= _GEN_2261;
        end else begin
          meta_208_valid_0 <= _GEN_7627;
        end
      end else begin
        meta_208_valid_0 <= _GEN_2261;
      end
    end else begin
      meta_208_valid_0 <= _GEN_2261;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_208_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_208_valid_1 <= _GEN_2773;
        end else begin
          meta_208_valid_1 <= _GEN_7628;
        end
      end else begin
        meta_208_valid_1 <= _GEN_2773;
      end
    end else begin
      meta_208_valid_1 <= _GEN_2773;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_208_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_208_lru <= _GEN_8444;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_209_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_209_valid_0 <= _GEN_2262;
        end else begin
          meta_209_valid_0 <= _GEN_7629;
        end
      end else begin
        meta_209_valid_0 <= _GEN_2262;
      end
    end else begin
      meta_209_valid_0 <= _GEN_2262;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_209_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_209_valid_1 <= _GEN_2774;
        end else begin
          meta_209_valid_1 <= _GEN_7630;
        end
      end else begin
        meta_209_valid_1 <= _GEN_2774;
      end
    end else begin
      meta_209_valid_1 <= _GEN_2774;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_209_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_209_lru <= _GEN_8445;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_210_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_210_valid_0 <= _GEN_2263;
        end else begin
          meta_210_valid_0 <= _GEN_7631;
        end
      end else begin
        meta_210_valid_0 <= _GEN_2263;
      end
    end else begin
      meta_210_valid_0 <= _GEN_2263;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_210_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_210_valid_1 <= _GEN_2775;
        end else begin
          meta_210_valid_1 <= _GEN_7632;
        end
      end else begin
        meta_210_valid_1 <= _GEN_2775;
      end
    end else begin
      meta_210_valid_1 <= _GEN_2775;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_210_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_210_lru <= _GEN_8446;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_211_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_211_valid_0 <= _GEN_2264;
        end else begin
          meta_211_valid_0 <= _GEN_7633;
        end
      end else begin
        meta_211_valid_0 <= _GEN_2264;
      end
    end else begin
      meta_211_valid_0 <= _GEN_2264;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_211_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_211_valid_1 <= _GEN_2776;
        end else begin
          meta_211_valid_1 <= _GEN_7634;
        end
      end else begin
        meta_211_valid_1 <= _GEN_2776;
      end
    end else begin
      meta_211_valid_1 <= _GEN_2776;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_211_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_211_lru <= _GEN_8447;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_212_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_212_valid_0 <= _GEN_2265;
        end else begin
          meta_212_valid_0 <= _GEN_7635;
        end
      end else begin
        meta_212_valid_0 <= _GEN_2265;
      end
    end else begin
      meta_212_valid_0 <= _GEN_2265;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_212_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_212_valid_1 <= _GEN_2777;
        end else begin
          meta_212_valid_1 <= _GEN_7636;
        end
      end else begin
        meta_212_valid_1 <= _GEN_2777;
      end
    end else begin
      meta_212_valid_1 <= _GEN_2777;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_212_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_212_lru <= _GEN_8448;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_213_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_213_valid_0 <= _GEN_2266;
        end else begin
          meta_213_valid_0 <= _GEN_7637;
        end
      end else begin
        meta_213_valid_0 <= _GEN_2266;
      end
    end else begin
      meta_213_valid_0 <= _GEN_2266;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_213_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_213_valid_1 <= _GEN_2778;
        end else begin
          meta_213_valid_1 <= _GEN_7638;
        end
      end else begin
        meta_213_valid_1 <= _GEN_2778;
      end
    end else begin
      meta_213_valid_1 <= _GEN_2778;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_213_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_213_lru <= _GEN_8449;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_214_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_214_valid_0 <= _GEN_2267;
        end else begin
          meta_214_valid_0 <= _GEN_7639;
        end
      end else begin
        meta_214_valid_0 <= _GEN_2267;
      end
    end else begin
      meta_214_valid_0 <= _GEN_2267;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_214_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_214_valid_1 <= _GEN_2779;
        end else begin
          meta_214_valid_1 <= _GEN_7640;
        end
      end else begin
        meta_214_valid_1 <= _GEN_2779;
      end
    end else begin
      meta_214_valid_1 <= _GEN_2779;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_214_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_214_lru <= _GEN_8450;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_215_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_215_valid_0 <= _GEN_2268;
        end else begin
          meta_215_valid_0 <= _GEN_7641;
        end
      end else begin
        meta_215_valid_0 <= _GEN_2268;
      end
    end else begin
      meta_215_valid_0 <= _GEN_2268;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_215_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_215_valid_1 <= _GEN_2780;
        end else begin
          meta_215_valid_1 <= _GEN_7642;
        end
      end else begin
        meta_215_valid_1 <= _GEN_2780;
      end
    end else begin
      meta_215_valid_1 <= _GEN_2780;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_215_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_215_lru <= _GEN_8451;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_216_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_216_valid_0 <= _GEN_2269;
        end else begin
          meta_216_valid_0 <= _GEN_7643;
        end
      end else begin
        meta_216_valid_0 <= _GEN_2269;
      end
    end else begin
      meta_216_valid_0 <= _GEN_2269;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_216_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_216_valid_1 <= _GEN_2781;
        end else begin
          meta_216_valid_1 <= _GEN_7644;
        end
      end else begin
        meta_216_valid_1 <= _GEN_2781;
      end
    end else begin
      meta_216_valid_1 <= _GEN_2781;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_216_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_216_lru <= _GEN_8452;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_217_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_217_valid_0 <= _GEN_2270;
        end else begin
          meta_217_valid_0 <= _GEN_7645;
        end
      end else begin
        meta_217_valid_0 <= _GEN_2270;
      end
    end else begin
      meta_217_valid_0 <= _GEN_2270;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_217_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_217_valid_1 <= _GEN_2782;
        end else begin
          meta_217_valid_1 <= _GEN_7646;
        end
      end else begin
        meta_217_valid_1 <= _GEN_2782;
      end
    end else begin
      meta_217_valid_1 <= _GEN_2782;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_217_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_217_lru <= _GEN_8453;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_218_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_218_valid_0 <= _GEN_2271;
        end else begin
          meta_218_valid_0 <= _GEN_7647;
        end
      end else begin
        meta_218_valid_0 <= _GEN_2271;
      end
    end else begin
      meta_218_valid_0 <= _GEN_2271;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_218_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_218_valid_1 <= _GEN_2783;
        end else begin
          meta_218_valid_1 <= _GEN_7648;
        end
      end else begin
        meta_218_valid_1 <= _GEN_2783;
      end
    end else begin
      meta_218_valid_1 <= _GEN_2783;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_218_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_218_lru <= _GEN_8454;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_219_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_219_valid_0 <= _GEN_2272;
        end else begin
          meta_219_valid_0 <= _GEN_7649;
        end
      end else begin
        meta_219_valid_0 <= _GEN_2272;
      end
    end else begin
      meta_219_valid_0 <= _GEN_2272;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_219_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_219_valid_1 <= _GEN_2784;
        end else begin
          meta_219_valid_1 <= _GEN_7650;
        end
      end else begin
        meta_219_valid_1 <= _GEN_2784;
      end
    end else begin
      meta_219_valid_1 <= _GEN_2784;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_219_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_219_lru <= _GEN_8455;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_220_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_220_valid_0 <= _GEN_2273;
        end else begin
          meta_220_valid_0 <= _GEN_7651;
        end
      end else begin
        meta_220_valid_0 <= _GEN_2273;
      end
    end else begin
      meta_220_valid_0 <= _GEN_2273;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_220_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_220_valid_1 <= _GEN_2785;
        end else begin
          meta_220_valid_1 <= _GEN_7652;
        end
      end else begin
        meta_220_valid_1 <= _GEN_2785;
      end
    end else begin
      meta_220_valid_1 <= _GEN_2785;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_220_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_220_lru <= _GEN_8456;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_221_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_221_valid_0 <= _GEN_2274;
        end else begin
          meta_221_valid_0 <= _GEN_7653;
        end
      end else begin
        meta_221_valid_0 <= _GEN_2274;
      end
    end else begin
      meta_221_valid_0 <= _GEN_2274;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_221_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_221_valid_1 <= _GEN_2786;
        end else begin
          meta_221_valid_1 <= _GEN_7654;
        end
      end else begin
        meta_221_valid_1 <= _GEN_2786;
      end
    end else begin
      meta_221_valid_1 <= _GEN_2786;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_221_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_221_lru <= _GEN_8457;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_222_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_222_valid_0 <= _GEN_2275;
        end else begin
          meta_222_valid_0 <= _GEN_7655;
        end
      end else begin
        meta_222_valid_0 <= _GEN_2275;
      end
    end else begin
      meta_222_valid_0 <= _GEN_2275;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_222_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_222_valid_1 <= _GEN_2787;
        end else begin
          meta_222_valid_1 <= _GEN_7656;
        end
      end else begin
        meta_222_valid_1 <= _GEN_2787;
      end
    end else begin
      meta_222_valid_1 <= _GEN_2787;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_222_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_222_lru <= _GEN_8458;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_223_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_223_valid_0 <= _GEN_2276;
        end else begin
          meta_223_valid_0 <= _GEN_7657;
        end
      end else begin
        meta_223_valid_0 <= _GEN_2276;
      end
    end else begin
      meta_223_valid_0 <= _GEN_2276;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_223_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_223_valid_1 <= _GEN_2788;
        end else begin
          meta_223_valid_1 <= _GEN_7658;
        end
      end else begin
        meta_223_valid_1 <= _GEN_2788;
      end
    end else begin
      meta_223_valid_1 <= _GEN_2788;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_223_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_223_lru <= _GEN_8459;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_224_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_224_valid_0 <= _GEN_2277;
        end else begin
          meta_224_valid_0 <= _GEN_7659;
        end
      end else begin
        meta_224_valid_0 <= _GEN_2277;
      end
    end else begin
      meta_224_valid_0 <= _GEN_2277;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_224_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_224_valid_1 <= _GEN_2789;
        end else begin
          meta_224_valid_1 <= _GEN_7660;
        end
      end else begin
        meta_224_valid_1 <= _GEN_2789;
      end
    end else begin
      meta_224_valid_1 <= _GEN_2789;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_224_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_224_lru <= _GEN_8460;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_225_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_225_valid_0 <= _GEN_2278;
        end else begin
          meta_225_valid_0 <= _GEN_7661;
        end
      end else begin
        meta_225_valid_0 <= _GEN_2278;
      end
    end else begin
      meta_225_valid_0 <= _GEN_2278;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_225_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_225_valid_1 <= _GEN_2790;
        end else begin
          meta_225_valid_1 <= _GEN_7662;
        end
      end else begin
        meta_225_valid_1 <= _GEN_2790;
      end
    end else begin
      meta_225_valid_1 <= _GEN_2790;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_225_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_225_lru <= _GEN_8461;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_226_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_226_valid_0 <= _GEN_2279;
        end else begin
          meta_226_valid_0 <= _GEN_7663;
        end
      end else begin
        meta_226_valid_0 <= _GEN_2279;
      end
    end else begin
      meta_226_valid_0 <= _GEN_2279;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_226_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_226_valid_1 <= _GEN_2791;
        end else begin
          meta_226_valid_1 <= _GEN_7664;
        end
      end else begin
        meta_226_valid_1 <= _GEN_2791;
      end
    end else begin
      meta_226_valid_1 <= _GEN_2791;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_226_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_226_lru <= _GEN_8462;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_227_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_227_valid_0 <= _GEN_2280;
        end else begin
          meta_227_valid_0 <= _GEN_7665;
        end
      end else begin
        meta_227_valid_0 <= _GEN_2280;
      end
    end else begin
      meta_227_valid_0 <= _GEN_2280;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_227_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_227_valid_1 <= _GEN_2792;
        end else begin
          meta_227_valid_1 <= _GEN_7666;
        end
      end else begin
        meta_227_valid_1 <= _GEN_2792;
      end
    end else begin
      meta_227_valid_1 <= _GEN_2792;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_227_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_227_lru <= _GEN_8463;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_228_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_228_valid_0 <= _GEN_2281;
        end else begin
          meta_228_valid_0 <= _GEN_7667;
        end
      end else begin
        meta_228_valid_0 <= _GEN_2281;
      end
    end else begin
      meta_228_valid_0 <= _GEN_2281;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_228_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_228_valid_1 <= _GEN_2793;
        end else begin
          meta_228_valid_1 <= _GEN_7668;
        end
      end else begin
        meta_228_valid_1 <= _GEN_2793;
      end
    end else begin
      meta_228_valid_1 <= _GEN_2793;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_228_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_228_lru <= _GEN_8464;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_229_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_229_valid_0 <= _GEN_2282;
        end else begin
          meta_229_valid_0 <= _GEN_7669;
        end
      end else begin
        meta_229_valid_0 <= _GEN_2282;
      end
    end else begin
      meta_229_valid_0 <= _GEN_2282;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_229_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_229_valid_1 <= _GEN_2794;
        end else begin
          meta_229_valid_1 <= _GEN_7670;
        end
      end else begin
        meta_229_valid_1 <= _GEN_2794;
      end
    end else begin
      meta_229_valid_1 <= _GEN_2794;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_229_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_229_lru <= _GEN_8465;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_230_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_230_valid_0 <= _GEN_2283;
        end else begin
          meta_230_valid_0 <= _GEN_7671;
        end
      end else begin
        meta_230_valid_0 <= _GEN_2283;
      end
    end else begin
      meta_230_valid_0 <= _GEN_2283;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_230_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_230_valid_1 <= _GEN_2795;
        end else begin
          meta_230_valid_1 <= _GEN_7672;
        end
      end else begin
        meta_230_valid_1 <= _GEN_2795;
      end
    end else begin
      meta_230_valid_1 <= _GEN_2795;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_230_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_230_lru <= _GEN_8466;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_231_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_231_valid_0 <= _GEN_2284;
        end else begin
          meta_231_valid_0 <= _GEN_7673;
        end
      end else begin
        meta_231_valid_0 <= _GEN_2284;
      end
    end else begin
      meta_231_valid_0 <= _GEN_2284;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_231_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_231_valid_1 <= _GEN_2796;
        end else begin
          meta_231_valid_1 <= _GEN_7674;
        end
      end else begin
        meta_231_valid_1 <= _GEN_2796;
      end
    end else begin
      meta_231_valid_1 <= _GEN_2796;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_231_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_231_lru <= _GEN_8467;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_232_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_232_valid_0 <= _GEN_2285;
        end else begin
          meta_232_valid_0 <= _GEN_7675;
        end
      end else begin
        meta_232_valid_0 <= _GEN_2285;
      end
    end else begin
      meta_232_valid_0 <= _GEN_2285;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_232_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_232_valid_1 <= _GEN_2797;
        end else begin
          meta_232_valid_1 <= _GEN_7676;
        end
      end else begin
        meta_232_valid_1 <= _GEN_2797;
      end
    end else begin
      meta_232_valid_1 <= _GEN_2797;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_232_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_232_lru <= _GEN_8468;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_233_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_233_valid_0 <= _GEN_2286;
        end else begin
          meta_233_valid_0 <= _GEN_7677;
        end
      end else begin
        meta_233_valid_0 <= _GEN_2286;
      end
    end else begin
      meta_233_valid_0 <= _GEN_2286;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_233_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_233_valid_1 <= _GEN_2798;
        end else begin
          meta_233_valid_1 <= _GEN_7678;
        end
      end else begin
        meta_233_valid_1 <= _GEN_2798;
      end
    end else begin
      meta_233_valid_1 <= _GEN_2798;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_233_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_233_lru <= _GEN_8469;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_234_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_234_valid_0 <= _GEN_2287;
        end else begin
          meta_234_valid_0 <= _GEN_7679;
        end
      end else begin
        meta_234_valid_0 <= _GEN_2287;
      end
    end else begin
      meta_234_valid_0 <= _GEN_2287;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_234_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_234_valid_1 <= _GEN_2799;
        end else begin
          meta_234_valid_1 <= _GEN_7680;
        end
      end else begin
        meta_234_valid_1 <= _GEN_2799;
      end
    end else begin
      meta_234_valid_1 <= _GEN_2799;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_234_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_234_lru <= _GEN_8470;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_235_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_235_valid_0 <= _GEN_2288;
        end else begin
          meta_235_valid_0 <= _GEN_7681;
        end
      end else begin
        meta_235_valid_0 <= _GEN_2288;
      end
    end else begin
      meta_235_valid_0 <= _GEN_2288;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_235_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_235_valid_1 <= _GEN_2800;
        end else begin
          meta_235_valid_1 <= _GEN_7682;
        end
      end else begin
        meta_235_valid_1 <= _GEN_2800;
      end
    end else begin
      meta_235_valid_1 <= _GEN_2800;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_235_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_235_lru <= _GEN_8471;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_236_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_236_valid_0 <= _GEN_2289;
        end else begin
          meta_236_valid_0 <= _GEN_7683;
        end
      end else begin
        meta_236_valid_0 <= _GEN_2289;
      end
    end else begin
      meta_236_valid_0 <= _GEN_2289;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_236_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_236_valid_1 <= _GEN_2801;
        end else begin
          meta_236_valid_1 <= _GEN_7684;
        end
      end else begin
        meta_236_valid_1 <= _GEN_2801;
      end
    end else begin
      meta_236_valid_1 <= _GEN_2801;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_236_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_236_lru <= _GEN_8472;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_237_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_237_valid_0 <= _GEN_2290;
        end else begin
          meta_237_valid_0 <= _GEN_7685;
        end
      end else begin
        meta_237_valid_0 <= _GEN_2290;
      end
    end else begin
      meta_237_valid_0 <= _GEN_2290;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_237_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_237_valid_1 <= _GEN_2802;
        end else begin
          meta_237_valid_1 <= _GEN_7686;
        end
      end else begin
        meta_237_valid_1 <= _GEN_2802;
      end
    end else begin
      meta_237_valid_1 <= _GEN_2802;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_237_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_237_lru <= _GEN_8473;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_238_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_238_valid_0 <= _GEN_2291;
        end else begin
          meta_238_valid_0 <= _GEN_7687;
        end
      end else begin
        meta_238_valid_0 <= _GEN_2291;
      end
    end else begin
      meta_238_valid_0 <= _GEN_2291;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_238_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_238_valid_1 <= _GEN_2803;
        end else begin
          meta_238_valid_1 <= _GEN_7688;
        end
      end else begin
        meta_238_valid_1 <= _GEN_2803;
      end
    end else begin
      meta_238_valid_1 <= _GEN_2803;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_238_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_238_lru <= _GEN_8474;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_239_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_239_valid_0 <= _GEN_2292;
        end else begin
          meta_239_valid_0 <= _GEN_7689;
        end
      end else begin
        meta_239_valid_0 <= _GEN_2292;
      end
    end else begin
      meta_239_valid_0 <= _GEN_2292;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_239_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_239_valid_1 <= _GEN_2804;
        end else begin
          meta_239_valid_1 <= _GEN_7690;
        end
      end else begin
        meta_239_valid_1 <= _GEN_2804;
      end
    end else begin
      meta_239_valid_1 <= _GEN_2804;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_239_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_239_lru <= _GEN_8475;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_240_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_240_valid_0 <= _GEN_2293;
        end else begin
          meta_240_valid_0 <= _GEN_7691;
        end
      end else begin
        meta_240_valid_0 <= _GEN_2293;
      end
    end else begin
      meta_240_valid_0 <= _GEN_2293;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_240_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_240_valid_1 <= _GEN_2805;
        end else begin
          meta_240_valid_1 <= _GEN_7692;
        end
      end else begin
        meta_240_valid_1 <= _GEN_2805;
      end
    end else begin
      meta_240_valid_1 <= _GEN_2805;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_240_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_240_lru <= _GEN_8476;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_241_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_241_valid_0 <= _GEN_2294;
        end else begin
          meta_241_valid_0 <= _GEN_7693;
        end
      end else begin
        meta_241_valid_0 <= _GEN_2294;
      end
    end else begin
      meta_241_valid_0 <= _GEN_2294;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_241_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_241_valid_1 <= _GEN_2806;
        end else begin
          meta_241_valid_1 <= _GEN_7694;
        end
      end else begin
        meta_241_valid_1 <= _GEN_2806;
      end
    end else begin
      meta_241_valid_1 <= _GEN_2806;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_241_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_241_lru <= _GEN_8477;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_242_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_242_valid_0 <= _GEN_2295;
        end else begin
          meta_242_valid_0 <= _GEN_7695;
        end
      end else begin
        meta_242_valid_0 <= _GEN_2295;
      end
    end else begin
      meta_242_valid_0 <= _GEN_2295;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_242_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_242_valid_1 <= _GEN_2807;
        end else begin
          meta_242_valid_1 <= _GEN_7696;
        end
      end else begin
        meta_242_valid_1 <= _GEN_2807;
      end
    end else begin
      meta_242_valid_1 <= _GEN_2807;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_242_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_242_lru <= _GEN_8478;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_243_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_243_valid_0 <= _GEN_2296;
        end else begin
          meta_243_valid_0 <= _GEN_7697;
        end
      end else begin
        meta_243_valid_0 <= _GEN_2296;
      end
    end else begin
      meta_243_valid_0 <= _GEN_2296;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_243_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_243_valid_1 <= _GEN_2808;
        end else begin
          meta_243_valid_1 <= _GEN_7698;
        end
      end else begin
        meta_243_valid_1 <= _GEN_2808;
      end
    end else begin
      meta_243_valid_1 <= _GEN_2808;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_243_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_243_lru <= _GEN_8479;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_244_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_244_valid_0 <= _GEN_2297;
        end else begin
          meta_244_valid_0 <= _GEN_7699;
        end
      end else begin
        meta_244_valid_0 <= _GEN_2297;
      end
    end else begin
      meta_244_valid_0 <= _GEN_2297;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_244_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_244_valid_1 <= _GEN_2809;
        end else begin
          meta_244_valid_1 <= _GEN_7700;
        end
      end else begin
        meta_244_valid_1 <= _GEN_2809;
      end
    end else begin
      meta_244_valid_1 <= _GEN_2809;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_244_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_244_lru <= _GEN_8480;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_245_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_245_valid_0 <= _GEN_2298;
        end else begin
          meta_245_valid_0 <= _GEN_7701;
        end
      end else begin
        meta_245_valid_0 <= _GEN_2298;
      end
    end else begin
      meta_245_valid_0 <= _GEN_2298;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_245_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_245_valid_1 <= _GEN_2810;
        end else begin
          meta_245_valid_1 <= _GEN_7702;
        end
      end else begin
        meta_245_valid_1 <= _GEN_2810;
      end
    end else begin
      meta_245_valid_1 <= _GEN_2810;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_245_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_245_lru <= _GEN_8481;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_246_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_246_valid_0 <= _GEN_2299;
        end else begin
          meta_246_valid_0 <= _GEN_7703;
        end
      end else begin
        meta_246_valid_0 <= _GEN_2299;
      end
    end else begin
      meta_246_valid_0 <= _GEN_2299;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_246_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_246_valid_1 <= _GEN_2811;
        end else begin
          meta_246_valid_1 <= _GEN_7704;
        end
      end else begin
        meta_246_valid_1 <= _GEN_2811;
      end
    end else begin
      meta_246_valid_1 <= _GEN_2811;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_246_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_246_lru <= _GEN_8482;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_247_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_247_valid_0 <= _GEN_2300;
        end else begin
          meta_247_valid_0 <= _GEN_7705;
        end
      end else begin
        meta_247_valid_0 <= _GEN_2300;
      end
    end else begin
      meta_247_valid_0 <= _GEN_2300;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_247_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_247_valid_1 <= _GEN_2812;
        end else begin
          meta_247_valid_1 <= _GEN_7706;
        end
      end else begin
        meta_247_valid_1 <= _GEN_2812;
      end
    end else begin
      meta_247_valid_1 <= _GEN_2812;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_247_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_247_lru <= _GEN_8483;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_248_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_248_valid_0 <= _GEN_2301;
        end else begin
          meta_248_valid_0 <= _GEN_7707;
        end
      end else begin
        meta_248_valid_0 <= _GEN_2301;
      end
    end else begin
      meta_248_valid_0 <= _GEN_2301;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_248_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_248_valid_1 <= _GEN_2813;
        end else begin
          meta_248_valid_1 <= _GEN_7708;
        end
      end else begin
        meta_248_valid_1 <= _GEN_2813;
      end
    end else begin
      meta_248_valid_1 <= _GEN_2813;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_248_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_248_lru <= _GEN_8484;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_249_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_249_valid_0 <= _GEN_2302;
        end else begin
          meta_249_valid_0 <= _GEN_7709;
        end
      end else begin
        meta_249_valid_0 <= _GEN_2302;
      end
    end else begin
      meta_249_valid_0 <= _GEN_2302;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_249_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_249_valid_1 <= _GEN_2814;
        end else begin
          meta_249_valid_1 <= _GEN_7710;
        end
      end else begin
        meta_249_valid_1 <= _GEN_2814;
      end
    end else begin
      meta_249_valid_1 <= _GEN_2814;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_249_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_249_lru <= _GEN_8485;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_250_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_250_valid_0 <= _GEN_2303;
        end else begin
          meta_250_valid_0 <= _GEN_7711;
        end
      end else begin
        meta_250_valid_0 <= _GEN_2303;
      end
    end else begin
      meta_250_valid_0 <= _GEN_2303;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_250_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_250_valid_1 <= _GEN_2815;
        end else begin
          meta_250_valid_1 <= _GEN_7712;
        end
      end else begin
        meta_250_valid_1 <= _GEN_2815;
      end
    end else begin
      meta_250_valid_1 <= _GEN_2815;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_250_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_250_lru <= _GEN_8486;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_251_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_251_valid_0 <= _GEN_2304;
        end else begin
          meta_251_valid_0 <= _GEN_7713;
        end
      end else begin
        meta_251_valid_0 <= _GEN_2304;
      end
    end else begin
      meta_251_valid_0 <= _GEN_2304;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_251_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_251_valid_1 <= _GEN_2816;
        end else begin
          meta_251_valid_1 <= _GEN_7714;
        end
      end else begin
        meta_251_valid_1 <= _GEN_2816;
      end
    end else begin
      meta_251_valid_1 <= _GEN_2816;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_251_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_251_lru <= _GEN_8487;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_252_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_252_valid_0 <= _GEN_2305;
        end else begin
          meta_252_valid_0 <= _GEN_7715;
        end
      end else begin
        meta_252_valid_0 <= _GEN_2305;
      end
    end else begin
      meta_252_valid_0 <= _GEN_2305;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_252_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_252_valid_1 <= _GEN_2817;
        end else begin
          meta_252_valid_1 <= _GEN_7716;
        end
      end else begin
        meta_252_valid_1 <= _GEN_2817;
      end
    end else begin
      meta_252_valid_1 <= _GEN_2817;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_252_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_252_lru <= _GEN_8488;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_253_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_253_valid_0 <= _GEN_2306;
        end else begin
          meta_253_valid_0 <= _GEN_7717;
        end
      end else begin
        meta_253_valid_0 <= _GEN_2306;
      end
    end else begin
      meta_253_valid_0 <= _GEN_2306;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_253_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_253_valid_1 <= _GEN_2818;
        end else begin
          meta_253_valid_1 <= _GEN_7718;
        end
      end else begin
        meta_253_valid_1 <= _GEN_2818;
      end
    end else begin
      meta_253_valid_1 <= _GEN_2818;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_253_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_253_lru <= _GEN_8489;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_254_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_254_valid_0 <= _GEN_2307;
        end else begin
          meta_254_valid_0 <= _GEN_7719;
        end
      end else begin
        meta_254_valid_0 <= _GEN_2307;
      end
    end else begin
      meta_254_valid_0 <= _GEN_2307;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_254_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_254_valid_1 <= _GEN_2819;
        end else begin
          meta_254_valid_1 <= _GEN_7720;
        end
      end else begin
        meta_254_valid_1 <= _GEN_2819;
      end
    end else begin
      meta_254_valid_1 <= _GEN_2819;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_254_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_254_lru <= _GEN_8490;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_255_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_255_valid_0 <= _GEN_2308;
        end else begin
          meta_255_valid_0 <= _GEN_7721;
        end
      end else begin
        meta_255_valid_0 <= _GEN_2308;
      end
    end else begin
      meta_255_valid_0 <= _GEN_2308;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_255_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_255_valid_1 <= _GEN_2820;
        end else begin
          meta_255_valid_1 <= _GEN_7722;
        end
      end else begin
        meta_255_valid_1 <= _GEN_2820;
      end
    end else begin
      meta_255_valid_1 <= _GEN_2820;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_255_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_255_lru <= _GEN_8491;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_256_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_256_valid_0 <= _GEN_2309;
        end else begin
          meta_256_valid_0 <= _GEN_7723;
        end
      end else begin
        meta_256_valid_0 <= _GEN_2309;
      end
    end else begin
      meta_256_valid_0 <= _GEN_2309;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_256_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_256_valid_1 <= _GEN_2821;
        end else begin
          meta_256_valid_1 <= _GEN_7724;
        end
      end else begin
        meta_256_valid_1 <= _GEN_2821;
      end
    end else begin
      meta_256_valid_1 <= _GEN_2821;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_256_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_256_lru <= _GEN_8492;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_257_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_257_valid_0 <= _GEN_2310;
        end else begin
          meta_257_valid_0 <= _GEN_7725;
        end
      end else begin
        meta_257_valid_0 <= _GEN_2310;
      end
    end else begin
      meta_257_valid_0 <= _GEN_2310;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_257_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_257_valid_1 <= _GEN_2822;
        end else begin
          meta_257_valid_1 <= _GEN_7726;
        end
      end else begin
        meta_257_valid_1 <= _GEN_2822;
      end
    end else begin
      meta_257_valid_1 <= _GEN_2822;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_257_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_257_lru <= _GEN_8493;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_258_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_258_valid_0 <= _GEN_2311;
        end else begin
          meta_258_valid_0 <= _GEN_7727;
        end
      end else begin
        meta_258_valid_0 <= _GEN_2311;
      end
    end else begin
      meta_258_valid_0 <= _GEN_2311;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_258_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_258_valid_1 <= _GEN_2823;
        end else begin
          meta_258_valid_1 <= _GEN_7728;
        end
      end else begin
        meta_258_valid_1 <= _GEN_2823;
      end
    end else begin
      meta_258_valid_1 <= _GEN_2823;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_258_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_258_lru <= _GEN_8494;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_259_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_259_valid_0 <= _GEN_2312;
        end else begin
          meta_259_valid_0 <= _GEN_7729;
        end
      end else begin
        meta_259_valid_0 <= _GEN_2312;
      end
    end else begin
      meta_259_valid_0 <= _GEN_2312;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_259_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_259_valid_1 <= _GEN_2824;
        end else begin
          meta_259_valid_1 <= _GEN_7730;
        end
      end else begin
        meta_259_valid_1 <= _GEN_2824;
      end
    end else begin
      meta_259_valid_1 <= _GEN_2824;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_259_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_259_lru <= _GEN_8495;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_260_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_260_valid_0 <= _GEN_2313;
        end else begin
          meta_260_valid_0 <= _GEN_7731;
        end
      end else begin
        meta_260_valid_0 <= _GEN_2313;
      end
    end else begin
      meta_260_valid_0 <= _GEN_2313;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_260_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_260_valid_1 <= _GEN_2825;
        end else begin
          meta_260_valid_1 <= _GEN_7732;
        end
      end else begin
        meta_260_valid_1 <= _GEN_2825;
      end
    end else begin
      meta_260_valid_1 <= _GEN_2825;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_260_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_260_lru <= _GEN_8496;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_261_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_261_valid_0 <= _GEN_2314;
        end else begin
          meta_261_valid_0 <= _GEN_7733;
        end
      end else begin
        meta_261_valid_0 <= _GEN_2314;
      end
    end else begin
      meta_261_valid_0 <= _GEN_2314;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_261_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_261_valid_1 <= _GEN_2826;
        end else begin
          meta_261_valid_1 <= _GEN_7734;
        end
      end else begin
        meta_261_valid_1 <= _GEN_2826;
      end
    end else begin
      meta_261_valid_1 <= _GEN_2826;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_261_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_261_lru <= _GEN_8497;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_262_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_262_valid_0 <= _GEN_2315;
        end else begin
          meta_262_valid_0 <= _GEN_7735;
        end
      end else begin
        meta_262_valid_0 <= _GEN_2315;
      end
    end else begin
      meta_262_valid_0 <= _GEN_2315;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_262_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_262_valid_1 <= _GEN_2827;
        end else begin
          meta_262_valid_1 <= _GEN_7736;
        end
      end else begin
        meta_262_valid_1 <= _GEN_2827;
      end
    end else begin
      meta_262_valid_1 <= _GEN_2827;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_262_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_262_lru <= _GEN_8498;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_263_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_263_valid_0 <= _GEN_2316;
        end else begin
          meta_263_valid_0 <= _GEN_7737;
        end
      end else begin
        meta_263_valid_0 <= _GEN_2316;
      end
    end else begin
      meta_263_valid_0 <= _GEN_2316;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_263_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_263_valid_1 <= _GEN_2828;
        end else begin
          meta_263_valid_1 <= _GEN_7738;
        end
      end else begin
        meta_263_valid_1 <= _GEN_2828;
      end
    end else begin
      meta_263_valid_1 <= _GEN_2828;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_263_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_263_lru <= _GEN_8499;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_264_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_264_valid_0 <= _GEN_2317;
        end else begin
          meta_264_valid_0 <= _GEN_7739;
        end
      end else begin
        meta_264_valid_0 <= _GEN_2317;
      end
    end else begin
      meta_264_valid_0 <= _GEN_2317;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_264_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_264_valid_1 <= _GEN_2829;
        end else begin
          meta_264_valid_1 <= _GEN_7740;
        end
      end else begin
        meta_264_valid_1 <= _GEN_2829;
      end
    end else begin
      meta_264_valid_1 <= _GEN_2829;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_264_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_264_lru <= _GEN_8500;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_265_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_265_valid_0 <= _GEN_2318;
        end else begin
          meta_265_valid_0 <= _GEN_7741;
        end
      end else begin
        meta_265_valid_0 <= _GEN_2318;
      end
    end else begin
      meta_265_valid_0 <= _GEN_2318;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_265_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_265_valid_1 <= _GEN_2830;
        end else begin
          meta_265_valid_1 <= _GEN_7742;
        end
      end else begin
        meta_265_valid_1 <= _GEN_2830;
      end
    end else begin
      meta_265_valid_1 <= _GEN_2830;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_265_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_265_lru <= _GEN_8501;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_266_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_266_valid_0 <= _GEN_2319;
        end else begin
          meta_266_valid_0 <= _GEN_7743;
        end
      end else begin
        meta_266_valid_0 <= _GEN_2319;
      end
    end else begin
      meta_266_valid_0 <= _GEN_2319;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_266_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_266_valid_1 <= _GEN_2831;
        end else begin
          meta_266_valid_1 <= _GEN_7744;
        end
      end else begin
        meta_266_valid_1 <= _GEN_2831;
      end
    end else begin
      meta_266_valid_1 <= _GEN_2831;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_266_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_266_lru <= _GEN_8502;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_267_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_267_valid_0 <= _GEN_2320;
        end else begin
          meta_267_valid_0 <= _GEN_7745;
        end
      end else begin
        meta_267_valid_0 <= _GEN_2320;
      end
    end else begin
      meta_267_valid_0 <= _GEN_2320;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_267_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_267_valid_1 <= _GEN_2832;
        end else begin
          meta_267_valid_1 <= _GEN_7746;
        end
      end else begin
        meta_267_valid_1 <= _GEN_2832;
      end
    end else begin
      meta_267_valid_1 <= _GEN_2832;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_267_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_267_lru <= _GEN_8503;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_268_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_268_valid_0 <= _GEN_2321;
        end else begin
          meta_268_valid_0 <= _GEN_7747;
        end
      end else begin
        meta_268_valid_0 <= _GEN_2321;
      end
    end else begin
      meta_268_valid_0 <= _GEN_2321;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_268_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_268_valid_1 <= _GEN_2833;
        end else begin
          meta_268_valid_1 <= _GEN_7748;
        end
      end else begin
        meta_268_valid_1 <= _GEN_2833;
      end
    end else begin
      meta_268_valid_1 <= _GEN_2833;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_268_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_268_lru <= _GEN_8504;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_269_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_269_valid_0 <= _GEN_2322;
        end else begin
          meta_269_valid_0 <= _GEN_7749;
        end
      end else begin
        meta_269_valid_0 <= _GEN_2322;
      end
    end else begin
      meta_269_valid_0 <= _GEN_2322;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_269_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_269_valid_1 <= _GEN_2834;
        end else begin
          meta_269_valid_1 <= _GEN_7750;
        end
      end else begin
        meta_269_valid_1 <= _GEN_2834;
      end
    end else begin
      meta_269_valid_1 <= _GEN_2834;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_269_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_269_lru <= _GEN_8505;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_270_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_270_valid_0 <= _GEN_2323;
        end else begin
          meta_270_valid_0 <= _GEN_7751;
        end
      end else begin
        meta_270_valid_0 <= _GEN_2323;
      end
    end else begin
      meta_270_valid_0 <= _GEN_2323;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_270_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_270_valid_1 <= _GEN_2835;
        end else begin
          meta_270_valid_1 <= _GEN_7752;
        end
      end else begin
        meta_270_valid_1 <= _GEN_2835;
      end
    end else begin
      meta_270_valid_1 <= _GEN_2835;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_270_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_270_lru <= _GEN_8506;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_271_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_271_valid_0 <= _GEN_2324;
        end else begin
          meta_271_valid_0 <= _GEN_7753;
        end
      end else begin
        meta_271_valid_0 <= _GEN_2324;
      end
    end else begin
      meta_271_valid_0 <= _GEN_2324;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_271_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_271_valid_1 <= _GEN_2836;
        end else begin
          meta_271_valid_1 <= _GEN_7754;
        end
      end else begin
        meta_271_valid_1 <= _GEN_2836;
      end
    end else begin
      meta_271_valid_1 <= _GEN_2836;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_271_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_271_lru <= _GEN_8507;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_272_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_272_valid_0 <= _GEN_2325;
        end else begin
          meta_272_valid_0 <= _GEN_7755;
        end
      end else begin
        meta_272_valid_0 <= _GEN_2325;
      end
    end else begin
      meta_272_valid_0 <= _GEN_2325;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_272_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_272_valid_1 <= _GEN_2837;
        end else begin
          meta_272_valid_1 <= _GEN_7756;
        end
      end else begin
        meta_272_valid_1 <= _GEN_2837;
      end
    end else begin
      meta_272_valid_1 <= _GEN_2837;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_272_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_272_lru <= _GEN_8508;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_273_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_273_valid_0 <= _GEN_2326;
        end else begin
          meta_273_valid_0 <= _GEN_7757;
        end
      end else begin
        meta_273_valid_0 <= _GEN_2326;
      end
    end else begin
      meta_273_valid_0 <= _GEN_2326;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_273_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_273_valid_1 <= _GEN_2838;
        end else begin
          meta_273_valid_1 <= _GEN_7758;
        end
      end else begin
        meta_273_valid_1 <= _GEN_2838;
      end
    end else begin
      meta_273_valid_1 <= _GEN_2838;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_273_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_273_lru <= _GEN_8509;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_274_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_274_valid_0 <= _GEN_2327;
        end else begin
          meta_274_valid_0 <= _GEN_7759;
        end
      end else begin
        meta_274_valid_0 <= _GEN_2327;
      end
    end else begin
      meta_274_valid_0 <= _GEN_2327;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_274_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_274_valid_1 <= _GEN_2839;
        end else begin
          meta_274_valid_1 <= _GEN_7760;
        end
      end else begin
        meta_274_valid_1 <= _GEN_2839;
      end
    end else begin
      meta_274_valid_1 <= _GEN_2839;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_274_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_274_lru <= _GEN_8510;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_275_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_275_valid_0 <= _GEN_2328;
        end else begin
          meta_275_valid_0 <= _GEN_7761;
        end
      end else begin
        meta_275_valid_0 <= _GEN_2328;
      end
    end else begin
      meta_275_valid_0 <= _GEN_2328;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_275_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_275_valid_1 <= _GEN_2840;
        end else begin
          meta_275_valid_1 <= _GEN_7762;
        end
      end else begin
        meta_275_valid_1 <= _GEN_2840;
      end
    end else begin
      meta_275_valid_1 <= _GEN_2840;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_275_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_275_lru <= _GEN_8511;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_276_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_276_valid_0 <= _GEN_2329;
        end else begin
          meta_276_valid_0 <= _GEN_7763;
        end
      end else begin
        meta_276_valid_0 <= _GEN_2329;
      end
    end else begin
      meta_276_valid_0 <= _GEN_2329;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_276_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_276_valid_1 <= _GEN_2841;
        end else begin
          meta_276_valid_1 <= _GEN_7764;
        end
      end else begin
        meta_276_valid_1 <= _GEN_2841;
      end
    end else begin
      meta_276_valid_1 <= _GEN_2841;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_276_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_276_lru <= _GEN_8512;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_277_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_277_valid_0 <= _GEN_2330;
        end else begin
          meta_277_valid_0 <= _GEN_7765;
        end
      end else begin
        meta_277_valid_0 <= _GEN_2330;
      end
    end else begin
      meta_277_valid_0 <= _GEN_2330;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_277_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_277_valid_1 <= _GEN_2842;
        end else begin
          meta_277_valid_1 <= _GEN_7766;
        end
      end else begin
        meta_277_valid_1 <= _GEN_2842;
      end
    end else begin
      meta_277_valid_1 <= _GEN_2842;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_277_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_277_lru <= _GEN_8513;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_278_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_278_valid_0 <= _GEN_2331;
        end else begin
          meta_278_valid_0 <= _GEN_7767;
        end
      end else begin
        meta_278_valid_0 <= _GEN_2331;
      end
    end else begin
      meta_278_valid_0 <= _GEN_2331;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_278_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_278_valid_1 <= _GEN_2843;
        end else begin
          meta_278_valid_1 <= _GEN_7768;
        end
      end else begin
        meta_278_valid_1 <= _GEN_2843;
      end
    end else begin
      meta_278_valid_1 <= _GEN_2843;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_278_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_278_lru <= _GEN_8514;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_279_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_279_valid_0 <= _GEN_2332;
        end else begin
          meta_279_valid_0 <= _GEN_7769;
        end
      end else begin
        meta_279_valid_0 <= _GEN_2332;
      end
    end else begin
      meta_279_valid_0 <= _GEN_2332;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_279_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_279_valid_1 <= _GEN_2844;
        end else begin
          meta_279_valid_1 <= _GEN_7770;
        end
      end else begin
        meta_279_valid_1 <= _GEN_2844;
      end
    end else begin
      meta_279_valid_1 <= _GEN_2844;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_279_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_279_lru <= _GEN_8515;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_280_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_280_valid_0 <= _GEN_2333;
        end else begin
          meta_280_valid_0 <= _GEN_7771;
        end
      end else begin
        meta_280_valid_0 <= _GEN_2333;
      end
    end else begin
      meta_280_valid_0 <= _GEN_2333;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_280_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_280_valid_1 <= _GEN_2845;
        end else begin
          meta_280_valid_1 <= _GEN_7772;
        end
      end else begin
        meta_280_valid_1 <= _GEN_2845;
      end
    end else begin
      meta_280_valid_1 <= _GEN_2845;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_280_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_280_lru <= _GEN_8516;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_281_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_281_valid_0 <= _GEN_2334;
        end else begin
          meta_281_valid_0 <= _GEN_7773;
        end
      end else begin
        meta_281_valid_0 <= _GEN_2334;
      end
    end else begin
      meta_281_valid_0 <= _GEN_2334;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_281_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_281_valid_1 <= _GEN_2846;
        end else begin
          meta_281_valid_1 <= _GEN_7774;
        end
      end else begin
        meta_281_valid_1 <= _GEN_2846;
      end
    end else begin
      meta_281_valid_1 <= _GEN_2846;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_281_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_281_lru <= _GEN_8517;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_282_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_282_valid_0 <= _GEN_2335;
        end else begin
          meta_282_valid_0 <= _GEN_7775;
        end
      end else begin
        meta_282_valid_0 <= _GEN_2335;
      end
    end else begin
      meta_282_valid_0 <= _GEN_2335;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_282_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_282_valid_1 <= _GEN_2847;
        end else begin
          meta_282_valid_1 <= _GEN_7776;
        end
      end else begin
        meta_282_valid_1 <= _GEN_2847;
      end
    end else begin
      meta_282_valid_1 <= _GEN_2847;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_282_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_282_lru <= _GEN_8518;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_283_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_283_valid_0 <= _GEN_2336;
        end else begin
          meta_283_valid_0 <= _GEN_7777;
        end
      end else begin
        meta_283_valid_0 <= _GEN_2336;
      end
    end else begin
      meta_283_valid_0 <= _GEN_2336;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_283_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_283_valid_1 <= _GEN_2848;
        end else begin
          meta_283_valid_1 <= _GEN_7778;
        end
      end else begin
        meta_283_valid_1 <= _GEN_2848;
      end
    end else begin
      meta_283_valid_1 <= _GEN_2848;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_283_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_283_lru <= _GEN_8519;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_284_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_284_valid_0 <= _GEN_2337;
        end else begin
          meta_284_valid_0 <= _GEN_7779;
        end
      end else begin
        meta_284_valid_0 <= _GEN_2337;
      end
    end else begin
      meta_284_valid_0 <= _GEN_2337;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_284_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_284_valid_1 <= _GEN_2849;
        end else begin
          meta_284_valid_1 <= _GEN_7780;
        end
      end else begin
        meta_284_valid_1 <= _GEN_2849;
      end
    end else begin
      meta_284_valid_1 <= _GEN_2849;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_284_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_284_lru <= _GEN_8520;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_285_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_285_valid_0 <= _GEN_2338;
        end else begin
          meta_285_valid_0 <= _GEN_7781;
        end
      end else begin
        meta_285_valid_0 <= _GEN_2338;
      end
    end else begin
      meta_285_valid_0 <= _GEN_2338;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_285_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_285_valid_1 <= _GEN_2850;
        end else begin
          meta_285_valid_1 <= _GEN_7782;
        end
      end else begin
        meta_285_valid_1 <= _GEN_2850;
      end
    end else begin
      meta_285_valid_1 <= _GEN_2850;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_285_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_285_lru <= _GEN_8521;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_286_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_286_valid_0 <= _GEN_2339;
        end else begin
          meta_286_valid_0 <= _GEN_7783;
        end
      end else begin
        meta_286_valid_0 <= _GEN_2339;
      end
    end else begin
      meta_286_valid_0 <= _GEN_2339;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_286_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_286_valid_1 <= _GEN_2851;
        end else begin
          meta_286_valid_1 <= _GEN_7784;
        end
      end else begin
        meta_286_valid_1 <= _GEN_2851;
      end
    end else begin
      meta_286_valid_1 <= _GEN_2851;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_286_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_286_lru <= _GEN_8522;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_287_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_287_valid_0 <= _GEN_2340;
        end else begin
          meta_287_valid_0 <= _GEN_7785;
        end
      end else begin
        meta_287_valid_0 <= _GEN_2340;
      end
    end else begin
      meta_287_valid_0 <= _GEN_2340;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_287_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_287_valid_1 <= _GEN_2852;
        end else begin
          meta_287_valid_1 <= _GEN_7786;
        end
      end else begin
        meta_287_valid_1 <= _GEN_2852;
      end
    end else begin
      meta_287_valid_1 <= _GEN_2852;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_287_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_287_lru <= _GEN_8523;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_288_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_288_valid_0 <= _GEN_2341;
        end else begin
          meta_288_valid_0 <= _GEN_7787;
        end
      end else begin
        meta_288_valid_0 <= _GEN_2341;
      end
    end else begin
      meta_288_valid_0 <= _GEN_2341;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_288_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_288_valid_1 <= _GEN_2853;
        end else begin
          meta_288_valid_1 <= _GEN_7788;
        end
      end else begin
        meta_288_valid_1 <= _GEN_2853;
      end
    end else begin
      meta_288_valid_1 <= _GEN_2853;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_288_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_288_lru <= _GEN_8524;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_289_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_289_valid_0 <= _GEN_2342;
        end else begin
          meta_289_valid_0 <= _GEN_7789;
        end
      end else begin
        meta_289_valid_0 <= _GEN_2342;
      end
    end else begin
      meta_289_valid_0 <= _GEN_2342;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_289_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_289_valid_1 <= _GEN_2854;
        end else begin
          meta_289_valid_1 <= _GEN_7790;
        end
      end else begin
        meta_289_valid_1 <= _GEN_2854;
      end
    end else begin
      meta_289_valid_1 <= _GEN_2854;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_289_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_289_lru <= _GEN_8525;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_290_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_290_valid_0 <= _GEN_2343;
        end else begin
          meta_290_valid_0 <= _GEN_7791;
        end
      end else begin
        meta_290_valid_0 <= _GEN_2343;
      end
    end else begin
      meta_290_valid_0 <= _GEN_2343;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_290_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_290_valid_1 <= _GEN_2855;
        end else begin
          meta_290_valid_1 <= _GEN_7792;
        end
      end else begin
        meta_290_valid_1 <= _GEN_2855;
      end
    end else begin
      meta_290_valid_1 <= _GEN_2855;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_290_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_290_lru <= _GEN_8526;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_291_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_291_valid_0 <= _GEN_2344;
        end else begin
          meta_291_valid_0 <= _GEN_7793;
        end
      end else begin
        meta_291_valid_0 <= _GEN_2344;
      end
    end else begin
      meta_291_valid_0 <= _GEN_2344;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_291_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_291_valid_1 <= _GEN_2856;
        end else begin
          meta_291_valid_1 <= _GEN_7794;
        end
      end else begin
        meta_291_valid_1 <= _GEN_2856;
      end
    end else begin
      meta_291_valid_1 <= _GEN_2856;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_291_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_291_lru <= _GEN_8527;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_292_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_292_valid_0 <= _GEN_2345;
        end else begin
          meta_292_valid_0 <= _GEN_7795;
        end
      end else begin
        meta_292_valid_0 <= _GEN_2345;
      end
    end else begin
      meta_292_valid_0 <= _GEN_2345;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_292_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_292_valid_1 <= _GEN_2857;
        end else begin
          meta_292_valid_1 <= _GEN_7796;
        end
      end else begin
        meta_292_valid_1 <= _GEN_2857;
      end
    end else begin
      meta_292_valid_1 <= _GEN_2857;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_292_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_292_lru <= _GEN_8528;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_293_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_293_valid_0 <= _GEN_2346;
        end else begin
          meta_293_valid_0 <= _GEN_7797;
        end
      end else begin
        meta_293_valid_0 <= _GEN_2346;
      end
    end else begin
      meta_293_valid_0 <= _GEN_2346;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_293_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_293_valid_1 <= _GEN_2858;
        end else begin
          meta_293_valid_1 <= _GEN_7798;
        end
      end else begin
        meta_293_valid_1 <= _GEN_2858;
      end
    end else begin
      meta_293_valid_1 <= _GEN_2858;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_293_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_293_lru <= _GEN_8529;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_294_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_294_valid_0 <= _GEN_2347;
        end else begin
          meta_294_valid_0 <= _GEN_7799;
        end
      end else begin
        meta_294_valid_0 <= _GEN_2347;
      end
    end else begin
      meta_294_valid_0 <= _GEN_2347;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_294_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_294_valid_1 <= _GEN_2859;
        end else begin
          meta_294_valid_1 <= _GEN_7800;
        end
      end else begin
        meta_294_valid_1 <= _GEN_2859;
      end
    end else begin
      meta_294_valid_1 <= _GEN_2859;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_294_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_294_lru <= _GEN_8530;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_295_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_295_valid_0 <= _GEN_2348;
        end else begin
          meta_295_valid_0 <= _GEN_7801;
        end
      end else begin
        meta_295_valid_0 <= _GEN_2348;
      end
    end else begin
      meta_295_valid_0 <= _GEN_2348;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_295_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_295_valid_1 <= _GEN_2860;
        end else begin
          meta_295_valid_1 <= _GEN_7802;
        end
      end else begin
        meta_295_valid_1 <= _GEN_2860;
      end
    end else begin
      meta_295_valid_1 <= _GEN_2860;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_295_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_295_lru <= _GEN_8531;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_296_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_296_valid_0 <= _GEN_2349;
        end else begin
          meta_296_valid_0 <= _GEN_7803;
        end
      end else begin
        meta_296_valid_0 <= _GEN_2349;
      end
    end else begin
      meta_296_valid_0 <= _GEN_2349;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_296_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_296_valid_1 <= _GEN_2861;
        end else begin
          meta_296_valid_1 <= _GEN_7804;
        end
      end else begin
        meta_296_valid_1 <= _GEN_2861;
      end
    end else begin
      meta_296_valid_1 <= _GEN_2861;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_296_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_296_lru <= _GEN_8532;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_297_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_297_valid_0 <= _GEN_2350;
        end else begin
          meta_297_valid_0 <= _GEN_7805;
        end
      end else begin
        meta_297_valid_0 <= _GEN_2350;
      end
    end else begin
      meta_297_valid_0 <= _GEN_2350;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_297_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_297_valid_1 <= _GEN_2862;
        end else begin
          meta_297_valid_1 <= _GEN_7806;
        end
      end else begin
        meta_297_valid_1 <= _GEN_2862;
      end
    end else begin
      meta_297_valid_1 <= _GEN_2862;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_297_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_297_lru <= _GEN_8533;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_298_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_298_valid_0 <= _GEN_2351;
        end else begin
          meta_298_valid_0 <= _GEN_7807;
        end
      end else begin
        meta_298_valid_0 <= _GEN_2351;
      end
    end else begin
      meta_298_valid_0 <= _GEN_2351;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_298_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_298_valid_1 <= _GEN_2863;
        end else begin
          meta_298_valid_1 <= _GEN_7808;
        end
      end else begin
        meta_298_valid_1 <= _GEN_2863;
      end
    end else begin
      meta_298_valid_1 <= _GEN_2863;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_298_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_298_lru <= _GEN_8534;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_299_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_299_valid_0 <= _GEN_2352;
        end else begin
          meta_299_valid_0 <= _GEN_7809;
        end
      end else begin
        meta_299_valid_0 <= _GEN_2352;
      end
    end else begin
      meta_299_valid_0 <= _GEN_2352;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_299_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_299_valid_1 <= _GEN_2864;
        end else begin
          meta_299_valid_1 <= _GEN_7810;
        end
      end else begin
        meta_299_valid_1 <= _GEN_2864;
      end
    end else begin
      meta_299_valid_1 <= _GEN_2864;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_299_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_299_lru <= _GEN_8535;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_300_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_300_valid_0 <= _GEN_2353;
        end else begin
          meta_300_valid_0 <= _GEN_7811;
        end
      end else begin
        meta_300_valid_0 <= _GEN_2353;
      end
    end else begin
      meta_300_valid_0 <= _GEN_2353;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_300_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_300_valid_1 <= _GEN_2865;
        end else begin
          meta_300_valid_1 <= _GEN_7812;
        end
      end else begin
        meta_300_valid_1 <= _GEN_2865;
      end
    end else begin
      meta_300_valid_1 <= _GEN_2865;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_300_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_300_lru <= _GEN_8536;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_301_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_301_valid_0 <= _GEN_2354;
        end else begin
          meta_301_valid_0 <= _GEN_7813;
        end
      end else begin
        meta_301_valid_0 <= _GEN_2354;
      end
    end else begin
      meta_301_valid_0 <= _GEN_2354;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_301_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_301_valid_1 <= _GEN_2866;
        end else begin
          meta_301_valid_1 <= _GEN_7814;
        end
      end else begin
        meta_301_valid_1 <= _GEN_2866;
      end
    end else begin
      meta_301_valid_1 <= _GEN_2866;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_301_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_301_lru <= _GEN_8537;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_302_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_302_valid_0 <= _GEN_2355;
        end else begin
          meta_302_valid_0 <= _GEN_7815;
        end
      end else begin
        meta_302_valid_0 <= _GEN_2355;
      end
    end else begin
      meta_302_valid_0 <= _GEN_2355;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_302_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_302_valid_1 <= _GEN_2867;
        end else begin
          meta_302_valid_1 <= _GEN_7816;
        end
      end else begin
        meta_302_valid_1 <= _GEN_2867;
      end
    end else begin
      meta_302_valid_1 <= _GEN_2867;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_302_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_302_lru <= _GEN_8538;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_303_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_303_valid_0 <= _GEN_2356;
        end else begin
          meta_303_valid_0 <= _GEN_7817;
        end
      end else begin
        meta_303_valid_0 <= _GEN_2356;
      end
    end else begin
      meta_303_valid_0 <= _GEN_2356;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_303_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_303_valid_1 <= _GEN_2868;
        end else begin
          meta_303_valid_1 <= _GEN_7818;
        end
      end else begin
        meta_303_valid_1 <= _GEN_2868;
      end
    end else begin
      meta_303_valid_1 <= _GEN_2868;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_303_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_303_lru <= _GEN_8539;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_304_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_304_valid_0 <= _GEN_2357;
        end else begin
          meta_304_valid_0 <= _GEN_7819;
        end
      end else begin
        meta_304_valid_0 <= _GEN_2357;
      end
    end else begin
      meta_304_valid_0 <= _GEN_2357;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_304_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_304_valid_1 <= _GEN_2869;
        end else begin
          meta_304_valid_1 <= _GEN_7820;
        end
      end else begin
        meta_304_valid_1 <= _GEN_2869;
      end
    end else begin
      meta_304_valid_1 <= _GEN_2869;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_304_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_304_lru <= _GEN_8540;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_305_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_305_valid_0 <= _GEN_2358;
        end else begin
          meta_305_valid_0 <= _GEN_7821;
        end
      end else begin
        meta_305_valid_0 <= _GEN_2358;
      end
    end else begin
      meta_305_valid_0 <= _GEN_2358;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_305_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_305_valid_1 <= _GEN_2870;
        end else begin
          meta_305_valid_1 <= _GEN_7822;
        end
      end else begin
        meta_305_valid_1 <= _GEN_2870;
      end
    end else begin
      meta_305_valid_1 <= _GEN_2870;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_305_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_305_lru <= _GEN_8541;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_306_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_306_valid_0 <= _GEN_2359;
        end else begin
          meta_306_valid_0 <= _GEN_7823;
        end
      end else begin
        meta_306_valid_0 <= _GEN_2359;
      end
    end else begin
      meta_306_valid_0 <= _GEN_2359;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_306_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_306_valid_1 <= _GEN_2871;
        end else begin
          meta_306_valid_1 <= _GEN_7824;
        end
      end else begin
        meta_306_valid_1 <= _GEN_2871;
      end
    end else begin
      meta_306_valid_1 <= _GEN_2871;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_306_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_306_lru <= _GEN_8542;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_307_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_307_valid_0 <= _GEN_2360;
        end else begin
          meta_307_valid_0 <= _GEN_7825;
        end
      end else begin
        meta_307_valid_0 <= _GEN_2360;
      end
    end else begin
      meta_307_valid_0 <= _GEN_2360;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_307_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_307_valid_1 <= _GEN_2872;
        end else begin
          meta_307_valid_1 <= _GEN_7826;
        end
      end else begin
        meta_307_valid_1 <= _GEN_2872;
      end
    end else begin
      meta_307_valid_1 <= _GEN_2872;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_307_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_307_lru <= _GEN_8543;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_308_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_308_valid_0 <= _GEN_2361;
        end else begin
          meta_308_valid_0 <= _GEN_7827;
        end
      end else begin
        meta_308_valid_0 <= _GEN_2361;
      end
    end else begin
      meta_308_valid_0 <= _GEN_2361;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_308_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_308_valid_1 <= _GEN_2873;
        end else begin
          meta_308_valid_1 <= _GEN_7828;
        end
      end else begin
        meta_308_valid_1 <= _GEN_2873;
      end
    end else begin
      meta_308_valid_1 <= _GEN_2873;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_308_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_308_lru <= _GEN_8544;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_309_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_309_valid_0 <= _GEN_2362;
        end else begin
          meta_309_valid_0 <= _GEN_7829;
        end
      end else begin
        meta_309_valid_0 <= _GEN_2362;
      end
    end else begin
      meta_309_valid_0 <= _GEN_2362;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_309_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_309_valid_1 <= _GEN_2874;
        end else begin
          meta_309_valid_1 <= _GEN_7830;
        end
      end else begin
        meta_309_valid_1 <= _GEN_2874;
      end
    end else begin
      meta_309_valid_1 <= _GEN_2874;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_309_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_309_lru <= _GEN_8545;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_310_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_310_valid_0 <= _GEN_2363;
        end else begin
          meta_310_valid_0 <= _GEN_7831;
        end
      end else begin
        meta_310_valid_0 <= _GEN_2363;
      end
    end else begin
      meta_310_valid_0 <= _GEN_2363;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_310_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_310_valid_1 <= _GEN_2875;
        end else begin
          meta_310_valid_1 <= _GEN_7832;
        end
      end else begin
        meta_310_valid_1 <= _GEN_2875;
      end
    end else begin
      meta_310_valid_1 <= _GEN_2875;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_310_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_310_lru <= _GEN_8546;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_311_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_311_valid_0 <= _GEN_2364;
        end else begin
          meta_311_valid_0 <= _GEN_7833;
        end
      end else begin
        meta_311_valid_0 <= _GEN_2364;
      end
    end else begin
      meta_311_valid_0 <= _GEN_2364;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_311_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_311_valid_1 <= _GEN_2876;
        end else begin
          meta_311_valid_1 <= _GEN_7834;
        end
      end else begin
        meta_311_valid_1 <= _GEN_2876;
      end
    end else begin
      meta_311_valid_1 <= _GEN_2876;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_311_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_311_lru <= _GEN_8547;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_312_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_312_valid_0 <= _GEN_2365;
        end else begin
          meta_312_valid_0 <= _GEN_7835;
        end
      end else begin
        meta_312_valid_0 <= _GEN_2365;
      end
    end else begin
      meta_312_valid_0 <= _GEN_2365;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_312_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_312_valid_1 <= _GEN_2877;
        end else begin
          meta_312_valid_1 <= _GEN_7836;
        end
      end else begin
        meta_312_valid_1 <= _GEN_2877;
      end
    end else begin
      meta_312_valid_1 <= _GEN_2877;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_312_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_312_lru <= _GEN_8548;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_313_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_313_valid_0 <= _GEN_2366;
        end else begin
          meta_313_valid_0 <= _GEN_7837;
        end
      end else begin
        meta_313_valid_0 <= _GEN_2366;
      end
    end else begin
      meta_313_valid_0 <= _GEN_2366;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_313_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_313_valid_1 <= _GEN_2878;
        end else begin
          meta_313_valid_1 <= _GEN_7838;
        end
      end else begin
        meta_313_valid_1 <= _GEN_2878;
      end
    end else begin
      meta_313_valid_1 <= _GEN_2878;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_313_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_313_lru <= _GEN_8549;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_314_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_314_valid_0 <= _GEN_2367;
        end else begin
          meta_314_valid_0 <= _GEN_7839;
        end
      end else begin
        meta_314_valid_0 <= _GEN_2367;
      end
    end else begin
      meta_314_valid_0 <= _GEN_2367;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_314_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_314_valid_1 <= _GEN_2879;
        end else begin
          meta_314_valid_1 <= _GEN_7840;
        end
      end else begin
        meta_314_valid_1 <= _GEN_2879;
      end
    end else begin
      meta_314_valid_1 <= _GEN_2879;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_314_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_314_lru <= _GEN_8550;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_315_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_315_valid_0 <= _GEN_2368;
        end else begin
          meta_315_valid_0 <= _GEN_7841;
        end
      end else begin
        meta_315_valid_0 <= _GEN_2368;
      end
    end else begin
      meta_315_valid_0 <= _GEN_2368;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_315_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_315_valid_1 <= _GEN_2880;
        end else begin
          meta_315_valid_1 <= _GEN_7842;
        end
      end else begin
        meta_315_valid_1 <= _GEN_2880;
      end
    end else begin
      meta_315_valid_1 <= _GEN_2880;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_315_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_315_lru <= _GEN_8551;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_316_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_316_valid_0 <= _GEN_2369;
        end else begin
          meta_316_valid_0 <= _GEN_7843;
        end
      end else begin
        meta_316_valid_0 <= _GEN_2369;
      end
    end else begin
      meta_316_valid_0 <= _GEN_2369;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_316_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_316_valid_1 <= _GEN_2881;
        end else begin
          meta_316_valid_1 <= _GEN_7844;
        end
      end else begin
        meta_316_valid_1 <= _GEN_2881;
      end
    end else begin
      meta_316_valid_1 <= _GEN_2881;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_316_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_316_lru <= _GEN_8552;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_317_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_317_valid_0 <= _GEN_2370;
        end else begin
          meta_317_valid_0 <= _GEN_7845;
        end
      end else begin
        meta_317_valid_0 <= _GEN_2370;
      end
    end else begin
      meta_317_valid_0 <= _GEN_2370;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_317_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_317_valid_1 <= _GEN_2882;
        end else begin
          meta_317_valid_1 <= _GEN_7846;
        end
      end else begin
        meta_317_valid_1 <= _GEN_2882;
      end
    end else begin
      meta_317_valid_1 <= _GEN_2882;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_317_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_317_lru <= _GEN_8553;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_318_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_318_valid_0 <= _GEN_2371;
        end else begin
          meta_318_valid_0 <= _GEN_7847;
        end
      end else begin
        meta_318_valid_0 <= _GEN_2371;
      end
    end else begin
      meta_318_valid_0 <= _GEN_2371;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_318_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_318_valid_1 <= _GEN_2883;
        end else begin
          meta_318_valid_1 <= _GEN_7848;
        end
      end else begin
        meta_318_valid_1 <= _GEN_2883;
      end
    end else begin
      meta_318_valid_1 <= _GEN_2883;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_318_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_318_lru <= _GEN_8554;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_319_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_319_valid_0 <= _GEN_2372;
        end else begin
          meta_319_valid_0 <= _GEN_7849;
        end
      end else begin
        meta_319_valid_0 <= _GEN_2372;
      end
    end else begin
      meta_319_valid_0 <= _GEN_2372;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_319_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_319_valid_1 <= _GEN_2884;
        end else begin
          meta_319_valid_1 <= _GEN_7850;
        end
      end else begin
        meta_319_valid_1 <= _GEN_2884;
      end
    end else begin
      meta_319_valid_1 <= _GEN_2884;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_319_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_319_lru <= _GEN_8555;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_320_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_320_valid_0 <= _GEN_2373;
        end else begin
          meta_320_valid_0 <= _GEN_7851;
        end
      end else begin
        meta_320_valid_0 <= _GEN_2373;
      end
    end else begin
      meta_320_valid_0 <= _GEN_2373;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_320_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_320_valid_1 <= _GEN_2885;
        end else begin
          meta_320_valid_1 <= _GEN_7852;
        end
      end else begin
        meta_320_valid_1 <= _GEN_2885;
      end
    end else begin
      meta_320_valid_1 <= _GEN_2885;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_320_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_320_lru <= _GEN_8556;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_321_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_321_valid_0 <= _GEN_2374;
        end else begin
          meta_321_valid_0 <= _GEN_7853;
        end
      end else begin
        meta_321_valid_0 <= _GEN_2374;
      end
    end else begin
      meta_321_valid_0 <= _GEN_2374;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_321_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_321_valid_1 <= _GEN_2886;
        end else begin
          meta_321_valid_1 <= _GEN_7854;
        end
      end else begin
        meta_321_valid_1 <= _GEN_2886;
      end
    end else begin
      meta_321_valid_1 <= _GEN_2886;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_321_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_321_lru <= _GEN_8557;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_322_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_322_valid_0 <= _GEN_2375;
        end else begin
          meta_322_valid_0 <= _GEN_7855;
        end
      end else begin
        meta_322_valid_0 <= _GEN_2375;
      end
    end else begin
      meta_322_valid_0 <= _GEN_2375;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_322_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_322_valid_1 <= _GEN_2887;
        end else begin
          meta_322_valid_1 <= _GEN_7856;
        end
      end else begin
        meta_322_valid_1 <= _GEN_2887;
      end
    end else begin
      meta_322_valid_1 <= _GEN_2887;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_322_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_322_lru <= _GEN_8558;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_323_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_323_valid_0 <= _GEN_2376;
        end else begin
          meta_323_valid_0 <= _GEN_7857;
        end
      end else begin
        meta_323_valid_0 <= _GEN_2376;
      end
    end else begin
      meta_323_valid_0 <= _GEN_2376;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_323_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_323_valid_1 <= _GEN_2888;
        end else begin
          meta_323_valid_1 <= _GEN_7858;
        end
      end else begin
        meta_323_valid_1 <= _GEN_2888;
      end
    end else begin
      meta_323_valid_1 <= _GEN_2888;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_323_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_323_lru <= _GEN_8559;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_324_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_324_valid_0 <= _GEN_2377;
        end else begin
          meta_324_valid_0 <= _GEN_7859;
        end
      end else begin
        meta_324_valid_0 <= _GEN_2377;
      end
    end else begin
      meta_324_valid_0 <= _GEN_2377;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_324_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_324_valid_1 <= _GEN_2889;
        end else begin
          meta_324_valid_1 <= _GEN_7860;
        end
      end else begin
        meta_324_valid_1 <= _GEN_2889;
      end
    end else begin
      meta_324_valid_1 <= _GEN_2889;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_324_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_324_lru <= _GEN_8560;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_325_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_325_valid_0 <= _GEN_2378;
        end else begin
          meta_325_valid_0 <= _GEN_7861;
        end
      end else begin
        meta_325_valid_0 <= _GEN_2378;
      end
    end else begin
      meta_325_valid_0 <= _GEN_2378;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_325_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_325_valid_1 <= _GEN_2890;
        end else begin
          meta_325_valid_1 <= _GEN_7862;
        end
      end else begin
        meta_325_valid_1 <= _GEN_2890;
      end
    end else begin
      meta_325_valid_1 <= _GEN_2890;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_325_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_325_lru <= _GEN_8561;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_326_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_326_valid_0 <= _GEN_2379;
        end else begin
          meta_326_valid_0 <= _GEN_7863;
        end
      end else begin
        meta_326_valid_0 <= _GEN_2379;
      end
    end else begin
      meta_326_valid_0 <= _GEN_2379;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_326_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_326_valid_1 <= _GEN_2891;
        end else begin
          meta_326_valid_1 <= _GEN_7864;
        end
      end else begin
        meta_326_valid_1 <= _GEN_2891;
      end
    end else begin
      meta_326_valid_1 <= _GEN_2891;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_326_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_326_lru <= _GEN_8562;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_327_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_327_valid_0 <= _GEN_2380;
        end else begin
          meta_327_valid_0 <= _GEN_7865;
        end
      end else begin
        meta_327_valid_0 <= _GEN_2380;
      end
    end else begin
      meta_327_valid_0 <= _GEN_2380;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_327_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_327_valid_1 <= _GEN_2892;
        end else begin
          meta_327_valid_1 <= _GEN_7866;
        end
      end else begin
        meta_327_valid_1 <= _GEN_2892;
      end
    end else begin
      meta_327_valid_1 <= _GEN_2892;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_327_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_327_lru <= _GEN_8563;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_328_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_328_valid_0 <= _GEN_2381;
        end else begin
          meta_328_valid_0 <= _GEN_7867;
        end
      end else begin
        meta_328_valid_0 <= _GEN_2381;
      end
    end else begin
      meta_328_valid_0 <= _GEN_2381;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_328_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_328_valid_1 <= _GEN_2893;
        end else begin
          meta_328_valid_1 <= _GEN_7868;
        end
      end else begin
        meta_328_valid_1 <= _GEN_2893;
      end
    end else begin
      meta_328_valid_1 <= _GEN_2893;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_328_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_328_lru <= _GEN_8564;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_329_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_329_valid_0 <= _GEN_2382;
        end else begin
          meta_329_valid_0 <= _GEN_7869;
        end
      end else begin
        meta_329_valid_0 <= _GEN_2382;
      end
    end else begin
      meta_329_valid_0 <= _GEN_2382;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_329_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_329_valid_1 <= _GEN_2894;
        end else begin
          meta_329_valid_1 <= _GEN_7870;
        end
      end else begin
        meta_329_valid_1 <= _GEN_2894;
      end
    end else begin
      meta_329_valid_1 <= _GEN_2894;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_329_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_329_lru <= _GEN_8565;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_330_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_330_valid_0 <= _GEN_2383;
        end else begin
          meta_330_valid_0 <= _GEN_7871;
        end
      end else begin
        meta_330_valid_0 <= _GEN_2383;
      end
    end else begin
      meta_330_valid_0 <= _GEN_2383;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_330_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_330_valid_1 <= _GEN_2895;
        end else begin
          meta_330_valid_1 <= _GEN_7872;
        end
      end else begin
        meta_330_valid_1 <= _GEN_2895;
      end
    end else begin
      meta_330_valid_1 <= _GEN_2895;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_330_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_330_lru <= _GEN_8566;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_331_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_331_valid_0 <= _GEN_2384;
        end else begin
          meta_331_valid_0 <= _GEN_7873;
        end
      end else begin
        meta_331_valid_0 <= _GEN_2384;
      end
    end else begin
      meta_331_valid_0 <= _GEN_2384;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_331_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_331_valid_1 <= _GEN_2896;
        end else begin
          meta_331_valid_1 <= _GEN_7874;
        end
      end else begin
        meta_331_valid_1 <= _GEN_2896;
      end
    end else begin
      meta_331_valid_1 <= _GEN_2896;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_331_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_331_lru <= _GEN_8567;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_332_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_332_valid_0 <= _GEN_2385;
        end else begin
          meta_332_valid_0 <= _GEN_7875;
        end
      end else begin
        meta_332_valid_0 <= _GEN_2385;
      end
    end else begin
      meta_332_valid_0 <= _GEN_2385;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_332_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_332_valid_1 <= _GEN_2897;
        end else begin
          meta_332_valid_1 <= _GEN_7876;
        end
      end else begin
        meta_332_valid_1 <= _GEN_2897;
      end
    end else begin
      meta_332_valid_1 <= _GEN_2897;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_332_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_332_lru <= _GEN_8568;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_333_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_333_valid_0 <= _GEN_2386;
        end else begin
          meta_333_valid_0 <= _GEN_7877;
        end
      end else begin
        meta_333_valid_0 <= _GEN_2386;
      end
    end else begin
      meta_333_valid_0 <= _GEN_2386;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_333_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_333_valid_1 <= _GEN_2898;
        end else begin
          meta_333_valid_1 <= _GEN_7878;
        end
      end else begin
        meta_333_valid_1 <= _GEN_2898;
      end
    end else begin
      meta_333_valid_1 <= _GEN_2898;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_333_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_333_lru <= _GEN_8569;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_334_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_334_valid_0 <= _GEN_2387;
        end else begin
          meta_334_valid_0 <= _GEN_7879;
        end
      end else begin
        meta_334_valid_0 <= _GEN_2387;
      end
    end else begin
      meta_334_valid_0 <= _GEN_2387;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_334_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_334_valid_1 <= _GEN_2899;
        end else begin
          meta_334_valid_1 <= _GEN_7880;
        end
      end else begin
        meta_334_valid_1 <= _GEN_2899;
      end
    end else begin
      meta_334_valid_1 <= _GEN_2899;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_334_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_334_lru <= _GEN_8570;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_335_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_335_valid_0 <= _GEN_2388;
        end else begin
          meta_335_valid_0 <= _GEN_7881;
        end
      end else begin
        meta_335_valid_0 <= _GEN_2388;
      end
    end else begin
      meta_335_valid_0 <= _GEN_2388;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_335_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_335_valid_1 <= _GEN_2900;
        end else begin
          meta_335_valid_1 <= _GEN_7882;
        end
      end else begin
        meta_335_valid_1 <= _GEN_2900;
      end
    end else begin
      meta_335_valid_1 <= _GEN_2900;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_335_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_335_lru <= _GEN_8571;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_336_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_336_valid_0 <= _GEN_2389;
        end else begin
          meta_336_valid_0 <= _GEN_7883;
        end
      end else begin
        meta_336_valid_0 <= _GEN_2389;
      end
    end else begin
      meta_336_valid_0 <= _GEN_2389;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_336_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_336_valid_1 <= _GEN_2901;
        end else begin
          meta_336_valid_1 <= _GEN_7884;
        end
      end else begin
        meta_336_valid_1 <= _GEN_2901;
      end
    end else begin
      meta_336_valid_1 <= _GEN_2901;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_336_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_336_lru <= _GEN_8572;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_337_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_337_valid_0 <= _GEN_2390;
        end else begin
          meta_337_valid_0 <= _GEN_7885;
        end
      end else begin
        meta_337_valid_0 <= _GEN_2390;
      end
    end else begin
      meta_337_valid_0 <= _GEN_2390;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_337_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_337_valid_1 <= _GEN_2902;
        end else begin
          meta_337_valid_1 <= _GEN_7886;
        end
      end else begin
        meta_337_valid_1 <= _GEN_2902;
      end
    end else begin
      meta_337_valid_1 <= _GEN_2902;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_337_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_337_lru <= _GEN_8573;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_338_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_338_valid_0 <= _GEN_2391;
        end else begin
          meta_338_valid_0 <= _GEN_7887;
        end
      end else begin
        meta_338_valid_0 <= _GEN_2391;
      end
    end else begin
      meta_338_valid_0 <= _GEN_2391;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_338_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_338_valid_1 <= _GEN_2903;
        end else begin
          meta_338_valid_1 <= _GEN_7888;
        end
      end else begin
        meta_338_valid_1 <= _GEN_2903;
      end
    end else begin
      meta_338_valid_1 <= _GEN_2903;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_338_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_338_lru <= _GEN_8574;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_339_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_339_valid_0 <= _GEN_2392;
        end else begin
          meta_339_valid_0 <= _GEN_7889;
        end
      end else begin
        meta_339_valid_0 <= _GEN_2392;
      end
    end else begin
      meta_339_valid_0 <= _GEN_2392;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_339_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_339_valid_1 <= _GEN_2904;
        end else begin
          meta_339_valid_1 <= _GEN_7890;
        end
      end else begin
        meta_339_valid_1 <= _GEN_2904;
      end
    end else begin
      meta_339_valid_1 <= _GEN_2904;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_339_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_339_lru <= _GEN_8575;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_340_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_340_valid_0 <= _GEN_2393;
        end else begin
          meta_340_valid_0 <= _GEN_7891;
        end
      end else begin
        meta_340_valid_0 <= _GEN_2393;
      end
    end else begin
      meta_340_valid_0 <= _GEN_2393;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_340_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_340_valid_1 <= _GEN_2905;
        end else begin
          meta_340_valid_1 <= _GEN_7892;
        end
      end else begin
        meta_340_valid_1 <= _GEN_2905;
      end
    end else begin
      meta_340_valid_1 <= _GEN_2905;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_340_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_340_lru <= _GEN_8576;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_341_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_341_valid_0 <= _GEN_2394;
        end else begin
          meta_341_valid_0 <= _GEN_7893;
        end
      end else begin
        meta_341_valid_0 <= _GEN_2394;
      end
    end else begin
      meta_341_valid_0 <= _GEN_2394;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_341_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_341_valid_1 <= _GEN_2906;
        end else begin
          meta_341_valid_1 <= _GEN_7894;
        end
      end else begin
        meta_341_valid_1 <= _GEN_2906;
      end
    end else begin
      meta_341_valid_1 <= _GEN_2906;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_341_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_341_lru <= _GEN_8577;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_342_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_342_valid_0 <= _GEN_2395;
        end else begin
          meta_342_valid_0 <= _GEN_7895;
        end
      end else begin
        meta_342_valid_0 <= _GEN_2395;
      end
    end else begin
      meta_342_valid_0 <= _GEN_2395;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_342_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_342_valid_1 <= _GEN_2907;
        end else begin
          meta_342_valid_1 <= _GEN_7896;
        end
      end else begin
        meta_342_valid_1 <= _GEN_2907;
      end
    end else begin
      meta_342_valid_1 <= _GEN_2907;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_342_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_342_lru <= _GEN_8578;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_343_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_343_valid_0 <= _GEN_2396;
        end else begin
          meta_343_valid_0 <= _GEN_7897;
        end
      end else begin
        meta_343_valid_0 <= _GEN_2396;
      end
    end else begin
      meta_343_valid_0 <= _GEN_2396;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_343_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_343_valid_1 <= _GEN_2908;
        end else begin
          meta_343_valid_1 <= _GEN_7898;
        end
      end else begin
        meta_343_valid_1 <= _GEN_2908;
      end
    end else begin
      meta_343_valid_1 <= _GEN_2908;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_343_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_343_lru <= _GEN_8579;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_344_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_344_valid_0 <= _GEN_2397;
        end else begin
          meta_344_valid_0 <= _GEN_7899;
        end
      end else begin
        meta_344_valid_0 <= _GEN_2397;
      end
    end else begin
      meta_344_valid_0 <= _GEN_2397;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_344_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_344_valid_1 <= _GEN_2909;
        end else begin
          meta_344_valid_1 <= _GEN_7900;
        end
      end else begin
        meta_344_valid_1 <= _GEN_2909;
      end
    end else begin
      meta_344_valid_1 <= _GEN_2909;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_344_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_344_lru <= _GEN_8580;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_345_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_345_valid_0 <= _GEN_2398;
        end else begin
          meta_345_valid_0 <= _GEN_7901;
        end
      end else begin
        meta_345_valid_0 <= _GEN_2398;
      end
    end else begin
      meta_345_valid_0 <= _GEN_2398;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_345_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_345_valid_1 <= _GEN_2910;
        end else begin
          meta_345_valid_1 <= _GEN_7902;
        end
      end else begin
        meta_345_valid_1 <= _GEN_2910;
      end
    end else begin
      meta_345_valid_1 <= _GEN_2910;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_345_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_345_lru <= _GEN_8581;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_346_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_346_valid_0 <= _GEN_2399;
        end else begin
          meta_346_valid_0 <= _GEN_7903;
        end
      end else begin
        meta_346_valid_0 <= _GEN_2399;
      end
    end else begin
      meta_346_valid_0 <= _GEN_2399;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_346_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_346_valid_1 <= _GEN_2911;
        end else begin
          meta_346_valid_1 <= _GEN_7904;
        end
      end else begin
        meta_346_valid_1 <= _GEN_2911;
      end
    end else begin
      meta_346_valid_1 <= _GEN_2911;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_346_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_346_lru <= _GEN_8582;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_347_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_347_valid_0 <= _GEN_2400;
        end else begin
          meta_347_valid_0 <= _GEN_7905;
        end
      end else begin
        meta_347_valid_0 <= _GEN_2400;
      end
    end else begin
      meta_347_valid_0 <= _GEN_2400;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_347_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_347_valid_1 <= _GEN_2912;
        end else begin
          meta_347_valid_1 <= _GEN_7906;
        end
      end else begin
        meta_347_valid_1 <= _GEN_2912;
      end
    end else begin
      meta_347_valid_1 <= _GEN_2912;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_347_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_347_lru <= _GEN_8583;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_348_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_348_valid_0 <= _GEN_2401;
        end else begin
          meta_348_valid_0 <= _GEN_7907;
        end
      end else begin
        meta_348_valid_0 <= _GEN_2401;
      end
    end else begin
      meta_348_valid_0 <= _GEN_2401;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_348_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_348_valid_1 <= _GEN_2913;
        end else begin
          meta_348_valid_1 <= _GEN_7908;
        end
      end else begin
        meta_348_valid_1 <= _GEN_2913;
      end
    end else begin
      meta_348_valid_1 <= _GEN_2913;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_348_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_348_lru <= _GEN_8584;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_349_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_349_valid_0 <= _GEN_2402;
        end else begin
          meta_349_valid_0 <= _GEN_7909;
        end
      end else begin
        meta_349_valid_0 <= _GEN_2402;
      end
    end else begin
      meta_349_valid_0 <= _GEN_2402;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_349_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_349_valid_1 <= _GEN_2914;
        end else begin
          meta_349_valid_1 <= _GEN_7910;
        end
      end else begin
        meta_349_valid_1 <= _GEN_2914;
      end
    end else begin
      meta_349_valid_1 <= _GEN_2914;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_349_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_349_lru <= _GEN_8585;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_350_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_350_valid_0 <= _GEN_2403;
        end else begin
          meta_350_valid_0 <= _GEN_7911;
        end
      end else begin
        meta_350_valid_0 <= _GEN_2403;
      end
    end else begin
      meta_350_valid_0 <= _GEN_2403;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_350_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_350_valid_1 <= _GEN_2915;
        end else begin
          meta_350_valid_1 <= _GEN_7912;
        end
      end else begin
        meta_350_valid_1 <= _GEN_2915;
      end
    end else begin
      meta_350_valid_1 <= _GEN_2915;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_350_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_350_lru <= _GEN_8586;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_351_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_351_valid_0 <= _GEN_2404;
        end else begin
          meta_351_valid_0 <= _GEN_7913;
        end
      end else begin
        meta_351_valid_0 <= _GEN_2404;
      end
    end else begin
      meta_351_valid_0 <= _GEN_2404;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_351_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_351_valid_1 <= _GEN_2916;
        end else begin
          meta_351_valid_1 <= _GEN_7914;
        end
      end else begin
        meta_351_valid_1 <= _GEN_2916;
      end
    end else begin
      meta_351_valid_1 <= _GEN_2916;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_351_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_351_lru <= _GEN_8587;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_352_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_352_valid_0 <= _GEN_2405;
        end else begin
          meta_352_valid_0 <= _GEN_7915;
        end
      end else begin
        meta_352_valid_0 <= _GEN_2405;
      end
    end else begin
      meta_352_valid_0 <= _GEN_2405;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_352_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_352_valid_1 <= _GEN_2917;
        end else begin
          meta_352_valid_1 <= _GEN_7916;
        end
      end else begin
        meta_352_valid_1 <= _GEN_2917;
      end
    end else begin
      meta_352_valid_1 <= _GEN_2917;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_352_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_352_lru <= _GEN_8588;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_353_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_353_valid_0 <= _GEN_2406;
        end else begin
          meta_353_valid_0 <= _GEN_7917;
        end
      end else begin
        meta_353_valid_0 <= _GEN_2406;
      end
    end else begin
      meta_353_valid_0 <= _GEN_2406;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_353_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_353_valid_1 <= _GEN_2918;
        end else begin
          meta_353_valid_1 <= _GEN_7918;
        end
      end else begin
        meta_353_valid_1 <= _GEN_2918;
      end
    end else begin
      meta_353_valid_1 <= _GEN_2918;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_353_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_353_lru <= _GEN_8589;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_354_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_354_valid_0 <= _GEN_2407;
        end else begin
          meta_354_valid_0 <= _GEN_7919;
        end
      end else begin
        meta_354_valid_0 <= _GEN_2407;
      end
    end else begin
      meta_354_valid_0 <= _GEN_2407;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_354_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_354_valid_1 <= _GEN_2919;
        end else begin
          meta_354_valid_1 <= _GEN_7920;
        end
      end else begin
        meta_354_valid_1 <= _GEN_2919;
      end
    end else begin
      meta_354_valid_1 <= _GEN_2919;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_354_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_354_lru <= _GEN_8590;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_355_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_355_valid_0 <= _GEN_2408;
        end else begin
          meta_355_valid_0 <= _GEN_7921;
        end
      end else begin
        meta_355_valid_0 <= _GEN_2408;
      end
    end else begin
      meta_355_valid_0 <= _GEN_2408;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_355_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_355_valid_1 <= _GEN_2920;
        end else begin
          meta_355_valid_1 <= _GEN_7922;
        end
      end else begin
        meta_355_valid_1 <= _GEN_2920;
      end
    end else begin
      meta_355_valid_1 <= _GEN_2920;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_355_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_355_lru <= _GEN_8591;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_356_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_356_valid_0 <= _GEN_2409;
        end else begin
          meta_356_valid_0 <= _GEN_7923;
        end
      end else begin
        meta_356_valid_0 <= _GEN_2409;
      end
    end else begin
      meta_356_valid_0 <= _GEN_2409;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_356_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_356_valid_1 <= _GEN_2921;
        end else begin
          meta_356_valid_1 <= _GEN_7924;
        end
      end else begin
        meta_356_valid_1 <= _GEN_2921;
      end
    end else begin
      meta_356_valid_1 <= _GEN_2921;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_356_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_356_lru <= _GEN_8592;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_357_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_357_valid_0 <= _GEN_2410;
        end else begin
          meta_357_valid_0 <= _GEN_7925;
        end
      end else begin
        meta_357_valid_0 <= _GEN_2410;
      end
    end else begin
      meta_357_valid_0 <= _GEN_2410;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_357_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_357_valid_1 <= _GEN_2922;
        end else begin
          meta_357_valid_1 <= _GEN_7926;
        end
      end else begin
        meta_357_valid_1 <= _GEN_2922;
      end
    end else begin
      meta_357_valid_1 <= _GEN_2922;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_357_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_357_lru <= _GEN_8593;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_358_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_358_valid_0 <= _GEN_2411;
        end else begin
          meta_358_valid_0 <= _GEN_7927;
        end
      end else begin
        meta_358_valid_0 <= _GEN_2411;
      end
    end else begin
      meta_358_valid_0 <= _GEN_2411;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_358_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_358_valid_1 <= _GEN_2923;
        end else begin
          meta_358_valid_1 <= _GEN_7928;
        end
      end else begin
        meta_358_valid_1 <= _GEN_2923;
      end
    end else begin
      meta_358_valid_1 <= _GEN_2923;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_358_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_358_lru <= _GEN_8594;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_359_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_359_valid_0 <= _GEN_2412;
        end else begin
          meta_359_valid_0 <= _GEN_7929;
        end
      end else begin
        meta_359_valid_0 <= _GEN_2412;
      end
    end else begin
      meta_359_valid_0 <= _GEN_2412;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_359_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_359_valid_1 <= _GEN_2924;
        end else begin
          meta_359_valid_1 <= _GEN_7930;
        end
      end else begin
        meta_359_valid_1 <= _GEN_2924;
      end
    end else begin
      meta_359_valid_1 <= _GEN_2924;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_359_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_359_lru <= _GEN_8595;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_360_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_360_valid_0 <= _GEN_2413;
        end else begin
          meta_360_valid_0 <= _GEN_7931;
        end
      end else begin
        meta_360_valid_0 <= _GEN_2413;
      end
    end else begin
      meta_360_valid_0 <= _GEN_2413;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_360_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_360_valid_1 <= _GEN_2925;
        end else begin
          meta_360_valid_1 <= _GEN_7932;
        end
      end else begin
        meta_360_valid_1 <= _GEN_2925;
      end
    end else begin
      meta_360_valid_1 <= _GEN_2925;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_360_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_360_lru <= _GEN_8596;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_361_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_361_valid_0 <= _GEN_2414;
        end else begin
          meta_361_valid_0 <= _GEN_7933;
        end
      end else begin
        meta_361_valid_0 <= _GEN_2414;
      end
    end else begin
      meta_361_valid_0 <= _GEN_2414;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_361_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_361_valid_1 <= _GEN_2926;
        end else begin
          meta_361_valid_1 <= _GEN_7934;
        end
      end else begin
        meta_361_valid_1 <= _GEN_2926;
      end
    end else begin
      meta_361_valid_1 <= _GEN_2926;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_361_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_361_lru <= _GEN_8597;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_362_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_362_valid_0 <= _GEN_2415;
        end else begin
          meta_362_valid_0 <= _GEN_7935;
        end
      end else begin
        meta_362_valid_0 <= _GEN_2415;
      end
    end else begin
      meta_362_valid_0 <= _GEN_2415;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_362_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_362_valid_1 <= _GEN_2927;
        end else begin
          meta_362_valid_1 <= _GEN_7936;
        end
      end else begin
        meta_362_valid_1 <= _GEN_2927;
      end
    end else begin
      meta_362_valid_1 <= _GEN_2927;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_362_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_362_lru <= _GEN_8598;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_363_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_363_valid_0 <= _GEN_2416;
        end else begin
          meta_363_valid_0 <= _GEN_7937;
        end
      end else begin
        meta_363_valid_0 <= _GEN_2416;
      end
    end else begin
      meta_363_valid_0 <= _GEN_2416;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_363_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_363_valid_1 <= _GEN_2928;
        end else begin
          meta_363_valid_1 <= _GEN_7938;
        end
      end else begin
        meta_363_valid_1 <= _GEN_2928;
      end
    end else begin
      meta_363_valid_1 <= _GEN_2928;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_363_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_363_lru <= _GEN_8599;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_364_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_364_valid_0 <= _GEN_2417;
        end else begin
          meta_364_valid_0 <= _GEN_7939;
        end
      end else begin
        meta_364_valid_0 <= _GEN_2417;
      end
    end else begin
      meta_364_valid_0 <= _GEN_2417;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_364_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_364_valid_1 <= _GEN_2929;
        end else begin
          meta_364_valid_1 <= _GEN_7940;
        end
      end else begin
        meta_364_valid_1 <= _GEN_2929;
      end
    end else begin
      meta_364_valid_1 <= _GEN_2929;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_364_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_364_lru <= _GEN_8600;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_365_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_365_valid_0 <= _GEN_2418;
        end else begin
          meta_365_valid_0 <= _GEN_7941;
        end
      end else begin
        meta_365_valid_0 <= _GEN_2418;
      end
    end else begin
      meta_365_valid_0 <= _GEN_2418;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_365_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_365_valid_1 <= _GEN_2930;
        end else begin
          meta_365_valid_1 <= _GEN_7942;
        end
      end else begin
        meta_365_valid_1 <= _GEN_2930;
      end
    end else begin
      meta_365_valid_1 <= _GEN_2930;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_365_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_365_lru <= _GEN_8601;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_366_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_366_valid_0 <= _GEN_2419;
        end else begin
          meta_366_valid_0 <= _GEN_7943;
        end
      end else begin
        meta_366_valid_0 <= _GEN_2419;
      end
    end else begin
      meta_366_valid_0 <= _GEN_2419;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_366_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_366_valid_1 <= _GEN_2931;
        end else begin
          meta_366_valid_1 <= _GEN_7944;
        end
      end else begin
        meta_366_valid_1 <= _GEN_2931;
      end
    end else begin
      meta_366_valid_1 <= _GEN_2931;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_366_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_366_lru <= _GEN_8602;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_367_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_367_valid_0 <= _GEN_2420;
        end else begin
          meta_367_valid_0 <= _GEN_7945;
        end
      end else begin
        meta_367_valid_0 <= _GEN_2420;
      end
    end else begin
      meta_367_valid_0 <= _GEN_2420;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_367_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_367_valid_1 <= _GEN_2932;
        end else begin
          meta_367_valid_1 <= _GEN_7946;
        end
      end else begin
        meta_367_valid_1 <= _GEN_2932;
      end
    end else begin
      meta_367_valid_1 <= _GEN_2932;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_367_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_367_lru <= _GEN_8603;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_368_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_368_valid_0 <= _GEN_2421;
        end else begin
          meta_368_valid_0 <= _GEN_7947;
        end
      end else begin
        meta_368_valid_0 <= _GEN_2421;
      end
    end else begin
      meta_368_valid_0 <= _GEN_2421;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_368_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_368_valid_1 <= _GEN_2933;
        end else begin
          meta_368_valid_1 <= _GEN_7948;
        end
      end else begin
        meta_368_valid_1 <= _GEN_2933;
      end
    end else begin
      meta_368_valid_1 <= _GEN_2933;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_368_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_368_lru <= _GEN_8604;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_369_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_369_valid_0 <= _GEN_2422;
        end else begin
          meta_369_valid_0 <= _GEN_7949;
        end
      end else begin
        meta_369_valid_0 <= _GEN_2422;
      end
    end else begin
      meta_369_valid_0 <= _GEN_2422;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_369_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_369_valid_1 <= _GEN_2934;
        end else begin
          meta_369_valid_1 <= _GEN_7950;
        end
      end else begin
        meta_369_valid_1 <= _GEN_2934;
      end
    end else begin
      meta_369_valid_1 <= _GEN_2934;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_369_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_369_lru <= _GEN_8605;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_370_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_370_valid_0 <= _GEN_2423;
        end else begin
          meta_370_valid_0 <= _GEN_7951;
        end
      end else begin
        meta_370_valid_0 <= _GEN_2423;
      end
    end else begin
      meta_370_valid_0 <= _GEN_2423;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_370_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_370_valid_1 <= _GEN_2935;
        end else begin
          meta_370_valid_1 <= _GEN_7952;
        end
      end else begin
        meta_370_valid_1 <= _GEN_2935;
      end
    end else begin
      meta_370_valid_1 <= _GEN_2935;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_370_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_370_lru <= _GEN_8606;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_371_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_371_valid_0 <= _GEN_2424;
        end else begin
          meta_371_valid_0 <= _GEN_7953;
        end
      end else begin
        meta_371_valid_0 <= _GEN_2424;
      end
    end else begin
      meta_371_valid_0 <= _GEN_2424;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_371_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_371_valid_1 <= _GEN_2936;
        end else begin
          meta_371_valid_1 <= _GEN_7954;
        end
      end else begin
        meta_371_valid_1 <= _GEN_2936;
      end
    end else begin
      meta_371_valid_1 <= _GEN_2936;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_371_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_371_lru <= _GEN_8607;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_372_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_372_valid_0 <= _GEN_2425;
        end else begin
          meta_372_valid_0 <= _GEN_7955;
        end
      end else begin
        meta_372_valid_0 <= _GEN_2425;
      end
    end else begin
      meta_372_valid_0 <= _GEN_2425;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_372_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_372_valid_1 <= _GEN_2937;
        end else begin
          meta_372_valid_1 <= _GEN_7956;
        end
      end else begin
        meta_372_valid_1 <= _GEN_2937;
      end
    end else begin
      meta_372_valid_1 <= _GEN_2937;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_372_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_372_lru <= _GEN_8608;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_373_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_373_valid_0 <= _GEN_2426;
        end else begin
          meta_373_valid_0 <= _GEN_7957;
        end
      end else begin
        meta_373_valid_0 <= _GEN_2426;
      end
    end else begin
      meta_373_valid_0 <= _GEN_2426;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_373_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_373_valid_1 <= _GEN_2938;
        end else begin
          meta_373_valid_1 <= _GEN_7958;
        end
      end else begin
        meta_373_valid_1 <= _GEN_2938;
      end
    end else begin
      meta_373_valid_1 <= _GEN_2938;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_373_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_373_lru <= _GEN_8609;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_374_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_374_valid_0 <= _GEN_2427;
        end else begin
          meta_374_valid_0 <= _GEN_7959;
        end
      end else begin
        meta_374_valid_0 <= _GEN_2427;
      end
    end else begin
      meta_374_valid_0 <= _GEN_2427;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_374_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_374_valid_1 <= _GEN_2939;
        end else begin
          meta_374_valid_1 <= _GEN_7960;
        end
      end else begin
        meta_374_valid_1 <= _GEN_2939;
      end
    end else begin
      meta_374_valid_1 <= _GEN_2939;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_374_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_374_lru <= _GEN_8610;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_375_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_375_valid_0 <= _GEN_2428;
        end else begin
          meta_375_valid_0 <= _GEN_7961;
        end
      end else begin
        meta_375_valid_0 <= _GEN_2428;
      end
    end else begin
      meta_375_valid_0 <= _GEN_2428;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_375_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_375_valid_1 <= _GEN_2940;
        end else begin
          meta_375_valid_1 <= _GEN_7962;
        end
      end else begin
        meta_375_valid_1 <= _GEN_2940;
      end
    end else begin
      meta_375_valid_1 <= _GEN_2940;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_375_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_375_lru <= _GEN_8611;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_376_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_376_valid_0 <= _GEN_2429;
        end else begin
          meta_376_valid_0 <= _GEN_7963;
        end
      end else begin
        meta_376_valid_0 <= _GEN_2429;
      end
    end else begin
      meta_376_valid_0 <= _GEN_2429;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_376_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_376_valid_1 <= _GEN_2941;
        end else begin
          meta_376_valid_1 <= _GEN_7964;
        end
      end else begin
        meta_376_valid_1 <= _GEN_2941;
      end
    end else begin
      meta_376_valid_1 <= _GEN_2941;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_376_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_376_lru <= _GEN_8612;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_377_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_377_valid_0 <= _GEN_2430;
        end else begin
          meta_377_valid_0 <= _GEN_7965;
        end
      end else begin
        meta_377_valid_0 <= _GEN_2430;
      end
    end else begin
      meta_377_valid_0 <= _GEN_2430;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_377_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_377_valid_1 <= _GEN_2942;
        end else begin
          meta_377_valid_1 <= _GEN_7966;
        end
      end else begin
        meta_377_valid_1 <= _GEN_2942;
      end
    end else begin
      meta_377_valid_1 <= _GEN_2942;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_377_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_377_lru <= _GEN_8613;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_378_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_378_valid_0 <= _GEN_2431;
        end else begin
          meta_378_valid_0 <= _GEN_7967;
        end
      end else begin
        meta_378_valid_0 <= _GEN_2431;
      end
    end else begin
      meta_378_valid_0 <= _GEN_2431;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_378_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_378_valid_1 <= _GEN_2943;
        end else begin
          meta_378_valid_1 <= _GEN_7968;
        end
      end else begin
        meta_378_valid_1 <= _GEN_2943;
      end
    end else begin
      meta_378_valid_1 <= _GEN_2943;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_378_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_378_lru <= _GEN_8614;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_379_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_379_valid_0 <= _GEN_2432;
        end else begin
          meta_379_valid_0 <= _GEN_7969;
        end
      end else begin
        meta_379_valid_0 <= _GEN_2432;
      end
    end else begin
      meta_379_valid_0 <= _GEN_2432;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_379_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_379_valid_1 <= _GEN_2944;
        end else begin
          meta_379_valid_1 <= _GEN_7970;
        end
      end else begin
        meta_379_valid_1 <= _GEN_2944;
      end
    end else begin
      meta_379_valid_1 <= _GEN_2944;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_379_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_379_lru <= _GEN_8615;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_380_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_380_valid_0 <= _GEN_2433;
        end else begin
          meta_380_valid_0 <= _GEN_7971;
        end
      end else begin
        meta_380_valid_0 <= _GEN_2433;
      end
    end else begin
      meta_380_valid_0 <= _GEN_2433;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_380_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_380_valid_1 <= _GEN_2945;
        end else begin
          meta_380_valid_1 <= _GEN_7972;
        end
      end else begin
        meta_380_valid_1 <= _GEN_2945;
      end
    end else begin
      meta_380_valid_1 <= _GEN_2945;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_380_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_380_lru <= _GEN_8616;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_381_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_381_valid_0 <= _GEN_2434;
        end else begin
          meta_381_valid_0 <= _GEN_7973;
        end
      end else begin
        meta_381_valid_0 <= _GEN_2434;
      end
    end else begin
      meta_381_valid_0 <= _GEN_2434;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_381_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_381_valid_1 <= _GEN_2946;
        end else begin
          meta_381_valid_1 <= _GEN_7974;
        end
      end else begin
        meta_381_valid_1 <= _GEN_2946;
      end
    end else begin
      meta_381_valid_1 <= _GEN_2946;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_381_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_381_lru <= _GEN_8617;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_382_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_382_valid_0 <= _GEN_2435;
        end else begin
          meta_382_valid_0 <= _GEN_7975;
        end
      end else begin
        meta_382_valid_0 <= _GEN_2435;
      end
    end else begin
      meta_382_valid_0 <= _GEN_2435;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_382_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_382_valid_1 <= _GEN_2947;
        end else begin
          meta_382_valid_1 <= _GEN_7976;
        end
      end else begin
        meta_382_valid_1 <= _GEN_2947;
      end
    end else begin
      meta_382_valid_1 <= _GEN_2947;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_382_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_382_lru <= _GEN_8618;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_383_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_383_valid_0 <= _GEN_2436;
        end else begin
          meta_383_valid_0 <= _GEN_7977;
        end
      end else begin
        meta_383_valid_0 <= _GEN_2436;
      end
    end else begin
      meta_383_valid_0 <= _GEN_2436;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_383_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_383_valid_1 <= _GEN_2948;
        end else begin
          meta_383_valid_1 <= _GEN_7978;
        end
      end else begin
        meta_383_valid_1 <= _GEN_2948;
      end
    end else begin
      meta_383_valid_1 <= _GEN_2948;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_383_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_383_lru <= _GEN_8619;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_384_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_384_valid_0 <= _GEN_2437;
        end else begin
          meta_384_valid_0 <= _GEN_7979;
        end
      end else begin
        meta_384_valid_0 <= _GEN_2437;
      end
    end else begin
      meta_384_valid_0 <= _GEN_2437;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_384_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_384_valid_1 <= _GEN_2949;
        end else begin
          meta_384_valid_1 <= _GEN_7980;
        end
      end else begin
        meta_384_valid_1 <= _GEN_2949;
      end
    end else begin
      meta_384_valid_1 <= _GEN_2949;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_384_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_384_lru <= _GEN_8620;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_385_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_385_valid_0 <= _GEN_2438;
        end else begin
          meta_385_valid_0 <= _GEN_7981;
        end
      end else begin
        meta_385_valid_0 <= _GEN_2438;
      end
    end else begin
      meta_385_valid_0 <= _GEN_2438;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_385_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_385_valid_1 <= _GEN_2950;
        end else begin
          meta_385_valid_1 <= _GEN_7982;
        end
      end else begin
        meta_385_valid_1 <= _GEN_2950;
      end
    end else begin
      meta_385_valid_1 <= _GEN_2950;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_385_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_385_lru <= _GEN_8621;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_386_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_386_valid_0 <= _GEN_2439;
        end else begin
          meta_386_valid_0 <= _GEN_7983;
        end
      end else begin
        meta_386_valid_0 <= _GEN_2439;
      end
    end else begin
      meta_386_valid_0 <= _GEN_2439;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_386_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_386_valid_1 <= _GEN_2951;
        end else begin
          meta_386_valid_1 <= _GEN_7984;
        end
      end else begin
        meta_386_valid_1 <= _GEN_2951;
      end
    end else begin
      meta_386_valid_1 <= _GEN_2951;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_386_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_386_lru <= _GEN_8622;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_387_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_387_valid_0 <= _GEN_2440;
        end else begin
          meta_387_valid_0 <= _GEN_7985;
        end
      end else begin
        meta_387_valid_0 <= _GEN_2440;
      end
    end else begin
      meta_387_valid_0 <= _GEN_2440;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_387_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_387_valid_1 <= _GEN_2952;
        end else begin
          meta_387_valid_1 <= _GEN_7986;
        end
      end else begin
        meta_387_valid_1 <= _GEN_2952;
      end
    end else begin
      meta_387_valid_1 <= _GEN_2952;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_387_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_387_lru <= _GEN_8623;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_388_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_388_valid_0 <= _GEN_2441;
        end else begin
          meta_388_valid_0 <= _GEN_7987;
        end
      end else begin
        meta_388_valid_0 <= _GEN_2441;
      end
    end else begin
      meta_388_valid_0 <= _GEN_2441;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_388_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_388_valid_1 <= _GEN_2953;
        end else begin
          meta_388_valid_1 <= _GEN_7988;
        end
      end else begin
        meta_388_valid_1 <= _GEN_2953;
      end
    end else begin
      meta_388_valid_1 <= _GEN_2953;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_388_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_388_lru <= _GEN_8624;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_389_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_389_valid_0 <= _GEN_2442;
        end else begin
          meta_389_valid_0 <= _GEN_7989;
        end
      end else begin
        meta_389_valid_0 <= _GEN_2442;
      end
    end else begin
      meta_389_valid_0 <= _GEN_2442;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_389_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_389_valid_1 <= _GEN_2954;
        end else begin
          meta_389_valid_1 <= _GEN_7990;
        end
      end else begin
        meta_389_valid_1 <= _GEN_2954;
      end
    end else begin
      meta_389_valid_1 <= _GEN_2954;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_389_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_389_lru <= _GEN_8625;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_390_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_390_valid_0 <= _GEN_2443;
        end else begin
          meta_390_valid_0 <= _GEN_7991;
        end
      end else begin
        meta_390_valid_0 <= _GEN_2443;
      end
    end else begin
      meta_390_valid_0 <= _GEN_2443;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_390_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_390_valid_1 <= _GEN_2955;
        end else begin
          meta_390_valid_1 <= _GEN_7992;
        end
      end else begin
        meta_390_valid_1 <= _GEN_2955;
      end
    end else begin
      meta_390_valid_1 <= _GEN_2955;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_390_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_390_lru <= _GEN_8626;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_391_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_391_valid_0 <= _GEN_2444;
        end else begin
          meta_391_valid_0 <= _GEN_7993;
        end
      end else begin
        meta_391_valid_0 <= _GEN_2444;
      end
    end else begin
      meta_391_valid_0 <= _GEN_2444;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_391_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_391_valid_1 <= _GEN_2956;
        end else begin
          meta_391_valid_1 <= _GEN_7994;
        end
      end else begin
        meta_391_valid_1 <= _GEN_2956;
      end
    end else begin
      meta_391_valid_1 <= _GEN_2956;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_391_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_391_lru <= _GEN_8627;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_392_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_392_valid_0 <= _GEN_2445;
        end else begin
          meta_392_valid_0 <= _GEN_7995;
        end
      end else begin
        meta_392_valid_0 <= _GEN_2445;
      end
    end else begin
      meta_392_valid_0 <= _GEN_2445;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_392_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_392_valid_1 <= _GEN_2957;
        end else begin
          meta_392_valid_1 <= _GEN_7996;
        end
      end else begin
        meta_392_valid_1 <= _GEN_2957;
      end
    end else begin
      meta_392_valid_1 <= _GEN_2957;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_392_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_392_lru <= _GEN_8628;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_393_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_393_valid_0 <= _GEN_2446;
        end else begin
          meta_393_valid_0 <= _GEN_7997;
        end
      end else begin
        meta_393_valid_0 <= _GEN_2446;
      end
    end else begin
      meta_393_valid_0 <= _GEN_2446;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_393_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_393_valid_1 <= _GEN_2958;
        end else begin
          meta_393_valid_1 <= _GEN_7998;
        end
      end else begin
        meta_393_valid_1 <= _GEN_2958;
      end
    end else begin
      meta_393_valid_1 <= _GEN_2958;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_393_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_393_lru <= _GEN_8629;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_394_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_394_valid_0 <= _GEN_2447;
        end else begin
          meta_394_valid_0 <= _GEN_7999;
        end
      end else begin
        meta_394_valid_0 <= _GEN_2447;
      end
    end else begin
      meta_394_valid_0 <= _GEN_2447;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_394_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_394_valid_1 <= _GEN_2959;
        end else begin
          meta_394_valid_1 <= _GEN_8000;
        end
      end else begin
        meta_394_valid_1 <= _GEN_2959;
      end
    end else begin
      meta_394_valid_1 <= _GEN_2959;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_394_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_394_lru <= _GEN_8630;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_395_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_395_valid_0 <= _GEN_2448;
        end else begin
          meta_395_valid_0 <= _GEN_8001;
        end
      end else begin
        meta_395_valid_0 <= _GEN_2448;
      end
    end else begin
      meta_395_valid_0 <= _GEN_2448;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_395_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_395_valid_1 <= _GEN_2960;
        end else begin
          meta_395_valid_1 <= _GEN_8002;
        end
      end else begin
        meta_395_valid_1 <= _GEN_2960;
      end
    end else begin
      meta_395_valid_1 <= _GEN_2960;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_395_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_395_lru <= _GEN_8631;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_396_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_396_valid_0 <= _GEN_2449;
        end else begin
          meta_396_valid_0 <= _GEN_8003;
        end
      end else begin
        meta_396_valid_0 <= _GEN_2449;
      end
    end else begin
      meta_396_valid_0 <= _GEN_2449;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_396_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_396_valid_1 <= _GEN_2961;
        end else begin
          meta_396_valid_1 <= _GEN_8004;
        end
      end else begin
        meta_396_valid_1 <= _GEN_2961;
      end
    end else begin
      meta_396_valid_1 <= _GEN_2961;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_396_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_396_lru <= _GEN_8632;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_397_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_397_valid_0 <= _GEN_2450;
        end else begin
          meta_397_valid_0 <= _GEN_8005;
        end
      end else begin
        meta_397_valid_0 <= _GEN_2450;
      end
    end else begin
      meta_397_valid_0 <= _GEN_2450;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_397_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_397_valid_1 <= _GEN_2962;
        end else begin
          meta_397_valid_1 <= _GEN_8006;
        end
      end else begin
        meta_397_valid_1 <= _GEN_2962;
      end
    end else begin
      meta_397_valid_1 <= _GEN_2962;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_397_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_397_lru <= _GEN_8633;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_398_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_398_valid_0 <= _GEN_2451;
        end else begin
          meta_398_valid_0 <= _GEN_8007;
        end
      end else begin
        meta_398_valid_0 <= _GEN_2451;
      end
    end else begin
      meta_398_valid_0 <= _GEN_2451;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_398_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_398_valid_1 <= _GEN_2963;
        end else begin
          meta_398_valid_1 <= _GEN_8008;
        end
      end else begin
        meta_398_valid_1 <= _GEN_2963;
      end
    end else begin
      meta_398_valid_1 <= _GEN_2963;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_398_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_398_lru <= _GEN_8634;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_399_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_399_valid_0 <= _GEN_2452;
        end else begin
          meta_399_valid_0 <= _GEN_8009;
        end
      end else begin
        meta_399_valid_0 <= _GEN_2452;
      end
    end else begin
      meta_399_valid_0 <= _GEN_2452;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_399_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_399_valid_1 <= _GEN_2964;
        end else begin
          meta_399_valid_1 <= _GEN_8010;
        end
      end else begin
        meta_399_valid_1 <= _GEN_2964;
      end
    end else begin
      meta_399_valid_1 <= _GEN_2964;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_399_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_399_lru <= _GEN_8635;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_400_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_400_valid_0 <= _GEN_2453;
        end else begin
          meta_400_valid_0 <= _GEN_8011;
        end
      end else begin
        meta_400_valid_0 <= _GEN_2453;
      end
    end else begin
      meta_400_valid_0 <= _GEN_2453;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_400_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_400_valid_1 <= _GEN_2965;
        end else begin
          meta_400_valid_1 <= _GEN_8012;
        end
      end else begin
        meta_400_valid_1 <= _GEN_2965;
      end
    end else begin
      meta_400_valid_1 <= _GEN_2965;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_400_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_400_lru <= _GEN_8636;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_401_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_401_valid_0 <= _GEN_2454;
        end else begin
          meta_401_valid_0 <= _GEN_8013;
        end
      end else begin
        meta_401_valid_0 <= _GEN_2454;
      end
    end else begin
      meta_401_valid_0 <= _GEN_2454;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_401_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_401_valid_1 <= _GEN_2966;
        end else begin
          meta_401_valid_1 <= _GEN_8014;
        end
      end else begin
        meta_401_valid_1 <= _GEN_2966;
      end
    end else begin
      meta_401_valid_1 <= _GEN_2966;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_401_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_401_lru <= _GEN_8637;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_402_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_402_valid_0 <= _GEN_2455;
        end else begin
          meta_402_valid_0 <= _GEN_8015;
        end
      end else begin
        meta_402_valid_0 <= _GEN_2455;
      end
    end else begin
      meta_402_valid_0 <= _GEN_2455;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_402_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_402_valid_1 <= _GEN_2967;
        end else begin
          meta_402_valid_1 <= _GEN_8016;
        end
      end else begin
        meta_402_valid_1 <= _GEN_2967;
      end
    end else begin
      meta_402_valid_1 <= _GEN_2967;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_402_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_402_lru <= _GEN_8638;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_403_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_403_valid_0 <= _GEN_2456;
        end else begin
          meta_403_valid_0 <= _GEN_8017;
        end
      end else begin
        meta_403_valid_0 <= _GEN_2456;
      end
    end else begin
      meta_403_valid_0 <= _GEN_2456;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_403_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_403_valid_1 <= _GEN_2968;
        end else begin
          meta_403_valid_1 <= _GEN_8018;
        end
      end else begin
        meta_403_valid_1 <= _GEN_2968;
      end
    end else begin
      meta_403_valid_1 <= _GEN_2968;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_403_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_403_lru <= _GEN_8639;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_404_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_404_valid_0 <= _GEN_2457;
        end else begin
          meta_404_valid_0 <= _GEN_8019;
        end
      end else begin
        meta_404_valid_0 <= _GEN_2457;
      end
    end else begin
      meta_404_valid_0 <= _GEN_2457;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_404_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_404_valid_1 <= _GEN_2969;
        end else begin
          meta_404_valid_1 <= _GEN_8020;
        end
      end else begin
        meta_404_valid_1 <= _GEN_2969;
      end
    end else begin
      meta_404_valid_1 <= _GEN_2969;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_404_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_404_lru <= _GEN_8640;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_405_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_405_valid_0 <= _GEN_2458;
        end else begin
          meta_405_valid_0 <= _GEN_8021;
        end
      end else begin
        meta_405_valid_0 <= _GEN_2458;
      end
    end else begin
      meta_405_valid_0 <= _GEN_2458;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_405_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_405_valid_1 <= _GEN_2970;
        end else begin
          meta_405_valid_1 <= _GEN_8022;
        end
      end else begin
        meta_405_valid_1 <= _GEN_2970;
      end
    end else begin
      meta_405_valid_1 <= _GEN_2970;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_405_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_405_lru <= _GEN_8641;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_406_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_406_valid_0 <= _GEN_2459;
        end else begin
          meta_406_valid_0 <= _GEN_8023;
        end
      end else begin
        meta_406_valid_0 <= _GEN_2459;
      end
    end else begin
      meta_406_valid_0 <= _GEN_2459;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_406_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_406_valid_1 <= _GEN_2971;
        end else begin
          meta_406_valid_1 <= _GEN_8024;
        end
      end else begin
        meta_406_valid_1 <= _GEN_2971;
      end
    end else begin
      meta_406_valid_1 <= _GEN_2971;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_406_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_406_lru <= _GEN_8642;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_407_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_407_valid_0 <= _GEN_2460;
        end else begin
          meta_407_valid_0 <= _GEN_8025;
        end
      end else begin
        meta_407_valid_0 <= _GEN_2460;
      end
    end else begin
      meta_407_valid_0 <= _GEN_2460;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_407_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_407_valid_1 <= _GEN_2972;
        end else begin
          meta_407_valid_1 <= _GEN_8026;
        end
      end else begin
        meta_407_valid_1 <= _GEN_2972;
      end
    end else begin
      meta_407_valid_1 <= _GEN_2972;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_407_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_407_lru <= _GEN_8643;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_408_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_408_valid_0 <= _GEN_2461;
        end else begin
          meta_408_valid_0 <= _GEN_8027;
        end
      end else begin
        meta_408_valid_0 <= _GEN_2461;
      end
    end else begin
      meta_408_valid_0 <= _GEN_2461;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_408_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_408_valid_1 <= _GEN_2973;
        end else begin
          meta_408_valid_1 <= _GEN_8028;
        end
      end else begin
        meta_408_valid_1 <= _GEN_2973;
      end
    end else begin
      meta_408_valid_1 <= _GEN_2973;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_408_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_408_lru <= _GEN_8644;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_409_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_409_valid_0 <= _GEN_2462;
        end else begin
          meta_409_valid_0 <= _GEN_8029;
        end
      end else begin
        meta_409_valid_0 <= _GEN_2462;
      end
    end else begin
      meta_409_valid_0 <= _GEN_2462;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_409_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_409_valid_1 <= _GEN_2974;
        end else begin
          meta_409_valid_1 <= _GEN_8030;
        end
      end else begin
        meta_409_valid_1 <= _GEN_2974;
      end
    end else begin
      meta_409_valid_1 <= _GEN_2974;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_409_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_409_lru <= _GEN_8645;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_410_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_410_valid_0 <= _GEN_2463;
        end else begin
          meta_410_valid_0 <= _GEN_8031;
        end
      end else begin
        meta_410_valid_0 <= _GEN_2463;
      end
    end else begin
      meta_410_valid_0 <= _GEN_2463;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_410_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_410_valid_1 <= _GEN_2975;
        end else begin
          meta_410_valid_1 <= _GEN_8032;
        end
      end else begin
        meta_410_valid_1 <= _GEN_2975;
      end
    end else begin
      meta_410_valid_1 <= _GEN_2975;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_410_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_410_lru <= _GEN_8646;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_411_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_411_valid_0 <= _GEN_2464;
        end else begin
          meta_411_valid_0 <= _GEN_8033;
        end
      end else begin
        meta_411_valid_0 <= _GEN_2464;
      end
    end else begin
      meta_411_valid_0 <= _GEN_2464;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_411_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_411_valid_1 <= _GEN_2976;
        end else begin
          meta_411_valid_1 <= _GEN_8034;
        end
      end else begin
        meta_411_valid_1 <= _GEN_2976;
      end
    end else begin
      meta_411_valid_1 <= _GEN_2976;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_411_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_411_lru <= _GEN_8647;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_412_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_412_valid_0 <= _GEN_2465;
        end else begin
          meta_412_valid_0 <= _GEN_8035;
        end
      end else begin
        meta_412_valid_0 <= _GEN_2465;
      end
    end else begin
      meta_412_valid_0 <= _GEN_2465;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_412_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_412_valid_1 <= _GEN_2977;
        end else begin
          meta_412_valid_1 <= _GEN_8036;
        end
      end else begin
        meta_412_valid_1 <= _GEN_2977;
      end
    end else begin
      meta_412_valid_1 <= _GEN_2977;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_412_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_412_lru <= _GEN_8648;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_413_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_413_valid_0 <= _GEN_2466;
        end else begin
          meta_413_valid_0 <= _GEN_8037;
        end
      end else begin
        meta_413_valid_0 <= _GEN_2466;
      end
    end else begin
      meta_413_valid_0 <= _GEN_2466;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_413_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_413_valid_1 <= _GEN_2978;
        end else begin
          meta_413_valid_1 <= _GEN_8038;
        end
      end else begin
        meta_413_valid_1 <= _GEN_2978;
      end
    end else begin
      meta_413_valid_1 <= _GEN_2978;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_413_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_413_lru <= _GEN_8649;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_414_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_414_valid_0 <= _GEN_2467;
        end else begin
          meta_414_valid_0 <= _GEN_8039;
        end
      end else begin
        meta_414_valid_0 <= _GEN_2467;
      end
    end else begin
      meta_414_valid_0 <= _GEN_2467;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_414_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_414_valid_1 <= _GEN_2979;
        end else begin
          meta_414_valid_1 <= _GEN_8040;
        end
      end else begin
        meta_414_valid_1 <= _GEN_2979;
      end
    end else begin
      meta_414_valid_1 <= _GEN_2979;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_414_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_414_lru <= _GEN_8650;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_415_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_415_valid_0 <= _GEN_2468;
        end else begin
          meta_415_valid_0 <= _GEN_8041;
        end
      end else begin
        meta_415_valid_0 <= _GEN_2468;
      end
    end else begin
      meta_415_valid_0 <= _GEN_2468;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_415_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_415_valid_1 <= _GEN_2980;
        end else begin
          meta_415_valid_1 <= _GEN_8042;
        end
      end else begin
        meta_415_valid_1 <= _GEN_2980;
      end
    end else begin
      meta_415_valid_1 <= _GEN_2980;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_415_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_415_lru <= _GEN_8651;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_416_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_416_valid_0 <= _GEN_2469;
        end else begin
          meta_416_valid_0 <= _GEN_8043;
        end
      end else begin
        meta_416_valid_0 <= _GEN_2469;
      end
    end else begin
      meta_416_valid_0 <= _GEN_2469;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_416_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_416_valid_1 <= _GEN_2981;
        end else begin
          meta_416_valid_1 <= _GEN_8044;
        end
      end else begin
        meta_416_valid_1 <= _GEN_2981;
      end
    end else begin
      meta_416_valid_1 <= _GEN_2981;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_416_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_416_lru <= _GEN_8652;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_417_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_417_valid_0 <= _GEN_2470;
        end else begin
          meta_417_valid_0 <= _GEN_8045;
        end
      end else begin
        meta_417_valid_0 <= _GEN_2470;
      end
    end else begin
      meta_417_valid_0 <= _GEN_2470;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_417_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_417_valid_1 <= _GEN_2982;
        end else begin
          meta_417_valid_1 <= _GEN_8046;
        end
      end else begin
        meta_417_valid_1 <= _GEN_2982;
      end
    end else begin
      meta_417_valid_1 <= _GEN_2982;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_417_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_417_lru <= _GEN_8653;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_418_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_418_valid_0 <= _GEN_2471;
        end else begin
          meta_418_valid_0 <= _GEN_8047;
        end
      end else begin
        meta_418_valid_0 <= _GEN_2471;
      end
    end else begin
      meta_418_valid_0 <= _GEN_2471;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_418_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_418_valid_1 <= _GEN_2983;
        end else begin
          meta_418_valid_1 <= _GEN_8048;
        end
      end else begin
        meta_418_valid_1 <= _GEN_2983;
      end
    end else begin
      meta_418_valid_1 <= _GEN_2983;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_418_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_418_lru <= _GEN_8654;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_419_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_419_valid_0 <= _GEN_2472;
        end else begin
          meta_419_valid_0 <= _GEN_8049;
        end
      end else begin
        meta_419_valid_0 <= _GEN_2472;
      end
    end else begin
      meta_419_valid_0 <= _GEN_2472;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_419_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_419_valid_1 <= _GEN_2984;
        end else begin
          meta_419_valid_1 <= _GEN_8050;
        end
      end else begin
        meta_419_valid_1 <= _GEN_2984;
      end
    end else begin
      meta_419_valid_1 <= _GEN_2984;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_419_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_419_lru <= _GEN_8655;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_420_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_420_valid_0 <= _GEN_2473;
        end else begin
          meta_420_valid_0 <= _GEN_8051;
        end
      end else begin
        meta_420_valid_0 <= _GEN_2473;
      end
    end else begin
      meta_420_valid_0 <= _GEN_2473;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_420_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_420_valid_1 <= _GEN_2985;
        end else begin
          meta_420_valid_1 <= _GEN_8052;
        end
      end else begin
        meta_420_valid_1 <= _GEN_2985;
      end
    end else begin
      meta_420_valid_1 <= _GEN_2985;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_420_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_420_lru <= _GEN_8656;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_421_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_421_valid_0 <= _GEN_2474;
        end else begin
          meta_421_valid_0 <= _GEN_8053;
        end
      end else begin
        meta_421_valid_0 <= _GEN_2474;
      end
    end else begin
      meta_421_valid_0 <= _GEN_2474;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_421_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_421_valid_1 <= _GEN_2986;
        end else begin
          meta_421_valid_1 <= _GEN_8054;
        end
      end else begin
        meta_421_valid_1 <= _GEN_2986;
      end
    end else begin
      meta_421_valid_1 <= _GEN_2986;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_421_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_421_lru <= _GEN_8657;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_422_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_422_valid_0 <= _GEN_2475;
        end else begin
          meta_422_valid_0 <= _GEN_8055;
        end
      end else begin
        meta_422_valid_0 <= _GEN_2475;
      end
    end else begin
      meta_422_valid_0 <= _GEN_2475;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_422_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_422_valid_1 <= _GEN_2987;
        end else begin
          meta_422_valid_1 <= _GEN_8056;
        end
      end else begin
        meta_422_valid_1 <= _GEN_2987;
      end
    end else begin
      meta_422_valid_1 <= _GEN_2987;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_422_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_422_lru <= _GEN_8658;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_423_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_423_valid_0 <= _GEN_2476;
        end else begin
          meta_423_valid_0 <= _GEN_8057;
        end
      end else begin
        meta_423_valid_0 <= _GEN_2476;
      end
    end else begin
      meta_423_valid_0 <= _GEN_2476;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_423_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_423_valid_1 <= _GEN_2988;
        end else begin
          meta_423_valid_1 <= _GEN_8058;
        end
      end else begin
        meta_423_valid_1 <= _GEN_2988;
      end
    end else begin
      meta_423_valid_1 <= _GEN_2988;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_423_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_423_lru <= _GEN_8659;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_424_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_424_valid_0 <= _GEN_2477;
        end else begin
          meta_424_valid_0 <= _GEN_8059;
        end
      end else begin
        meta_424_valid_0 <= _GEN_2477;
      end
    end else begin
      meta_424_valid_0 <= _GEN_2477;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_424_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_424_valid_1 <= _GEN_2989;
        end else begin
          meta_424_valid_1 <= _GEN_8060;
        end
      end else begin
        meta_424_valid_1 <= _GEN_2989;
      end
    end else begin
      meta_424_valid_1 <= _GEN_2989;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_424_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_424_lru <= _GEN_8660;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_425_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_425_valid_0 <= _GEN_2478;
        end else begin
          meta_425_valid_0 <= _GEN_8061;
        end
      end else begin
        meta_425_valid_0 <= _GEN_2478;
      end
    end else begin
      meta_425_valid_0 <= _GEN_2478;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_425_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_425_valid_1 <= _GEN_2990;
        end else begin
          meta_425_valid_1 <= _GEN_8062;
        end
      end else begin
        meta_425_valid_1 <= _GEN_2990;
      end
    end else begin
      meta_425_valid_1 <= _GEN_2990;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_425_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_425_lru <= _GEN_8661;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_426_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_426_valid_0 <= _GEN_2479;
        end else begin
          meta_426_valid_0 <= _GEN_8063;
        end
      end else begin
        meta_426_valid_0 <= _GEN_2479;
      end
    end else begin
      meta_426_valid_0 <= _GEN_2479;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_426_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_426_valid_1 <= _GEN_2991;
        end else begin
          meta_426_valid_1 <= _GEN_8064;
        end
      end else begin
        meta_426_valid_1 <= _GEN_2991;
      end
    end else begin
      meta_426_valid_1 <= _GEN_2991;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_426_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_426_lru <= _GEN_8662;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_427_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_427_valid_0 <= _GEN_2480;
        end else begin
          meta_427_valid_0 <= _GEN_8065;
        end
      end else begin
        meta_427_valid_0 <= _GEN_2480;
      end
    end else begin
      meta_427_valid_0 <= _GEN_2480;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_427_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_427_valid_1 <= _GEN_2992;
        end else begin
          meta_427_valid_1 <= _GEN_8066;
        end
      end else begin
        meta_427_valid_1 <= _GEN_2992;
      end
    end else begin
      meta_427_valid_1 <= _GEN_2992;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_427_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_427_lru <= _GEN_8663;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_428_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_428_valid_0 <= _GEN_2481;
        end else begin
          meta_428_valid_0 <= _GEN_8067;
        end
      end else begin
        meta_428_valid_0 <= _GEN_2481;
      end
    end else begin
      meta_428_valid_0 <= _GEN_2481;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_428_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_428_valid_1 <= _GEN_2993;
        end else begin
          meta_428_valid_1 <= _GEN_8068;
        end
      end else begin
        meta_428_valid_1 <= _GEN_2993;
      end
    end else begin
      meta_428_valid_1 <= _GEN_2993;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_428_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_428_lru <= _GEN_8664;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_429_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_429_valid_0 <= _GEN_2482;
        end else begin
          meta_429_valid_0 <= _GEN_8069;
        end
      end else begin
        meta_429_valid_0 <= _GEN_2482;
      end
    end else begin
      meta_429_valid_0 <= _GEN_2482;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_429_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_429_valid_1 <= _GEN_2994;
        end else begin
          meta_429_valid_1 <= _GEN_8070;
        end
      end else begin
        meta_429_valid_1 <= _GEN_2994;
      end
    end else begin
      meta_429_valid_1 <= _GEN_2994;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_429_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_429_lru <= _GEN_8665;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_430_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_430_valid_0 <= _GEN_2483;
        end else begin
          meta_430_valid_0 <= _GEN_8071;
        end
      end else begin
        meta_430_valid_0 <= _GEN_2483;
      end
    end else begin
      meta_430_valid_0 <= _GEN_2483;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_430_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_430_valid_1 <= _GEN_2995;
        end else begin
          meta_430_valid_1 <= _GEN_8072;
        end
      end else begin
        meta_430_valid_1 <= _GEN_2995;
      end
    end else begin
      meta_430_valid_1 <= _GEN_2995;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_430_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_430_lru <= _GEN_8666;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_431_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_431_valid_0 <= _GEN_2484;
        end else begin
          meta_431_valid_0 <= _GEN_8073;
        end
      end else begin
        meta_431_valid_0 <= _GEN_2484;
      end
    end else begin
      meta_431_valid_0 <= _GEN_2484;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_431_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_431_valid_1 <= _GEN_2996;
        end else begin
          meta_431_valid_1 <= _GEN_8074;
        end
      end else begin
        meta_431_valid_1 <= _GEN_2996;
      end
    end else begin
      meta_431_valid_1 <= _GEN_2996;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_431_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_431_lru <= _GEN_8667;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_432_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_432_valid_0 <= _GEN_2485;
        end else begin
          meta_432_valid_0 <= _GEN_8075;
        end
      end else begin
        meta_432_valid_0 <= _GEN_2485;
      end
    end else begin
      meta_432_valid_0 <= _GEN_2485;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_432_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_432_valid_1 <= _GEN_2997;
        end else begin
          meta_432_valid_1 <= _GEN_8076;
        end
      end else begin
        meta_432_valid_1 <= _GEN_2997;
      end
    end else begin
      meta_432_valid_1 <= _GEN_2997;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_432_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_432_lru <= _GEN_8668;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_433_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_433_valid_0 <= _GEN_2486;
        end else begin
          meta_433_valid_0 <= _GEN_8077;
        end
      end else begin
        meta_433_valid_0 <= _GEN_2486;
      end
    end else begin
      meta_433_valid_0 <= _GEN_2486;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_433_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_433_valid_1 <= _GEN_2998;
        end else begin
          meta_433_valid_1 <= _GEN_8078;
        end
      end else begin
        meta_433_valid_1 <= _GEN_2998;
      end
    end else begin
      meta_433_valid_1 <= _GEN_2998;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_433_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_433_lru <= _GEN_8669;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_434_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_434_valid_0 <= _GEN_2487;
        end else begin
          meta_434_valid_0 <= _GEN_8079;
        end
      end else begin
        meta_434_valid_0 <= _GEN_2487;
      end
    end else begin
      meta_434_valid_0 <= _GEN_2487;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_434_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_434_valid_1 <= _GEN_2999;
        end else begin
          meta_434_valid_1 <= _GEN_8080;
        end
      end else begin
        meta_434_valid_1 <= _GEN_2999;
      end
    end else begin
      meta_434_valid_1 <= _GEN_2999;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_434_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_434_lru <= _GEN_8670;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_435_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_435_valid_0 <= _GEN_2488;
        end else begin
          meta_435_valid_0 <= _GEN_8081;
        end
      end else begin
        meta_435_valid_0 <= _GEN_2488;
      end
    end else begin
      meta_435_valid_0 <= _GEN_2488;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_435_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_435_valid_1 <= _GEN_3000;
        end else begin
          meta_435_valid_1 <= _GEN_8082;
        end
      end else begin
        meta_435_valid_1 <= _GEN_3000;
      end
    end else begin
      meta_435_valid_1 <= _GEN_3000;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_435_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_435_lru <= _GEN_8671;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_436_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_436_valid_0 <= _GEN_2489;
        end else begin
          meta_436_valid_0 <= _GEN_8083;
        end
      end else begin
        meta_436_valid_0 <= _GEN_2489;
      end
    end else begin
      meta_436_valid_0 <= _GEN_2489;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_436_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_436_valid_1 <= _GEN_3001;
        end else begin
          meta_436_valid_1 <= _GEN_8084;
        end
      end else begin
        meta_436_valid_1 <= _GEN_3001;
      end
    end else begin
      meta_436_valid_1 <= _GEN_3001;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_436_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_436_lru <= _GEN_8672;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_437_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_437_valid_0 <= _GEN_2490;
        end else begin
          meta_437_valid_0 <= _GEN_8085;
        end
      end else begin
        meta_437_valid_0 <= _GEN_2490;
      end
    end else begin
      meta_437_valid_0 <= _GEN_2490;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_437_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_437_valid_1 <= _GEN_3002;
        end else begin
          meta_437_valid_1 <= _GEN_8086;
        end
      end else begin
        meta_437_valid_1 <= _GEN_3002;
      end
    end else begin
      meta_437_valid_1 <= _GEN_3002;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_437_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_437_lru <= _GEN_8673;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_438_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_438_valid_0 <= _GEN_2491;
        end else begin
          meta_438_valid_0 <= _GEN_8087;
        end
      end else begin
        meta_438_valid_0 <= _GEN_2491;
      end
    end else begin
      meta_438_valid_0 <= _GEN_2491;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_438_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_438_valid_1 <= _GEN_3003;
        end else begin
          meta_438_valid_1 <= _GEN_8088;
        end
      end else begin
        meta_438_valid_1 <= _GEN_3003;
      end
    end else begin
      meta_438_valid_1 <= _GEN_3003;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_438_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_438_lru <= _GEN_8674;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_439_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_439_valid_0 <= _GEN_2492;
        end else begin
          meta_439_valid_0 <= _GEN_8089;
        end
      end else begin
        meta_439_valid_0 <= _GEN_2492;
      end
    end else begin
      meta_439_valid_0 <= _GEN_2492;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_439_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_439_valid_1 <= _GEN_3004;
        end else begin
          meta_439_valid_1 <= _GEN_8090;
        end
      end else begin
        meta_439_valid_1 <= _GEN_3004;
      end
    end else begin
      meta_439_valid_1 <= _GEN_3004;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_439_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_439_lru <= _GEN_8675;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_440_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_440_valid_0 <= _GEN_2493;
        end else begin
          meta_440_valid_0 <= _GEN_8091;
        end
      end else begin
        meta_440_valid_0 <= _GEN_2493;
      end
    end else begin
      meta_440_valid_0 <= _GEN_2493;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_440_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_440_valid_1 <= _GEN_3005;
        end else begin
          meta_440_valid_1 <= _GEN_8092;
        end
      end else begin
        meta_440_valid_1 <= _GEN_3005;
      end
    end else begin
      meta_440_valid_1 <= _GEN_3005;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_440_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_440_lru <= _GEN_8676;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_441_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_441_valid_0 <= _GEN_2494;
        end else begin
          meta_441_valid_0 <= _GEN_8093;
        end
      end else begin
        meta_441_valid_0 <= _GEN_2494;
      end
    end else begin
      meta_441_valid_0 <= _GEN_2494;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_441_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_441_valid_1 <= _GEN_3006;
        end else begin
          meta_441_valid_1 <= _GEN_8094;
        end
      end else begin
        meta_441_valid_1 <= _GEN_3006;
      end
    end else begin
      meta_441_valid_1 <= _GEN_3006;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_441_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_441_lru <= _GEN_8677;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_442_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_442_valid_0 <= _GEN_2495;
        end else begin
          meta_442_valid_0 <= _GEN_8095;
        end
      end else begin
        meta_442_valid_0 <= _GEN_2495;
      end
    end else begin
      meta_442_valid_0 <= _GEN_2495;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_442_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_442_valid_1 <= _GEN_3007;
        end else begin
          meta_442_valid_1 <= _GEN_8096;
        end
      end else begin
        meta_442_valid_1 <= _GEN_3007;
      end
    end else begin
      meta_442_valid_1 <= _GEN_3007;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_442_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_442_lru <= _GEN_8678;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_443_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_443_valid_0 <= _GEN_2496;
        end else begin
          meta_443_valid_0 <= _GEN_8097;
        end
      end else begin
        meta_443_valid_0 <= _GEN_2496;
      end
    end else begin
      meta_443_valid_0 <= _GEN_2496;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_443_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_443_valid_1 <= _GEN_3008;
        end else begin
          meta_443_valid_1 <= _GEN_8098;
        end
      end else begin
        meta_443_valid_1 <= _GEN_3008;
      end
    end else begin
      meta_443_valid_1 <= _GEN_3008;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_443_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_443_lru <= _GEN_8679;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_444_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_444_valid_0 <= _GEN_2497;
        end else begin
          meta_444_valid_0 <= _GEN_8099;
        end
      end else begin
        meta_444_valid_0 <= _GEN_2497;
      end
    end else begin
      meta_444_valid_0 <= _GEN_2497;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_444_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_444_valid_1 <= _GEN_3009;
        end else begin
          meta_444_valid_1 <= _GEN_8100;
        end
      end else begin
        meta_444_valid_1 <= _GEN_3009;
      end
    end else begin
      meta_444_valid_1 <= _GEN_3009;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_444_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_444_lru <= _GEN_8680;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_445_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_445_valid_0 <= _GEN_2498;
        end else begin
          meta_445_valid_0 <= _GEN_8101;
        end
      end else begin
        meta_445_valid_0 <= _GEN_2498;
      end
    end else begin
      meta_445_valid_0 <= _GEN_2498;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_445_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_445_valid_1 <= _GEN_3010;
        end else begin
          meta_445_valid_1 <= _GEN_8102;
        end
      end else begin
        meta_445_valid_1 <= _GEN_3010;
      end
    end else begin
      meta_445_valid_1 <= _GEN_3010;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_445_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_445_lru <= _GEN_8681;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_446_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_446_valid_0 <= _GEN_2499;
        end else begin
          meta_446_valid_0 <= _GEN_8103;
        end
      end else begin
        meta_446_valid_0 <= _GEN_2499;
      end
    end else begin
      meta_446_valid_0 <= _GEN_2499;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_446_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_446_valid_1 <= _GEN_3011;
        end else begin
          meta_446_valid_1 <= _GEN_8104;
        end
      end else begin
        meta_446_valid_1 <= _GEN_3011;
      end
    end else begin
      meta_446_valid_1 <= _GEN_3011;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_446_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_446_lru <= _GEN_8682;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_447_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_447_valid_0 <= _GEN_2500;
        end else begin
          meta_447_valid_0 <= _GEN_8105;
        end
      end else begin
        meta_447_valid_0 <= _GEN_2500;
      end
    end else begin
      meta_447_valid_0 <= _GEN_2500;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_447_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_447_valid_1 <= _GEN_3012;
        end else begin
          meta_447_valid_1 <= _GEN_8106;
        end
      end else begin
        meta_447_valid_1 <= _GEN_3012;
      end
    end else begin
      meta_447_valid_1 <= _GEN_3012;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_447_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_447_lru <= _GEN_8683;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_448_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_448_valid_0 <= _GEN_2501;
        end else begin
          meta_448_valid_0 <= _GEN_8107;
        end
      end else begin
        meta_448_valid_0 <= _GEN_2501;
      end
    end else begin
      meta_448_valid_0 <= _GEN_2501;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_448_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_448_valid_1 <= _GEN_3013;
        end else begin
          meta_448_valid_1 <= _GEN_8108;
        end
      end else begin
        meta_448_valid_1 <= _GEN_3013;
      end
    end else begin
      meta_448_valid_1 <= _GEN_3013;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_448_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_448_lru <= _GEN_8684;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_449_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_449_valid_0 <= _GEN_2502;
        end else begin
          meta_449_valid_0 <= _GEN_8109;
        end
      end else begin
        meta_449_valid_0 <= _GEN_2502;
      end
    end else begin
      meta_449_valid_0 <= _GEN_2502;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_449_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_449_valid_1 <= _GEN_3014;
        end else begin
          meta_449_valid_1 <= _GEN_8110;
        end
      end else begin
        meta_449_valid_1 <= _GEN_3014;
      end
    end else begin
      meta_449_valid_1 <= _GEN_3014;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_449_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_449_lru <= _GEN_8685;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_450_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_450_valid_0 <= _GEN_2503;
        end else begin
          meta_450_valid_0 <= _GEN_8111;
        end
      end else begin
        meta_450_valid_0 <= _GEN_2503;
      end
    end else begin
      meta_450_valid_0 <= _GEN_2503;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_450_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_450_valid_1 <= _GEN_3015;
        end else begin
          meta_450_valid_1 <= _GEN_8112;
        end
      end else begin
        meta_450_valid_1 <= _GEN_3015;
      end
    end else begin
      meta_450_valid_1 <= _GEN_3015;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_450_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_450_lru <= _GEN_8686;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_451_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_451_valid_0 <= _GEN_2504;
        end else begin
          meta_451_valid_0 <= _GEN_8113;
        end
      end else begin
        meta_451_valid_0 <= _GEN_2504;
      end
    end else begin
      meta_451_valid_0 <= _GEN_2504;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_451_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_451_valid_1 <= _GEN_3016;
        end else begin
          meta_451_valid_1 <= _GEN_8114;
        end
      end else begin
        meta_451_valid_1 <= _GEN_3016;
      end
    end else begin
      meta_451_valid_1 <= _GEN_3016;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_451_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_451_lru <= _GEN_8687;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_452_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_452_valid_0 <= _GEN_2505;
        end else begin
          meta_452_valid_0 <= _GEN_8115;
        end
      end else begin
        meta_452_valid_0 <= _GEN_2505;
      end
    end else begin
      meta_452_valid_0 <= _GEN_2505;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_452_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_452_valid_1 <= _GEN_3017;
        end else begin
          meta_452_valid_1 <= _GEN_8116;
        end
      end else begin
        meta_452_valid_1 <= _GEN_3017;
      end
    end else begin
      meta_452_valid_1 <= _GEN_3017;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_452_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_452_lru <= _GEN_8688;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_453_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_453_valid_0 <= _GEN_2506;
        end else begin
          meta_453_valid_0 <= _GEN_8117;
        end
      end else begin
        meta_453_valid_0 <= _GEN_2506;
      end
    end else begin
      meta_453_valid_0 <= _GEN_2506;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_453_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_453_valid_1 <= _GEN_3018;
        end else begin
          meta_453_valid_1 <= _GEN_8118;
        end
      end else begin
        meta_453_valid_1 <= _GEN_3018;
      end
    end else begin
      meta_453_valid_1 <= _GEN_3018;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_453_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_453_lru <= _GEN_8689;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_454_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_454_valid_0 <= _GEN_2507;
        end else begin
          meta_454_valid_0 <= _GEN_8119;
        end
      end else begin
        meta_454_valid_0 <= _GEN_2507;
      end
    end else begin
      meta_454_valid_0 <= _GEN_2507;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_454_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_454_valid_1 <= _GEN_3019;
        end else begin
          meta_454_valid_1 <= _GEN_8120;
        end
      end else begin
        meta_454_valid_1 <= _GEN_3019;
      end
    end else begin
      meta_454_valid_1 <= _GEN_3019;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_454_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_454_lru <= _GEN_8690;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_455_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_455_valid_0 <= _GEN_2508;
        end else begin
          meta_455_valid_0 <= _GEN_8121;
        end
      end else begin
        meta_455_valid_0 <= _GEN_2508;
      end
    end else begin
      meta_455_valid_0 <= _GEN_2508;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_455_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_455_valid_1 <= _GEN_3020;
        end else begin
          meta_455_valid_1 <= _GEN_8122;
        end
      end else begin
        meta_455_valid_1 <= _GEN_3020;
      end
    end else begin
      meta_455_valid_1 <= _GEN_3020;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_455_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_455_lru <= _GEN_8691;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_456_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_456_valid_0 <= _GEN_2509;
        end else begin
          meta_456_valid_0 <= _GEN_8123;
        end
      end else begin
        meta_456_valid_0 <= _GEN_2509;
      end
    end else begin
      meta_456_valid_0 <= _GEN_2509;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_456_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_456_valid_1 <= _GEN_3021;
        end else begin
          meta_456_valid_1 <= _GEN_8124;
        end
      end else begin
        meta_456_valid_1 <= _GEN_3021;
      end
    end else begin
      meta_456_valid_1 <= _GEN_3021;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_456_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_456_lru <= _GEN_8692;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_457_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_457_valid_0 <= _GEN_2510;
        end else begin
          meta_457_valid_0 <= _GEN_8125;
        end
      end else begin
        meta_457_valid_0 <= _GEN_2510;
      end
    end else begin
      meta_457_valid_0 <= _GEN_2510;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_457_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_457_valid_1 <= _GEN_3022;
        end else begin
          meta_457_valid_1 <= _GEN_8126;
        end
      end else begin
        meta_457_valid_1 <= _GEN_3022;
      end
    end else begin
      meta_457_valid_1 <= _GEN_3022;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_457_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_457_lru <= _GEN_8693;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_458_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_458_valid_0 <= _GEN_2511;
        end else begin
          meta_458_valid_0 <= _GEN_8127;
        end
      end else begin
        meta_458_valid_0 <= _GEN_2511;
      end
    end else begin
      meta_458_valid_0 <= _GEN_2511;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_458_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_458_valid_1 <= _GEN_3023;
        end else begin
          meta_458_valid_1 <= _GEN_8128;
        end
      end else begin
        meta_458_valid_1 <= _GEN_3023;
      end
    end else begin
      meta_458_valid_1 <= _GEN_3023;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_458_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_458_lru <= _GEN_8694;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_459_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_459_valid_0 <= _GEN_2512;
        end else begin
          meta_459_valid_0 <= _GEN_8129;
        end
      end else begin
        meta_459_valid_0 <= _GEN_2512;
      end
    end else begin
      meta_459_valid_0 <= _GEN_2512;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_459_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_459_valid_1 <= _GEN_3024;
        end else begin
          meta_459_valid_1 <= _GEN_8130;
        end
      end else begin
        meta_459_valid_1 <= _GEN_3024;
      end
    end else begin
      meta_459_valid_1 <= _GEN_3024;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_459_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_459_lru <= _GEN_8695;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_460_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_460_valid_0 <= _GEN_2513;
        end else begin
          meta_460_valid_0 <= _GEN_8131;
        end
      end else begin
        meta_460_valid_0 <= _GEN_2513;
      end
    end else begin
      meta_460_valid_0 <= _GEN_2513;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_460_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_460_valid_1 <= _GEN_3025;
        end else begin
          meta_460_valid_1 <= _GEN_8132;
        end
      end else begin
        meta_460_valid_1 <= _GEN_3025;
      end
    end else begin
      meta_460_valid_1 <= _GEN_3025;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_460_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_460_lru <= _GEN_8696;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_461_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_461_valid_0 <= _GEN_2514;
        end else begin
          meta_461_valid_0 <= _GEN_8133;
        end
      end else begin
        meta_461_valid_0 <= _GEN_2514;
      end
    end else begin
      meta_461_valid_0 <= _GEN_2514;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_461_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_461_valid_1 <= _GEN_3026;
        end else begin
          meta_461_valid_1 <= _GEN_8134;
        end
      end else begin
        meta_461_valid_1 <= _GEN_3026;
      end
    end else begin
      meta_461_valid_1 <= _GEN_3026;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_461_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_461_lru <= _GEN_8697;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_462_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_462_valid_0 <= _GEN_2515;
        end else begin
          meta_462_valid_0 <= _GEN_8135;
        end
      end else begin
        meta_462_valid_0 <= _GEN_2515;
      end
    end else begin
      meta_462_valid_0 <= _GEN_2515;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_462_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_462_valid_1 <= _GEN_3027;
        end else begin
          meta_462_valid_1 <= _GEN_8136;
        end
      end else begin
        meta_462_valid_1 <= _GEN_3027;
      end
    end else begin
      meta_462_valid_1 <= _GEN_3027;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_462_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_462_lru <= _GEN_8698;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_463_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_463_valid_0 <= _GEN_2516;
        end else begin
          meta_463_valid_0 <= _GEN_8137;
        end
      end else begin
        meta_463_valid_0 <= _GEN_2516;
      end
    end else begin
      meta_463_valid_0 <= _GEN_2516;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_463_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_463_valid_1 <= _GEN_3028;
        end else begin
          meta_463_valid_1 <= _GEN_8138;
        end
      end else begin
        meta_463_valid_1 <= _GEN_3028;
      end
    end else begin
      meta_463_valid_1 <= _GEN_3028;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_463_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_463_lru <= _GEN_8699;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_464_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_464_valid_0 <= _GEN_2517;
        end else begin
          meta_464_valid_0 <= _GEN_8139;
        end
      end else begin
        meta_464_valid_0 <= _GEN_2517;
      end
    end else begin
      meta_464_valid_0 <= _GEN_2517;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_464_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_464_valid_1 <= _GEN_3029;
        end else begin
          meta_464_valid_1 <= _GEN_8140;
        end
      end else begin
        meta_464_valid_1 <= _GEN_3029;
      end
    end else begin
      meta_464_valid_1 <= _GEN_3029;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_464_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_464_lru <= _GEN_8700;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_465_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_465_valid_0 <= _GEN_2518;
        end else begin
          meta_465_valid_0 <= _GEN_8141;
        end
      end else begin
        meta_465_valid_0 <= _GEN_2518;
      end
    end else begin
      meta_465_valid_0 <= _GEN_2518;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_465_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_465_valid_1 <= _GEN_3030;
        end else begin
          meta_465_valid_1 <= _GEN_8142;
        end
      end else begin
        meta_465_valid_1 <= _GEN_3030;
      end
    end else begin
      meta_465_valid_1 <= _GEN_3030;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_465_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_465_lru <= _GEN_8701;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_466_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_466_valid_0 <= _GEN_2519;
        end else begin
          meta_466_valid_0 <= _GEN_8143;
        end
      end else begin
        meta_466_valid_0 <= _GEN_2519;
      end
    end else begin
      meta_466_valid_0 <= _GEN_2519;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_466_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_466_valid_1 <= _GEN_3031;
        end else begin
          meta_466_valid_1 <= _GEN_8144;
        end
      end else begin
        meta_466_valid_1 <= _GEN_3031;
      end
    end else begin
      meta_466_valid_1 <= _GEN_3031;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_466_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_466_lru <= _GEN_8702;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_467_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_467_valid_0 <= _GEN_2520;
        end else begin
          meta_467_valid_0 <= _GEN_8145;
        end
      end else begin
        meta_467_valid_0 <= _GEN_2520;
      end
    end else begin
      meta_467_valid_0 <= _GEN_2520;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_467_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_467_valid_1 <= _GEN_3032;
        end else begin
          meta_467_valid_1 <= _GEN_8146;
        end
      end else begin
        meta_467_valid_1 <= _GEN_3032;
      end
    end else begin
      meta_467_valid_1 <= _GEN_3032;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_467_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_467_lru <= _GEN_8703;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_468_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_468_valid_0 <= _GEN_2521;
        end else begin
          meta_468_valid_0 <= _GEN_8147;
        end
      end else begin
        meta_468_valid_0 <= _GEN_2521;
      end
    end else begin
      meta_468_valid_0 <= _GEN_2521;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_468_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_468_valid_1 <= _GEN_3033;
        end else begin
          meta_468_valid_1 <= _GEN_8148;
        end
      end else begin
        meta_468_valid_1 <= _GEN_3033;
      end
    end else begin
      meta_468_valid_1 <= _GEN_3033;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_468_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_468_lru <= _GEN_8704;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_469_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_469_valid_0 <= _GEN_2522;
        end else begin
          meta_469_valid_0 <= _GEN_8149;
        end
      end else begin
        meta_469_valid_0 <= _GEN_2522;
      end
    end else begin
      meta_469_valid_0 <= _GEN_2522;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_469_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_469_valid_1 <= _GEN_3034;
        end else begin
          meta_469_valid_1 <= _GEN_8150;
        end
      end else begin
        meta_469_valid_1 <= _GEN_3034;
      end
    end else begin
      meta_469_valid_1 <= _GEN_3034;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_469_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_469_lru <= _GEN_8705;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_470_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_470_valid_0 <= _GEN_2523;
        end else begin
          meta_470_valid_0 <= _GEN_8151;
        end
      end else begin
        meta_470_valid_0 <= _GEN_2523;
      end
    end else begin
      meta_470_valid_0 <= _GEN_2523;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_470_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_470_valid_1 <= _GEN_3035;
        end else begin
          meta_470_valid_1 <= _GEN_8152;
        end
      end else begin
        meta_470_valid_1 <= _GEN_3035;
      end
    end else begin
      meta_470_valid_1 <= _GEN_3035;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_470_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_470_lru <= _GEN_8706;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_471_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_471_valid_0 <= _GEN_2524;
        end else begin
          meta_471_valid_0 <= _GEN_8153;
        end
      end else begin
        meta_471_valid_0 <= _GEN_2524;
      end
    end else begin
      meta_471_valid_0 <= _GEN_2524;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_471_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_471_valid_1 <= _GEN_3036;
        end else begin
          meta_471_valid_1 <= _GEN_8154;
        end
      end else begin
        meta_471_valid_1 <= _GEN_3036;
      end
    end else begin
      meta_471_valid_1 <= _GEN_3036;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_471_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_471_lru <= _GEN_8707;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_472_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_472_valid_0 <= _GEN_2525;
        end else begin
          meta_472_valid_0 <= _GEN_8155;
        end
      end else begin
        meta_472_valid_0 <= _GEN_2525;
      end
    end else begin
      meta_472_valid_0 <= _GEN_2525;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_472_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_472_valid_1 <= _GEN_3037;
        end else begin
          meta_472_valid_1 <= _GEN_8156;
        end
      end else begin
        meta_472_valid_1 <= _GEN_3037;
      end
    end else begin
      meta_472_valid_1 <= _GEN_3037;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_472_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_472_lru <= _GEN_8708;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_473_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_473_valid_0 <= _GEN_2526;
        end else begin
          meta_473_valid_0 <= _GEN_8157;
        end
      end else begin
        meta_473_valid_0 <= _GEN_2526;
      end
    end else begin
      meta_473_valid_0 <= _GEN_2526;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_473_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_473_valid_1 <= _GEN_3038;
        end else begin
          meta_473_valid_1 <= _GEN_8158;
        end
      end else begin
        meta_473_valid_1 <= _GEN_3038;
      end
    end else begin
      meta_473_valid_1 <= _GEN_3038;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_473_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_473_lru <= _GEN_8709;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_474_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_474_valid_0 <= _GEN_2527;
        end else begin
          meta_474_valid_0 <= _GEN_8159;
        end
      end else begin
        meta_474_valid_0 <= _GEN_2527;
      end
    end else begin
      meta_474_valid_0 <= _GEN_2527;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_474_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_474_valid_1 <= _GEN_3039;
        end else begin
          meta_474_valid_1 <= _GEN_8160;
        end
      end else begin
        meta_474_valid_1 <= _GEN_3039;
      end
    end else begin
      meta_474_valid_1 <= _GEN_3039;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_474_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_474_lru <= _GEN_8710;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_475_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_475_valid_0 <= _GEN_2528;
        end else begin
          meta_475_valid_0 <= _GEN_8161;
        end
      end else begin
        meta_475_valid_0 <= _GEN_2528;
      end
    end else begin
      meta_475_valid_0 <= _GEN_2528;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_475_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_475_valid_1 <= _GEN_3040;
        end else begin
          meta_475_valid_1 <= _GEN_8162;
        end
      end else begin
        meta_475_valid_1 <= _GEN_3040;
      end
    end else begin
      meta_475_valid_1 <= _GEN_3040;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_475_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_475_lru <= _GEN_8711;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_476_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_476_valid_0 <= _GEN_2529;
        end else begin
          meta_476_valid_0 <= _GEN_8163;
        end
      end else begin
        meta_476_valid_0 <= _GEN_2529;
      end
    end else begin
      meta_476_valid_0 <= _GEN_2529;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_476_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_476_valid_1 <= _GEN_3041;
        end else begin
          meta_476_valid_1 <= _GEN_8164;
        end
      end else begin
        meta_476_valid_1 <= _GEN_3041;
      end
    end else begin
      meta_476_valid_1 <= _GEN_3041;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_476_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_476_lru <= _GEN_8712;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_477_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_477_valid_0 <= _GEN_2530;
        end else begin
          meta_477_valid_0 <= _GEN_8165;
        end
      end else begin
        meta_477_valid_0 <= _GEN_2530;
      end
    end else begin
      meta_477_valid_0 <= _GEN_2530;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_477_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_477_valid_1 <= _GEN_3042;
        end else begin
          meta_477_valid_1 <= _GEN_8166;
        end
      end else begin
        meta_477_valid_1 <= _GEN_3042;
      end
    end else begin
      meta_477_valid_1 <= _GEN_3042;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_477_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_477_lru <= _GEN_8713;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_478_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_478_valid_0 <= _GEN_2531;
        end else begin
          meta_478_valid_0 <= _GEN_8167;
        end
      end else begin
        meta_478_valid_0 <= _GEN_2531;
      end
    end else begin
      meta_478_valid_0 <= _GEN_2531;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_478_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_478_valid_1 <= _GEN_3043;
        end else begin
          meta_478_valid_1 <= _GEN_8168;
        end
      end else begin
        meta_478_valid_1 <= _GEN_3043;
      end
    end else begin
      meta_478_valid_1 <= _GEN_3043;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_478_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_478_lru <= _GEN_8714;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_479_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_479_valid_0 <= _GEN_2532;
        end else begin
          meta_479_valid_0 <= _GEN_8169;
        end
      end else begin
        meta_479_valid_0 <= _GEN_2532;
      end
    end else begin
      meta_479_valid_0 <= _GEN_2532;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_479_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_479_valid_1 <= _GEN_3044;
        end else begin
          meta_479_valid_1 <= _GEN_8170;
        end
      end else begin
        meta_479_valid_1 <= _GEN_3044;
      end
    end else begin
      meta_479_valid_1 <= _GEN_3044;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_479_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_479_lru <= _GEN_8715;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_480_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_480_valid_0 <= _GEN_2533;
        end else begin
          meta_480_valid_0 <= _GEN_8171;
        end
      end else begin
        meta_480_valid_0 <= _GEN_2533;
      end
    end else begin
      meta_480_valid_0 <= _GEN_2533;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_480_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_480_valid_1 <= _GEN_3045;
        end else begin
          meta_480_valid_1 <= _GEN_8172;
        end
      end else begin
        meta_480_valid_1 <= _GEN_3045;
      end
    end else begin
      meta_480_valid_1 <= _GEN_3045;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_480_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_480_lru <= _GEN_8716;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_481_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_481_valid_0 <= _GEN_2534;
        end else begin
          meta_481_valid_0 <= _GEN_8173;
        end
      end else begin
        meta_481_valid_0 <= _GEN_2534;
      end
    end else begin
      meta_481_valid_0 <= _GEN_2534;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_481_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_481_valid_1 <= _GEN_3046;
        end else begin
          meta_481_valid_1 <= _GEN_8174;
        end
      end else begin
        meta_481_valid_1 <= _GEN_3046;
      end
    end else begin
      meta_481_valid_1 <= _GEN_3046;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_481_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_481_lru <= _GEN_8717;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_482_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_482_valid_0 <= _GEN_2535;
        end else begin
          meta_482_valid_0 <= _GEN_8175;
        end
      end else begin
        meta_482_valid_0 <= _GEN_2535;
      end
    end else begin
      meta_482_valid_0 <= _GEN_2535;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_482_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_482_valid_1 <= _GEN_3047;
        end else begin
          meta_482_valid_1 <= _GEN_8176;
        end
      end else begin
        meta_482_valid_1 <= _GEN_3047;
      end
    end else begin
      meta_482_valid_1 <= _GEN_3047;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_482_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_482_lru <= _GEN_8718;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_483_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_483_valid_0 <= _GEN_2536;
        end else begin
          meta_483_valid_0 <= _GEN_8177;
        end
      end else begin
        meta_483_valid_0 <= _GEN_2536;
      end
    end else begin
      meta_483_valid_0 <= _GEN_2536;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_483_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_483_valid_1 <= _GEN_3048;
        end else begin
          meta_483_valid_1 <= _GEN_8178;
        end
      end else begin
        meta_483_valid_1 <= _GEN_3048;
      end
    end else begin
      meta_483_valid_1 <= _GEN_3048;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_483_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_483_lru <= _GEN_8719;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_484_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_484_valid_0 <= _GEN_2537;
        end else begin
          meta_484_valid_0 <= _GEN_8179;
        end
      end else begin
        meta_484_valid_0 <= _GEN_2537;
      end
    end else begin
      meta_484_valid_0 <= _GEN_2537;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_484_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_484_valid_1 <= _GEN_3049;
        end else begin
          meta_484_valid_1 <= _GEN_8180;
        end
      end else begin
        meta_484_valid_1 <= _GEN_3049;
      end
    end else begin
      meta_484_valid_1 <= _GEN_3049;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_484_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_484_lru <= _GEN_8720;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_485_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_485_valid_0 <= _GEN_2538;
        end else begin
          meta_485_valid_0 <= _GEN_8181;
        end
      end else begin
        meta_485_valid_0 <= _GEN_2538;
      end
    end else begin
      meta_485_valid_0 <= _GEN_2538;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_485_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_485_valid_1 <= _GEN_3050;
        end else begin
          meta_485_valid_1 <= _GEN_8182;
        end
      end else begin
        meta_485_valid_1 <= _GEN_3050;
      end
    end else begin
      meta_485_valid_1 <= _GEN_3050;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_485_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_485_lru <= _GEN_8721;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_486_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_486_valid_0 <= _GEN_2539;
        end else begin
          meta_486_valid_0 <= _GEN_8183;
        end
      end else begin
        meta_486_valid_0 <= _GEN_2539;
      end
    end else begin
      meta_486_valid_0 <= _GEN_2539;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_486_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_486_valid_1 <= _GEN_3051;
        end else begin
          meta_486_valid_1 <= _GEN_8184;
        end
      end else begin
        meta_486_valid_1 <= _GEN_3051;
      end
    end else begin
      meta_486_valid_1 <= _GEN_3051;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_486_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_486_lru <= _GEN_8722;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_487_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_487_valid_0 <= _GEN_2540;
        end else begin
          meta_487_valid_0 <= _GEN_8185;
        end
      end else begin
        meta_487_valid_0 <= _GEN_2540;
      end
    end else begin
      meta_487_valid_0 <= _GEN_2540;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_487_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_487_valid_1 <= _GEN_3052;
        end else begin
          meta_487_valid_1 <= _GEN_8186;
        end
      end else begin
        meta_487_valid_1 <= _GEN_3052;
      end
    end else begin
      meta_487_valid_1 <= _GEN_3052;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_487_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_487_lru <= _GEN_8723;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_488_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_488_valid_0 <= _GEN_2541;
        end else begin
          meta_488_valid_0 <= _GEN_8187;
        end
      end else begin
        meta_488_valid_0 <= _GEN_2541;
      end
    end else begin
      meta_488_valid_0 <= _GEN_2541;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_488_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_488_valid_1 <= _GEN_3053;
        end else begin
          meta_488_valid_1 <= _GEN_8188;
        end
      end else begin
        meta_488_valid_1 <= _GEN_3053;
      end
    end else begin
      meta_488_valid_1 <= _GEN_3053;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_488_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_488_lru <= _GEN_8724;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_489_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_489_valid_0 <= _GEN_2542;
        end else begin
          meta_489_valid_0 <= _GEN_8189;
        end
      end else begin
        meta_489_valid_0 <= _GEN_2542;
      end
    end else begin
      meta_489_valid_0 <= _GEN_2542;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_489_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_489_valid_1 <= _GEN_3054;
        end else begin
          meta_489_valid_1 <= _GEN_8190;
        end
      end else begin
        meta_489_valid_1 <= _GEN_3054;
      end
    end else begin
      meta_489_valid_1 <= _GEN_3054;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_489_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_489_lru <= _GEN_8725;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_490_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_490_valid_0 <= _GEN_2543;
        end else begin
          meta_490_valid_0 <= _GEN_8191;
        end
      end else begin
        meta_490_valid_0 <= _GEN_2543;
      end
    end else begin
      meta_490_valid_0 <= _GEN_2543;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_490_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_490_valid_1 <= _GEN_3055;
        end else begin
          meta_490_valid_1 <= _GEN_8192;
        end
      end else begin
        meta_490_valid_1 <= _GEN_3055;
      end
    end else begin
      meta_490_valid_1 <= _GEN_3055;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_490_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_490_lru <= _GEN_8726;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_491_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_491_valid_0 <= _GEN_2544;
        end else begin
          meta_491_valid_0 <= _GEN_8193;
        end
      end else begin
        meta_491_valid_0 <= _GEN_2544;
      end
    end else begin
      meta_491_valid_0 <= _GEN_2544;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_491_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_491_valid_1 <= _GEN_3056;
        end else begin
          meta_491_valid_1 <= _GEN_8194;
        end
      end else begin
        meta_491_valid_1 <= _GEN_3056;
      end
    end else begin
      meta_491_valid_1 <= _GEN_3056;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_491_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_491_lru <= _GEN_8727;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_492_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_492_valid_0 <= _GEN_2545;
        end else begin
          meta_492_valid_0 <= _GEN_8195;
        end
      end else begin
        meta_492_valid_0 <= _GEN_2545;
      end
    end else begin
      meta_492_valid_0 <= _GEN_2545;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_492_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_492_valid_1 <= _GEN_3057;
        end else begin
          meta_492_valid_1 <= _GEN_8196;
        end
      end else begin
        meta_492_valid_1 <= _GEN_3057;
      end
    end else begin
      meta_492_valid_1 <= _GEN_3057;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_492_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_492_lru <= _GEN_8728;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_493_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_493_valid_0 <= _GEN_2546;
        end else begin
          meta_493_valid_0 <= _GEN_8197;
        end
      end else begin
        meta_493_valid_0 <= _GEN_2546;
      end
    end else begin
      meta_493_valid_0 <= _GEN_2546;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_493_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_493_valid_1 <= _GEN_3058;
        end else begin
          meta_493_valid_1 <= _GEN_8198;
        end
      end else begin
        meta_493_valid_1 <= _GEN_3058;
      end
    end else begin
      meta_493_valid_1 <= _GEN_3058;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_493_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_493_lru <= _GEN_8729;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_494_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_494_valid_0 <= _GEN_2547;
        end else begin
          meta_494_valid_0 <= _GEN_8199;
        end
      end else begin
        meta_494_valid_0 <= _GEN_2547;
      end
    end else begin
      meta_494_valid_0 <= _GEN_2547;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_494_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_494_valid_1 <= _GEN_3059;
        end else begin
          meta_494_valid_1 <= _GEN_8200;
        end
      end else begin
        meta_494_valid_1 <= _GEN_3059;
      end
    end else begin
      meta_494_valid_1 <= _GEN_3059;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_494_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_494_lru <= _GEN_8730;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_495_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_495_valid_0 <= _GEN_2548;
        end else begin
          meta_495_valid_0 <= _GEN_8201;
        end
      end else begin
        meta_495_valid_0 <= _GEN_2548;
      end
    end else begin
      meta_495_valid_0 <= _GEN_2548;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_495_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_495_valid_1 <= _GEN_3060;
        end else begin
          meta_495_valid_1 <= _GEN_8202;
        end
      end else begin
        meta_495_valid_1 <= _GEN_3060;
      end
    end else begin
      meta_495_valid_1 <= _GEN_3060;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_495_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_495_lru <= _GEN_8731;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_496_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_496_valid_0 <= _GEN_2549;
        end else begin
          meta_496_valid_0 <= _GEN_8203;
        end
      end else begin
        meta_496_valid_0 <= _GEN_2549;
      end
    end else begin
      meta_496_valid_0 <= _GEN_2549;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_496_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_496_valid_1 <= _GEN_3061;
        end else begin
          meta_496_valid_1 <= _GEN_8204;
        end
      end else begin
        meta_496_valid_1 <= _GEN_3061;
      end
    end else begin
      meta_496_valid_1 <= _GEN_3061;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_496_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_496_lru <= _GEN_8732;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_497_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_497_valid_0 <= _GEN_2550;
        end else begin
          meta_497_valid_0 <= _GEN_8205;
        end
      end else begin
        meta_497_valid_0 <= _GEN_2550;
      end
    end else begin
      meta_497_valid_0 <= _GEN_2550;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_497_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_497_valid_1 <= _GEN_3062;
        end else begin
          meta_497_valid_1 <= _GEN_8206;
        end
      end else begin
        meta_497_valid_1 <= _GEN_3062;
      end
    end else begin
      meta_497_valid_1 <= _GEN_3062;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_497_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_497_lru <= _GEN_8733;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_498_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_498_valid_0 <= _GEN_2551;
        end else begin
          meta_498_valid_0 <= _GEN_8207;
        end
      end else begin
        meta_498_valid_0 <= _GEN_2551;
      end
    end else begin
      meta_498_valid_0 <= _GEN_2551;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_498_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_498_valid_1 <= _GEN_3063;
        end else begin
          meta_498_valid_1 <= _GEN_8208;
        end
      end else begin
        meta_498_valid_1 <= _GEN_3063;
      end
    end else begin
      meta_498_valid_1 <= _GEN_3063;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_498_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_498_lru <= _GEN_8734;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_499_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_499_valid_0 <= _GEN_2552;
        end else begin
          meta_499_valid_0 <= _GEN_8209;
        end
      end else begin
        meta_499_valid_0 <= _GEN_2552;
      end
    end else begin
      meta_499_valid_0 <= _GEN_2552;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_499_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_499_valid_1 <= _GEN_3064;
        end else begin
          meta_499_valid_1 <= _GEN_8210;
        end
      end else begin
        meta_499_valid_1 <= _GEN_3064;
      end
    end else begin
      meta_499_valid_1 <= _GEN_3064;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_499_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_499_lru <= _GEN_8735;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_500_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_500_valid_0 <= _GEN_2553;
        end else begin
          meta_500_valid_0 <= _GEN_8211;
        end
      end else begin
        meta_500_valid_0 <= _GEN_2553;
      end
    end else begin
      meta_500_valid_0 <= _GEN_2553;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_500_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_500_valid_1 <= _GEN_3065;
        end else begin
          meta_500_valid_1 <= _GEN_8212;
        end
      end else begin
        meta_500_valid_1 <= _GEN_3065;
      end
    end else begin
      meta_500_valid_1 <= _GEN_3065;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_500_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_500_lru <= _GEN_8736;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_501_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_501_valid_0 <= _GEN_2554;
        end else begin
          meta_501_valid_0 <= _GEN_8213;
        end
      end else begin
        meta_501_valid_0 <= _GEN_2554;
      end
    end else begin
      meta_501_valid_0 <= _GEN_2554;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_501_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_501_valid_1 <= _GEN_3066;
        end else begin
          meta_501_valid_1 <= _GEN_8214;
        end
      end else begin
        meta_501_valid_1 <= _GEN_3066;
      end
    end else begin
      meta_501_valid_1 <= _GEN_3066;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_501_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_501_lru <= _GEN_8737;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_502_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_502_valid_0 <= _GEN_2555;
        end else begin
          meta_502_valid_0 <= _GEN_8215;
        end
      end else begin
        meta_502_valid_0 <= _GEN_2555;
      end
    end else begin
      meta_502_valid_0 <= _GEN_2555;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_502_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_502_valid_1 <= _GEN_3067;
        end else begin
          meta_502_valid_1 <= _GEN_8216;
        end
      end else begin
        meta_502_valid_1 <= _GEN_3067;
      end
    end else begin
      meta_502_valid_1 <= _GEN_3067;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_502_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_502_lru <= _GEN_8738;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_503_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_503_valid_0 <= _GEN_2556;
        end else begin
          meta_503_valid_0 <= _GEN_8217;
        end
      end else begin
        meta_503_valid_0 <= _GEN_2556;
      end
    end else begin
      meta_503_valid_0 <= _GEN_2556;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_503_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_503_valid_1 <= _GEN_3068;
        end else begin
          meta_503_valid_1 <= _GEN_8218;
        end
      end else begin
        meta_503_valid_1 <= _GEN_3068;
      end
    end else begin
      meta_503_valid_1 <= _GEN_3068;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_503_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_503_lru <= _GEN_8739;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_504_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_504_valid_0 <= _GEN_2557;
        end else begin
          meta_504_valid_0 <= _GEN_8219;
        end
      end else begin
        meta_504_valid_0 <= _GEN_2557;
      end
    end else begin
      meta_504_valid_0 <= _GEN_2557;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_504_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_504_valid_1 <= _GEN_3069;
        end else begin
          meta_504_valid_1 <= _GEN_8220;
        end
      end else begin
        meta_504_valid_1 <= _GEN_3069;
      end
    end else begin
      meta_504_valid_1 <= _GEN_3069;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_504_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_504_lru <= _GEN_8740;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_505_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_505_valid_0 <= _GEN_2558;
        end else begin
          meta_505_valid_0 <= _GEN_8221;
        end
      end else begin
        meta_505_valid_0 <= _GEN_2558;
      end
    end else begin
      meta_505_valid_0 <= _GEN_2558;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_505_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_505_valid_1 <= _GEN_3070;
        end else begin
          meta_505_valid_1 <= _GEN_8222;
        end
      end else begin
        meta_505_valid_1 <= _GEN_3070;
      end
    end else begin
      meta_505_valid_1 <= _GEN_3070;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_505_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_505_lru <= _GEN_8741;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_506_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_506_valid_0 <= _GEN_2559;
        end else begin
          meta_506_valid_0 <= _GEN_8223;
        end
      end else begin
        meta_506_valid_0 <= _GEN_2559;
      end
    end else begin
      meta_506_valid_0 <= _GEN_2559;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_506_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_506_valid_1 <= _GEN_3071;
        end else begin
          meta_506_valid_1 <= _GEN_8224;
        end
      end else begin
        meta_506_valid_1 <= _GEN_3071;
      end
    end else begin
      meta_506_valid_1 <= _GEN_3071;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_506_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_506_lru <= _GEN_8742;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_507_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_507_valid_0 <= _GEN_2560;
        end else begin
          meta_507_valid_0 <= _GEN_8225;
        end
      end else begin
        meta_507_valid_0 <= _GEN_2560;
      end
    end else begin
      meta_507_valid_0 <= _GEN_2560;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_507_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_507_valid_1 <= _GEN_3072;
        end else begin
          meta_507_valid_1 <= _GEN_8226;
        end
      end else begin
        meta_507_valid_1 <= _GEN_3072;
      end
    end else begin
      meta_507_valid_1 <= _GEN_3072;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_507_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_507_lru <= _GEN_8743;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_508_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_508_valid_0 <= _GEN_2561;
        end else begin
          meta_508_valid_0 <= _GEN_8227;
        end
      end else begin
        meta_508_valid_0 <= _GEN_2561;
      end
    end else begin
      meta_508_valid_0 <= _GEN_2561;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_508_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_508_valid_1 <= _GEN_3073;
        end else begin
          meta_508_valid_1 <= _GEN_8228;
        end
      end else begin
        meta_508_valid_1 <= _GEN_3073;
      end
    end else begin
      meta_508_valid_1 <= _GEN_3073;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_508_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_508_lru <= _GEN_8744;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_509_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_509_valid_0 <= _GEN_2562;
        end else begin
          meta_509_valid_0 <= _GEN_8229;
        end
      end else begin
        meta_509_valid_0 <= _GEN_2562;
      end
    end else begin
      meta_509_valid_0 <= _GEN_2562;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_509_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_509_valid_1 <= _GEN_3074;
        end else begin
          meta_509_valid_1 <= _GEN_8230;
        end
      end else begin
        meta_509_valid_1 <= _GEN_3074;
      end
    end else begin
      meta_509_valid_1 <= _GEN_3074;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_509_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_509_lru <= _GEN_8745;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_510_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_510_valid_0 <= _GEN_2563;
        end else begin
          meta_510_valid_0 <= _GEN_8231;
        end
      end else begin
        meta_510_valid_0 <= _GEN_2563;
      end
    end else begin
      meta_510_valid_0 <= _GEN_2563;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_510_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_510_valid_1 <= _GEN_3075;
        end else begin
          meta_510_valid_1 <= _GEN_8232;
        end
      end else begin
        meta_510_valid_1 <= _GEN_3075;
      end
    end else begin
      meta_510_valid_1 <= _GEN_3075;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_510_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_510_lru <= _GEN_8746;
        end
      end
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_511_valid_0 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_511_valid_0 <= _GEN_2564;
        end else begin
          meta_511_valid_0 <= _GEN_8233;
        end
      end else begin
        meta_511_valid_0 <= _GEN_2564;
      end
    end else begin
      meta_511_valid_0 <= _GEN_2564;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_511_valid_1 <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          meta_511_valid_1 <= _GEN_3076;
        end else begin
          meta_511_valid_1 <= _GEN_8234;
        end
      end else begin
        meta_511_valid_1 <= _GEN_3076;
      end
    end else begin
      meta_511_valid_1 <= _GEN_3076;
    end
    if (reset) begin // @[ICache.scala 34:21]
      meta_511_lru <= 1'h0; // @[ICache.scala 34:21]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          meta_511_lru <= _GEN_8747;
        end
      end
    end
    tlb_vpn <= _GEN_19663[16:0]; // @[ICache.scala 40:{20,20}]
    tlb_ppn <= _GEN_19664[16:0]; // @[ICache.scala 40:{20,20}]
    if (reset) begin // @[ICache.scala 40:20]
      tlb_uncached <= 1'h0; // @[ICache.scala 40:20]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 163:17]
      if (3'h1 == state) begin // @[ICache.scala 163:17]
        if (_T_19) begin // @[ICache.scala 204:9]
          tlb_uncached <= _tlb_uncached_T_1; // @[ICache.scala 208:22]
        end
      end
    end
    if (reset) begin // @[ICache.scala 40:20]
      tlb_valid <= 1'h0; // @[ICache.scala 40:20]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      tlb_valid <= _GEN_1028;
    end else if (3'h1 == state) begin // @[ICache.scala 163:17]
      tlb_valid <= _GEN_11859;
    end else begin
      tlb_valid <= _GEN_1028;
    end
    if (reset) begin // @[ICache.scala 48:81]
      state <= 3'h0; // @[ICache.scala 48:81]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (~translation_ok) begin // @[ICache.scala 166:31]
          state <= 3'h1; // @[ICache.scala 167:20]
        end else begin
          state <= _GEN_7200;
        end
      end
    end else if (3'h1 == state) begin // @[ICache.scala 163:17]
      if (_T_19) begin // @[ICache.scala 204:9]
        state <= 3'h0; // @[ICache.scala 205:22]
      end else begin
        state <= 3'h4; // @[ICache.scala 211:24]
      end
    end else if (3'h2 == state) begin // @[ICache.scala 163:17]
      state <= _GEN_11871;
    end else begin
      state <= _GEN_11920;
    end
    if (reset) begin // @[ICache.scala 58:38]
      replace_line_addr <= 6'h0; // @[ICache.scala 58:38]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          replace_line_addr <= _GEN_7205;
        end
      end
    end
    if (reset) begin // @[ICache.scala 66:30]
      data_wen_0 <= 8'h0; // @[ICache.scala 66:30]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          data_wen_0 <= _GEN_7206;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 163:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 163:17]
        data_wen_0 <= _GEN_11916;
      end
    end
    if (reset) begin // @[ICache.scala 66:30]
      data_wen_1 <= 8'h0; // @[ICache.scala 66:30]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          data_wen_1 <= _GEN_7207;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 163:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 163:17]
        data_wen_1 <= _GEN_11917;
      end
    end
    if (reset) begin // @[ICache.scala 67:30]
      tag_wen_0 <= 1'h0; // @[ICache.scala 67:30]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          tag_wen_0 <= _GEN_7208;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 163:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 163:17]
        tag_wen_0 <= _GEN_11918;
      end
    end
    if (reset) begin // @[ICache.scala 67:30]
      tag_wen_1 <= 1'h0; // @[ICache.scala 67:30]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          tag_wen_1 <= _GEN_7209;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 163:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 163:17]
        tag_wen_1 <= _GEN_11919;
      end
    end
    tag_ram_wdata <= _GEN_19665[16:0]; // @[ICache.scala 68:{30,30}]
    if (reset) begin // @[ICache.scala 91:22]
      saved_0_inst <= 32'h0; // @[ICache.scala 91:22]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 163:17]
      if (3'h1 == state) begin // @[ICache.scala 163:17]
        if (!(_T_19)) begin // @[ICache.scala 204:9]
          saved_0_inst <= 32'h0; // @[ICache.scala 213:24]
        end
      end else if (3'h2 == state) begin // @[ICache.scala 163:17]
        saved_0_inst <= _GEN_11872;
      end
    end
    if (reset) begin // @[ICache.scala 91:22]
      saved_0_valid <= 1'h0; // @[ICache.scala 91:22]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          saved_0_valid <= _GEN_8749;
        end
      end
    end else if (3'h1 == state) begin // @[ICache.scala 163:17]
      if (!(_T_19)) begin // @[ICache.scala 204:9]
        saved_0_valid <= 1'h1; // @[ICache.scala 214:24]
      end
    end else if (3'h2 == state) begin // @[ICache.scala 163:17]
      saved_0_valid <= _GEN_11873;
    end else begin
      saved_0_valid <= _GEN_11923;
    end
    saved_1_inst <= _GEN_19666[31:0]; // @[ICache.scala 91:{22,22}]
    if (reset) begin // @[ICache.scala 91:22]
      saved_1_valid <= 1'h0; // @[ICache.scala 91:22]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          saved_1_valid <= _GEN_8750;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 163:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 163:17]
        saved_1_valid <= _GEN_11924;
      end
    end
    if (reset) begin // @[ICache.scala 109:24]
      axi_cnt <= 5'h0; // @[ICache.scala 109:24]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          axi_cnt <= _GEN_8235;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 163:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 163:17]
        axi_cnt <= _GEN_11915;
      end
    end
    if (reset) begin // @[ICache.scala 141:24]
      ar_addr <= 32'h0; // @[ICache.scala 141:24]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          ar_addr <= _GEN_7201;
        end
      end
    end
    if (reset) begin // @[ICache.scala 141:24]
      ar_len <= 8'h0; // @[ICache.scala 141:24]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          ar_len <= _GEN_7202;
        end
      end
    end
    if (reset) begin // @[ICache.scala 141:24]
      ar_size <= 3'h0; // @[ICache.scala 141:24]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          ar_size <= _GEN_7203;
        end
      end
    end
    if (reset) begin // @[ICache.scala 142:24]
      arvalid <= 1'h0; // @[ICache.scala 142:24]
    end else if (3'h0 == state) begin // @[ICache.scala 163:17]
      if (io_cpu_req) begin // @[ICache.scala 165:24]
        if (!(~translation_ok)) begin // @[ICache.scala 166:31]
          arvalid <= _GEN_7204;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 163:17]
      if (3'h2 == state) begin // @[ICache.scala 163:17]
        arvalid <= _GEN_11869;
      end else begin
        arvalid <= _GEN_11913;
      end
    end
    if (reset) begin // @[ICache.scala 147:23]
      rready <= 1'h0; // @[ICache.scala 147:23]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 163:17]
      if (!(3'h1 == state)) begin // @[ICache.scala 163:17]
        if (3'h2 == state) begin // @[ICache.scala 163:17]
          rready <= _GEN_11870;
        end else begin
          rready <= _GEN_11914;
        end
      end
    end
    if (reset) begin // @[ICache.scala 151:21]
      tlb1_invalid <= 1'h0; // @[ICache.scala 151:21]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 163:17]
      if (3'h1 == state) begin // @[ICache.scala 163:17]
        if (!(_T_19)) begin // @[ICache.scala 204:9]
          tlb1_invalid <= 1'h1; // @[ICache.scala 212:24]
        end
      end else if (!(3'h2 == state)) begin // @[ICache.scala 163:17]
        tlb1_invalid <= _GEN_11921;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  meta_0_valid_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  meta_0_valid_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  meta_0_lru = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  meta_1_valid_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  meta_1_valid_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  meta_1_lru = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  meta_2_valid_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  meta_2_valid_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  meta_2_lru = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  meta_3_valid_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  meta_3_valid_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  meta_3_lru = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  meta_4_valid_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  meta_4_valid_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  meta_4_lru = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  meta_5_valid_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  meta_5_valid_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  meta_5_lru = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  meta_6_valid_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  meta_6_valid_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  meta_6_lru = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  meta_7_valid_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  meta_7_valid_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  meta_7_lru = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  meta_8_valid_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  meta_8_valid_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  meta_8_lru = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  meta_9_valid_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  meta_9_valid_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  meta_9_lru = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  meta_10_valid_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  meta_10_valid_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  meta_10_lru = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  meta_11_valid_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  meta_11_valid_1 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  meta_11_lru = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  meta_12_valid_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  meta_12_valid_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  meta_12_lru = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  meta_13_valid_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  meta_13_valid_1 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  meta_13_lru = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  meta_14_valid_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  meta_14_valid_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  meta_14_lru = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  meta_15_valid_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  meta_15_valid_1 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  meta_15_lru = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  meta_16_valid_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  meta_16_valid_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  meta_16_lru = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  meta_17_valid_0 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  meta_17_valid_1 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  meta_17_lru = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  meta_18_valid_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  meta_18_valid_1 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  meta_18_lru = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  meta_19_valid_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  meta_19_valid_1 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  meta_19_lru = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  meta_20_valid_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  meta_20_valid_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  meta_20_lru = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  meta_21_valid_0 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  meta_21_valid_1 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  meta_21_lru = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  meta_22_valid_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  meta_22_valid_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  meta_22_lru = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  meta_23_valid_0 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  meta_23_valid_1 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  meta_23_lru = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  meta_24_valid_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  meta_24_valid_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  meta_24_lru = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  meta_25_valid_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  meta_25_valid_1 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  meta_25_lru = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  meta_26_valid_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  meta_26_valid_1 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  meta_26_lru = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  meta_27_valid_0 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  meta_27_valid_1 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  meta_27_lru = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  meta_28_valid_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  meta_28_valid_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  meta_28_lru = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  meta_29_valid_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  meta_29_valid_1 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  meta_29_lru = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  meta_30_valid_0 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  meta_30_valid_1 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  meta_30_lru = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  meta_31_valid_0 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  meta_31_valid_1 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  meta_31_lru = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  meta_32_valid_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  meta_32_valid_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  meta_32_lru = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  meta_33_valid_0 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  meta_33_valid_1 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  meta_33_lru = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  meta_34_valid_0 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  meta_34_valid_1 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  meta_34_lru = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  meta_35_valid_0 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  meta_35_valid_1 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  meta_35_lru = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  meta_36_valid_0 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  meta_36_valid_1 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  meta_36_lru = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  meta_37_valid_0 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  meta_37_valid_1 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  meta_37_lru = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  meta_38_valid_0 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  meta_38_valid_1 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  meta_38_lru = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  meta_39_valid_0 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  meta_39_valid_1 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  meta_39_lru = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  meta_40_valid_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  meta_40_valid_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  meta_40_lru = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  meta_41_valid_0 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  meta_41_valid_1 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  meta_41_lru = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  meta_42_valid_0 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  meta_42_valid_1 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  meta_42_lru = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  meta_43_valid_0 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  meta_43_valid_1 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  meta_43_lru = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  meta_44_valid_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  meta_44_valid_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  meta_44_lru = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  meta_45_valid_0 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  meta_45_valid_1 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  meta_45_lru = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  meta_46_valid_0 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  meta_46_valid_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  meta_46_lru = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  meta_47_valid_0 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  meta_47_valid_1 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  meta_47_lru = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  meta_48_valid_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  meta_48_valid_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  meta_48_lru = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  meta_49_valid_0 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  meta_49_valid_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  meta_49_lru = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  meta_50_valid_0 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  meta_50_valid_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  meta_50_lru = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  meta_51_valid_0 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  meta_51_valid_1 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  meta_51_lru = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  meta_52_valid_0 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  meta_52_valid_1 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  meta_52_lru = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  meta_53_valid_0 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  meta_53_valid_1 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  meta_53_lru = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  meta_54_valid_0 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  meta_54_valid_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  meta_54_lru = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  meta_55_valid_0 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  meta_55_valid_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  meta_55_lru = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  meta_56_valid_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  meta_56_valid_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  meta_56_lru = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  meta_57_valid_0 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  meta_57_valid_1 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  meta_57_lru = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  meta_58_valid_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  meta_58_valid_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  meta_58_lru = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  meta_59_valid_0 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  meta_59_valid_1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  meta_59_lru = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  meta_60_valid_0 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  meta_60_valid_1 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  meta_60_lru = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  meta_61_valid_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  meta_61_valid_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  meta_61_lru = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  meta_62_valid_0 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  meta_62_valid_1 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  meta_62_lru = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  meta_63_valid_0 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  meta_63_valid_1 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  meta_63_lru = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  meta_64_valid_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  meta_64_valid_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  meta_64_lru = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  meta_65_valid_0 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  meta_65_valid_1 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  meta_65_lru = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  meta_66_valid_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  meta_66_valid_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  meta_66_lru = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  meta_67_valid_0 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  meta_67_valid_1 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  meta_67_lru = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  meta_68_valid_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  meta_68_valid_1 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  meta_68_lru = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  meta_69_valid_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  meta_69_valid_1 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  meta_69_lru = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  meta_70_valid_0 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  meta_70_valid_1 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  meta_70_lru = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  meta_71_valid_0 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  meta_71_valid_1 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  meta_71_lru = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  meta_72_valid_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  meta_72_valid_1 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  meta_72_lru = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  meta_73_valid_0 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  meta_73_valid_1 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  meta_73_lru = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  meta_74_valid_0 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  meta_74_valid_1 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  meta_74_lru = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  meta_75_valid_0 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  meta_75_valid_1 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  meta_75_lru = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  meta_76_valid_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  meta_76_valid_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  meta_76_lru = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  meta_77_valid_0 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  meta_77_valid_1 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  meta_77_lru = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  meta_78_valid_0 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  meta_78_valid_1 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  meta_78_lru = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  meta_79_valid_0 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  meta_79_valid_1 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  meta_79_lru = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  meta_80_valid_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  meta_80_valid_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  meta_80_lru = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  meta_81_valid_0 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  meta_81_valid_1 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  meta_81_lru = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  meta_82_valid_0 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  meta_82_valid_1 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  meta_82_lru = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  meta_83_valid_0 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  meta_83_valid_1 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  meta_83_lru = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  meta_84_valid_0 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  meta_84_valid_1 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  meta_84_lru = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  meta_85_valid_0 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  meta_85_valid_1 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  meta_85_lru = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  meta_86_valid_0 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  meta_86_valid_1 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  meta_86_lru = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  meta_87_valid_0 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  meta_87_valid_1 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  meta_87_lru = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  meta_88_valid_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  meta_88_valid_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  meta_88_lru = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  meta_89_valid_0 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  meta_89_valid_1 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  meta_89_lru = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  meta_90_valid_0 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  meta_90_valid_1 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  meta_90_lru = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  meta_91_valid_0 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  meta_91_valid_1 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  meta_91_lru = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  meta_92_valid_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  meta_92_valid_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  meta_92_lru = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  meta_93_valid_0 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  meta_93_valid_1 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  meta_93_lru = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  meta_94_valid_0 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  meta_94_valid_1 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  meta_94_lru = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  meta_95_valid_0 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  meta_95_valid_1 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  meta_95_lru = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  meta_96_valid_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  meta_96_valid_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  meta_96_lru = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  meta_97_valid_0 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  meta_97_valid_1 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  meta_97_lru = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  meta_98_valid_0 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  meta_98_valid_1 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  meta_98_lru = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  meta_99_valid_0 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  meta_99_valid_1 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  meta_99_lru = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  meta_100_valid_0 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  meta_100_valid_1 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  meta_100_lru = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  meta_101_valid_0 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  meta_101_valid_1 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  meta_101_lru = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  meta_102_valid_0 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  meta_102_valid_1 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  meta_102_lru = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  meta_103_valid_0 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  meta_103_valid_1 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  meta_103_lru = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  meta_104_valid_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  meta_104_valid_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  meta_104_lru = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  meta_105_valid_0 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  meta_105_valid_1 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  meta_105_lru = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  meta_106_valid_0 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  meta_106_valid_1 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  meta_106_lru = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  meta_107_valid_0 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  meta_107_valid_1 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  meta_107_lru = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  meta_108_valid_0 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  meta_108_valid_1 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  meta_108_lru = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  meta_109_valid_0 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  meta_109_valid_1 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  meta_109_lru = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  meta_110_valid_0 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  meta_110_valid_1 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  meta_110_lru = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  meta_111_valid_0 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  meta_111_valid_1 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  meta_111_lru = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  meta_112_valid_0 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  meta_112_valid_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  meta_112_lru = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  meta_113_valid_0 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  meta_113_valid_1 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  meta_113_lru = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  meta_114_valid_0 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  meta_114_valid_1 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  meta_114_lru = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  meta_115_valid_0 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  meta_115_valid_1 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  meta_115_lru = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  meta_116_valid_0 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  meta_116_valid_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  meta_116_lru = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  meta_117_valid_0 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  meta_117_valid_1 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  meta_117_lru = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  meta_118_valid_0 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  meta_118_valid_1 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  meta_118_lru = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  meta_119_valid_0 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  meta_119_valid_1 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  meta_119_lru = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  meta_120_valid_0 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  meta_120_valid_1 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  meta_120_lru = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  meta_121_valid_0 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  meta_121_valid_1 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  meta_121_lru = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  meta_122_valid_0 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  meta_122_valid_1 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  meta_122_lru = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  meta_123_valid_0 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  meta_123_valid_1 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  meta_123_lru = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  meta_124_valid_0 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  meta_124_valid_1 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  meta_124_lru = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  meta_125_valid_0 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  meta_125_valid_1 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  meta_125_lru = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  meta_126_valid_0 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  meta_126_valid_1 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  meta_126_lru = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  meta_127_valid_0 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  meta_127_valid_1 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  meta_127_lru = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  meta_128_valid_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  meta_128_valid_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  meta_128_lru = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  meta_129_valid_0 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  meta_129_valid_1 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  meta_129_lru = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  meta_130_valid_0 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  meta_130_valid_1 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  meta_130_lru = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  meta_131_valid_0 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  meta_131_valid_1 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  meta_131_lru = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  meta_132_valid_0 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  meta_132_valid_1 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  meta_132_lru = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  meta_133_valid_0 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  meta_133_valid_1 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  meta_133_lru = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  meta_134_valid_0 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  meta_134_valid_1 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  meta_134_lru = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  meta_135_valid_0 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  meta_135_valid_1 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  meta_135_lru = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  meta_136_valid_0 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  meta_136_valid_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  meta_136_lru = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  meta_137_valid_0 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  meta_137_valid_1 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  meta_137_lru = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  meta_138_valid_0 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  meta_138_valid_1 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  meta_138_lru = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  meta_139_valid_0 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  meta_139_valid_1 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  meta_139_lru = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  meta_140_valid_0 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  meta_140_valid_1 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  meta_140_lru = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  meta_141_valid_0 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  meta_141_valid_1 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  meta_141_lru = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  meta_142_valid_0 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  meta_142_valid_1 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  meta_142_lru = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  meta_143_valid_0 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  meta_143_valid_1 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  meta_143_lru = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  meta_144_valid_0 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  meta_144_valid_1 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  meta_144_lru = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  meta_145_valid_0 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  meta_145_valid_1 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  meta_145_lru = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  meta_146_valid_0 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  meta_146_valid_1 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  meta_146_lru = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  meta_147_valid_0 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  meta_147_valid_1 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  meta_147_lru = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  meta_148_valid_0 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  meta_148_valid_1 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  meta_148_lru = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  meta_149_valid_0 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  meta_149_valid_1 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  meta_149_lru = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  meta_150_valid_0 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  meta_150_valid_1 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  meta_150_lru = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  meta_151_valid_0 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  meta_151_valid_1 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  meta_151_lru = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  meta_152_valid_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  meta_152_valid_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  meta_152_lru = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  meta_153_valid_0 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  meta_153_valid_1 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  meta_153_lru = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  meta_154_valid_0 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  meta_154_valid_1 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  meta_154_lru = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  meta_155_valid_0 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  meta_155_valid_1 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  meta_155_lru = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  meta_156_valid_0 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  meta_156_valid_1 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  meta_156_lru = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  meta_157_valid_0 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  meta_157_valid_1 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  meta_157_lru = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  meta_158_valid_0 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  meta_158_valid_1 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  meta_158_lru = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  meta_159_valid_0 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  meta_159_valid_1 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  meta_159_lru = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  meta_160_valid_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  meta_160_valid_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  meta_160_lru = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  meta_161_valid_0 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  meta_161_valid_1 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  meta_161_lru = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  meta_162_valid_0 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  meta_162_valid_1 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  meta_162_lru = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  meta_163_valid_0 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  meta_163_valid_1 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  meta_163_lru = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  meta_164_valid_0 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  meta_164_valid_1 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  meta_164_lru = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  meta_165_valid_0 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  meta_165_valid_1 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  meta_165_lru = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  meta_166_valid_0 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  meta_166_valid_1 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  meta_166_lru = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  meta_167_valid_0 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  meta_167_valid_1 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  meta_167_lru = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  meta_168_valid_0 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  meta_168_valid_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  meta_168_lru = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  meta_169_valid_0 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  meta_169_valid_1 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  meta_169_lru = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  meta_170_valid_0 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  meta_170_valid_1 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  meta_170_lru = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  meta_171_valid_0 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  meta_171_valid_1 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  meta_171_lru = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  meta_172_valid_0 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  meta_172_valid_1 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  meta_172_lru = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  meta_173_valid_0 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  meta_173_valid_1 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  meta_173_lru = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  meta_174_valid_0 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  meta_174_valid_1 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  meta_174_lru = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  meta_175_valid_0 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  meta_175_valid_1 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  meta_175_lru = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  meta_176_valid_0 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  meta_176_valid_1 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  meta_176_lru = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  meta_177_valid_0 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  meta_177_valid_1 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  meta_177_lru = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  meta_178_valid_0 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  meta_178_valid_1 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  meta_178_lru = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  meta_179_valid_0 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  meta_179_valid_1 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  meta_179_lru = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  meta_180_valid_0 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  meta_180_valid_1 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  meta_180_lru = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  meta_181_valid_0 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  meta_181_valid_1 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  meta_181_lru = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  meta_182_valid_0 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  meta_182_valid_1 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  meta_182_lru = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  meta_183_valid_0 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  meta_183_valid_1 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  meta_183_lru = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  meta_184_valid_0 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  meta_184_valid_1 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  meta_184_lru = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  meta_185_valid_0 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  meta_185_valid_1 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  meta_185_lru = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  meta_186_valid_0 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  meta_186_valid_1 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  meta_186_lru = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  meta_187_valid_0 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  meta_187_valid_1 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  meta_187_lru = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  meta_188_valid_0 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  meta_188_valid_1 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  meta_188_lru = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  meta_189_valid_0 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  meta_189_valid_1 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  meta_189_lru = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  meta_190_valid_0 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  meta_190_valid_1 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  meta_190_lru = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  meta_191_valid_0 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  meta_191_valid_1 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  meta_191_lru = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  meta_192_valid_0 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  meta_192_valid_1 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  meta_192_lru = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  meta_193_valid_0 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  meta_193_valid_1 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  meta_193_lru = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  meta_194_valid_0 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  meta_194_valid_1 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  meta_194_lru = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  meta_195_valid_0 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  meta_195_valid_1 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  meta_195_lru = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  meta_196_valid_0 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  meta_196_valid_1 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  meta_196_lru = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  meta_197_valid_0 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  meta_197_valid_1 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  meta_197_lru = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  meta_198_valid_0 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  meta_198_valid_1 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  meta_198_lru = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  meta_199_valid_0 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  meta_199_valid_1 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  meta_199_lru = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  meta_200_valid_0 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  meta_200_valid_1 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  meta_200_lru = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  meta_201_valid_0 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  meta_201_valid_1 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  meta_201_lru = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  meta_202_valid_0 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  meta_202_valid_1 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  meta_202_lru = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  meta_203_valid_0 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  meta_203_valid_1 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  meta_203_lru = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  meta_204_valid_0 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  meta_204_valid_1 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  meta_204_lru = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  meta_205_valid_0 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  meta_205_valid_1 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  meta_205_lru = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  meta_206_valid_0 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  meta_206_valid_1 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  meta_206_lru = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  meta_207_valid_0 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  meta_207_valid_1 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  meta_207_lru = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  meta_208_valid_0 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  meta_208_valid_1 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  meta_208_lru = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  meta_209_valid_0 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  meta_209_valid_1 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  meta_209_lru = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  meta_210_valid_0 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  meta_210_valid_1 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  meta_210_lru = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  meta_211_valid_0 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  meta_211_valid_1 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  meta_211_lru = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  meta_212_valid_0 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  meta_212_valid_1 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  meta_212_lru = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  meta_213_valid_0 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  meta_213_valid_1 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  meta_213_lru = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  meta_214_valid_0 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  meta_214_valid_1 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  meta_214_lru = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  meta_215_valid_0 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  meta_215_valid_1 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  meta_215_lru = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  meta_216_valid_0 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  meta_216_valid_1 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  meta_216_lru = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  meta_217_valid_0 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  meta_217_valid_1 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  meta_217_lru = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  meta_218_valid_0 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  meta_218_valid_1 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  meta_218_lru = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  meta_219_valid_0 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  meta_219_valid_1 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  meta_219_lru = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  meta_220_valid_0 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  meta_220_valid_1 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  meta_220_lru = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  meta_221_valid_0 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  meta_221_valid_1 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  meta_221_lru = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  meta_222_valid_0 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  meta_222_valid_1 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  meta_222_lru = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  meta_223_valid_0 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  meta_223_valid_1 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  meta_223_lru = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  meta_224_valid_0 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  meta_224_valid_1 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  meta_224_lru = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  meta_225_valid_0 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  meta_225_valid_1 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  meta_225_lru = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  meta_226_valid_0 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  meta_226_valid_1 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  meta_226_lru = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  meta_227_valid_0 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  meta_227_valid_1 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  meta_227_lru = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  meta_228_valid_0 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  meta_228_valid_1 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  meta_228_lru = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  meta_229_valid_0 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  meta_229_valid_1 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  meta_229_lru = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  meta_230_valid_0 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  meta_230_valid_1 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  meta_230_lru = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  meta_231_valid_0 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  meta_231_valid_1 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  meta_231_lru = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  meta_232_valid_0 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  meta_232_valid_1 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  meta_232_lru = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  meta_233_valid_0 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  meta_233_valid_1 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  meta_233_lru = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  meta_234_valid_0 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  meta_234_valid_1 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  meta_234_lru = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  meta_235_valid_0 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  meta_235_valid_1 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  meta_235_lru = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  meta_236_valid_0 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  meta_236_valid_1 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  meta_236_lru = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  meta_237_valid_0 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  meta_237_valid_1 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  meta_237_lru = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  meta_238_valid_0 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  meta_238_valid_1 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  meta_238_lru = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  meta_239_valid_0 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  meta_239_valid_1 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  meta_239_lru = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  meta_240_valid_0 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  meta_240_valid_1 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  meta_240_lru = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  meta_241_valid_0 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  meta_241_valid_1 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  meta_241_lru = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  meta_242_valid_0 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  meta_242_valid_1 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  meta_242_lru = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  meta_243_valid_0 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  meta_243_valid_1 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  meta_243_lru = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  meta_244_valid_0 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  meta_244_valid_1 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  meta_244_lru = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  meta_245_valid_0 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  meta_245_valid_1 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  meta_245_lru = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  meta_246_valid_0 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  meta_246_valid_1 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  meta_246_lru = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  meta_247_valid_0 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  meta_247_valid_1 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  meta_247_lru = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  meta_248_valid_0 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  meta_248_valid_1 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  meta_248_lru = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  meta_249_valid_0 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  meta_249_valid_1 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  meta_249_lru = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  meta_250_valid_0 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  meta_250_valid_1 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  meta_250_lru = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  meta_251_valid_0 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  meta_251_valid_1 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  meta_251_lru = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  meta_252_valid_0 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  meta_252_valid_1 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  meta_252_lru = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  meta_253_valid_0 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  meta_253_valid_1 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  meta_253_lru = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  meta_254_valid_0 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  meta_254_valid_1 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  meta_254_lru = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  meta_255_valid_0 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  meta_255_valid_1 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  meta_255_lru = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  meta_256_valid_0 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  meta_256_valid_1 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  meta_256_lru = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  meta_257_valid_0 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  meta_257_valid_1 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  meta_257_lru = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  meta_258_valid_0 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  meta_258_valid_1 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  meta_258_lru = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  meta_259_valid_0 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  meta_259_valid_1 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  meta_259_lru = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  meta_260_valid_0 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  meta_260_valid_1 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  meta_260_lru = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  meta_261_valid_0 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  meta_261_valid_1 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  meta_261_lru = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  meta_262_valid_0 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  meta_262_valid_1 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  meta_262_lru = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  meta_263_valid_0 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  meta_263_valid_1 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  meta_263_lru = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  meta_264_valid_0 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  meta_264_valid_1 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  meta_264_lru = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  meta_265_valid_0 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  meta_265_valid_1 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  meta_265_lru = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  meta_266_valid_0 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  meta_266_valid_1 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  meta_266_lru = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  meta_267_valid_0 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  meta_267_valid_1 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  meta_267_lru = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  meta_268_valid_0 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  meta_268_valid_1 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  meta_268_lru = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  meta_269_valid_0 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  meta_269_valid_1 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  meta_269_lru = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  meta_270_valid_0 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  meta_270_valid_1 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  meta_270_lru = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  meta_271_valid_0 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  meta_271_valid_1 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  meta_271_lru = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  meta_272_valid_0 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  meta_272_valid_1 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  meta_272_lru = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  meta_273_valid_0 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  meta_273_valid_1 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  meta_273_lru = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  meta_274_valid_0 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  meta_274_valid_1 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  meta_274_lru = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  meta_275_valid_0 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  meta_275_valid_1 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  meta_275_lru = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  meta_276_valid_0 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  meta_276_valid_1 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  meta_276_lru = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  meta_277_valid_0 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  meta_277_valid_1 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  meta_277_lru = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  meta_278_valid_0 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  meta_278_valid_1 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  meta_278_lru = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  meta_279_valid_0 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  meta_279_valid_1 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  meta_279_lru = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  meta_280_valid_0 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  meta_280_valid_1 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  meta_280_lru = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  meta_281_valid_0 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  meta_281_valid_1 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  meta_281_lru = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  meta_282_valid_0 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  meta_282_valid_1 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  meta_282_lru = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  meta_283_valid_0 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  meta_283_valid_1 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  meta_283_lru = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  meta_284_valid_0 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  meta_284_valid_1 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  meta_284_lru = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  meta_285_valid_0 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  meta_285_valid_1 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  meta_285_lru = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  meta_286_valid_0 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  meta_286_valid_1 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  meta_286_lru = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  meta_287_valid_0 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  meta_287_valid_1 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  meta_287_lru = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  meta_288_valid_0 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  meta_288_valid_1 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  meta_288_lru = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  meta_289_valid_0 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  meta_289_valid_1 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  meta_289_lru = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  meta_290_valid_0 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  meta_290_valid_1 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  meta_290_lru = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  meta_291_valid_0 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  meta_291_valid_1 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  meta_291_lru = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  meta_292_valid_0 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  meta_292_valid_1 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  meta_292_lru = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  meta_293_valid_0 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  meta_293_valid_1 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  meta_293_lru = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  meta_294_valid_0 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  meta_294_valid_1 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  meta_294_lru = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  meta_295_valid_0 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  meta_295_valid_1 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  meta_295_lru = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  meta_296_valid_0 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  meta_296_valid_1 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  meta_296_lru = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  meta_297_valid_0 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  meta_297_valid_1 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  meta_297_lru = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  meta_298_valid_0 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  meta_298_valid_1 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  meta_298_lru = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  meta_299_valid_0 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  meta_299_valid_1 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  meta_299_lru = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  meta_300_valid_0 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  meta_300_valid_1 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  meta_300_lru = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  meta_301_valid_0 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  meta_301_valid_1 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  meta_301_lru = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  meta_302_valid_0 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  meta_302_valid_1 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  meta_302_lru = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  meta_303_valid_0 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  meta_303_valid_1 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  meta_303_lru = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  meta_304_valid_0 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  meta_304_valid_1 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  meta_304_lru = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  meta_305_valid_0 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  meta_305_valid_1 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  meta_305_lru = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  meta_306_valid_0 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  meta_306_valid_1 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  meta_306_lru = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  meta_307_valid_0 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  meta_307_valid_1 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  meta_307_lru = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  meta_308_valid_0 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  meta_308_valid_1 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  meta_308_lru = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  meta_309_valid_0 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  meta_309_valid_1 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  meta_309_lru = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  meta_310_valid_0 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  meta_310_valid_1 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  meta_310_lru = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  meta_311_valid_0 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  meta_311_valid_1 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  meta_311_lru = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  meta_312_valid_0 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  meta_312_valid_1 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  meta_312_lru = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  meta_313_valid_0 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  meta_313_valid_1 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  meta_313_lru = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  meta_314_valid_0 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  meta_314_valid_1 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  meta_314_lru = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  meta_315_valid_0 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  meta_315_valid_1 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  meta_315_lru = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  meta_316_valid_0 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  meta_316_valid_1 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  meta_316_lru = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  meta_317_valid_0 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  meta_317_valid_1 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  meta_317_lru = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  meta_318_valid_0 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  meta_318_valid_1 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  meta_318_lru = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  meta_319_valid_0 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  meta_319_valid_1 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  meta_319_lru = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  meta_320_valid_0 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  meta_320_valid_1 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  meta_320_lru = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  meta_321_valid_0 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  meta_321_valid_1 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  meta_321_lru = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  meta_322_valid_0 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  meta_322_valid_1 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  meta_322_lru = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  meta_323_valid_0 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  meta_323_valid_1 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  meta_323_lru = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  meta_324_valid_0 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  meta_324_valid_1 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  meta_324_lru = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  meta_325_valid_0 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  meta_325_valid_1 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  meta_325_lru = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  meta_326_valid_0 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  meta_326_valid_1 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  meta_326_lru = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  meta_327_valid_0 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  meta_327_valid_1 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  meta_327_lru = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  meta_328_valid_0 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  meta_328_valid_1 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  meta_328_lru = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  meta_329_valid_0 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  meta_329_valid_1 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  meta_329_lru = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  meta_330_valid_0 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  meta_330_valid_1 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  meta_330_lru = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  meta_331_valid_0 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  meta_331_valid_1 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  meta_331_lru = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  meta_332_valid_0 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  meta_332_valid_1 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  meta_332_lru = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  meta_333_valid_0 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  meta_333_valid_1 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  meta_333_lru = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  meta_334_valid_0 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  meta_334_valid_1 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  meta_334_lru = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  meta_335_valid_0 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  meta_335_valid_1 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  meta_335_lru = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  meta_336_valid_0 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  meta_336_valid_1 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  meta_336_lru = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  meta_337_valid_0 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  meta_337_valid_1 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  meta_337_lru = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  meta_338_valid_0 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  meta_338_valid_1 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  meta_338_lru = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  meta_339_valid_0 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  meta_339_valid_1 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  meta_339_lru = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  meta_340_valid_0 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  meta_340_valid_1 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  meta_340_lru = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  meta_341_valid_0 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  meta_341_valid_1 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  meta_341_lru = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  meta_342_valid_0 = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  meta_342_valid_1 = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  meta_342_lru = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  meta_343_valid_0 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  meta_343_valid_1 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  meta_343_lru = _RAND_1031[0:0];
  _RAND_1032 = {1{`RANDOM}};
  meta_344_valid_0 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  meta_344_valid_1 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  meta_344_lru = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  meta_345_valid_0 = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  meta_345_valid_1 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  meta_345_lru = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  meta_346_valid_0 = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  meta_346_valid_1 = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  meta_346_lru = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  meta_347_valid_0 = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  meta_347_valid_1 = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  meta_347_lru = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  meta_348_valid_0 = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  meta_348_valid_1 = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  meta_348_lru = _RAND_1046[0:0];
  _RAND_1047 = {1{`RANDOM}};
  meta_349_valid_0 = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  meta_349_valid_1 = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  meta_349_lru = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  meta_350_valid_0 = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  meta_350_valid_1 = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  meta_350_lru = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  meta_351_valid_0 = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  meta_351_valid_1 = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  meta_351_lru = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  meta_352_valid_0 = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  meta_352_valid_1 = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  meta_352_lru = _RAND_1058[0:0];
  _RAND_1059 = {1{`RANDOM}};
  meta_353_valid_0 = _RAND_1059[0:0];
  _RAND_1060 = {1{`RANDOM}};
  meta_353_valid_1 = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  meta_353_lru = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  meta_354_valid_0 = _RAND_1062[0:0];
  _RAND_1063 = {1{`RANDOM}};
  meta_354_valid_1 = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  meta_354_lru = _RAND_1064[0:0];
  _RAND_1065 = {1{`RANDOM}};
  meta_355_valid_0 = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  meta_355_valid_1 = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  meta_355_lru = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  meta_356_valid_0 = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  meta_356_valid_1 = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  meta_356_lru = _RAND_1070[0:0];
  _RAND_1071 = {1{`RANDOM}};
  meta_357_valid_0 = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  meta_357_valid_1 = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  meta_357_lru = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  meta_358_valid_0 = _RAND_1074[0:0];
  _RAND_1075 = {1{`RANDOM}};
  meta_358_valid_1 = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  meta_358_lru = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  meta_359_valid_0 = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  meta_359_valid_1 = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  meta_359_lru = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  meta_360_valid_0 = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  meta_360_valid_1 = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  meta_360_lru = _RAND_1082[0:0];
  _RAND_1083 = {1{`RANDOM}};
  meta_361_valid_0 = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  meta_361_valid_1 = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  meta_361_lru = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  meta_362_valid_0 = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  meta_362_valid_1 = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  meta_362_lru = _RAND_1088[0:0];
  _RAND_1089 = {1{`RANDOM}};
  meta_363_valid_0 = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  meta_363_valid_1 = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  meta_363_lru = _RAND_1091[0:0];
  _RAND_1092 = {1{`RANDOM}};
  meta_364_valid_0 = _RAND_1092[0:0];
  _RAND_1093 = {1{`RANDOM}};
  meta_364_valid_1 = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  meta_364_lru = _RAND_1094[0:0];
  _RAND_1095 = {1{`RANDOM}};
  meta_365_valid_0 = _RAND_1095[0:0];
  _RAND_1096 = {1{`RANDOM}};
  meta_365_valid_1 = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  meta_365_lru = _RAND_1097[0:0];
  _RAND_1098 = {1{`RANDOM}};
  meta_366_valid_0 = _RAND_1098[0:0];
  _RAND_1099 = {1{`RANDOM}};
  meta_366_valid_1 = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  meta_366_lru = _RAND_1100[0:0];
  _RAND_1101 = {1{`RANDOM}};
  meta_367_valid_0 = _RAND_1101[0:0];
  _RAND_1102 = {1{`RANDOM}};
  meta_367_valid_1 = _RAND_1102[0:0];
  _RAND_1103 = {1{`RANDOM}};
  meta_367_lru = _RAND_1103[0:0];
  _RAND_1104 = {1{`RANDOM}};
  meta_368_valid_0 = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  meta_368_valid_1 = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  meta_368_lru = _RAND_1106[0:0];
  _RAND_1107 = {1{`RANDOM}};
  meta_369_valid_0 = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  meta_369_valid_1 = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  meta_369_lru = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  meta_370_valid_0 = _RAND_1110[0:0];
  _RAND_1111 = {1{`RANDOM}};
  meta_370_valid_1 = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  meta_370_lru = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  meta_371_valid_0 = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  meta_371_valid_1 = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  meta_371_lru = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  meta_372_valid_0 = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  meta_372_valid_1 = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  meta_372_lru = _RAND_1118[0:0];
  _RAND_1119 = {1{`RANDOM}};
  meta_373_valid_0 = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  meta_373_valid_1 = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  meta_373_lru = _RAND_1121[0:0];
  _RAND_1122 = {1{`RANDOM}};
  meta_374_valid_0 = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  meta_374_valid_1 = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  meta_374_lru = _RAND_1124[0:0];
  _RAND_1125 = {1{`RANDOM}};
  meta_375_valid_0 = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  meta_375_valid_1 = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  meta_375_lru = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  meta_376_valid_0 = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  meta_376_valid_1 = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  meta_376_lru = _RAND_1130[0:0];
  _RAND_1131 = {1{`RANDOM}};
  meta_377_valid_0 = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  meta_377_valid_1 = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  meta_377_lru = _RAND_1133[0:0];
  _RAND_1134 = {1{`RANDOM}};
  meta_378_valid_0 = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  meta_378_valid_1 = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  meta_378_lru = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  meta_379_valid_0 = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  meta_379_valid_1 = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  meta_379_lru = _RAND_1139[0:0];
  _RAND_1140 = {1{`RANDOM}};
  meta_380_valid_0 = _RAND_1140[0:0];
  _RAND_1141 = {1{`RANDOM}};
  meta_380_valid_1 = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  meta_380_lru = _RAND_1142[0:0];
  _RAND_1143 = {1{`RANDOM}};
  meta_381_valid_0 = _RAND_1143[0:0];
  _RAND_1144 = {1{`RANDOM}};
  meta_381_valid_1 = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  meta_381_lru = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  meta_382_valid_0 = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  meta_382_valid_1 = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  meta_382_lru = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  meta_383_valid_0 = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  meta_383_valid_1 = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  meta_383_lru = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  meta_384_valid_0 = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  meta_384_valid_1 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  meta_384_lru = _RAND_1154[0:0];
  _RAND_1155 = {1{`RANDOM}};
  meta_385_valid_0 = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  meta_385_valid_1 = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  meta_385_lru = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  meta_386_valid_0 = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  meta_386_valid_1 = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  meta_386_lru = _RAND_1160[0:0];
  _RAND_1161 = {1{`RANDOM}};
  meta_387_valid_0 = _RAND_1161[0:0];
  _RAND_1162 = {1{`RANDOM}};
  meta_387_valid_1 = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  meta_387_lru = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  meta_388_valid_0 = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  meta_388_valid_1 = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  meta_388_lru = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  meta_389_valid_0 = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  meta_389_valid_1 = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  meta_389_lru = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  meta_390_valid_0 = _RAND_1170[0:0];
  _RAND_1171 = {1{`RANDOM}};
  meta_390_valid_1 = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  meta_390_lru = _RAND_1172[0:0];
  _RAND_1173 = {1{`RANDOM}};
  meta_391_valid_0 = _RAND_1173[0:0];
  _RAND_1174 = {1{`RANDOM}};
  meta_391_valid_1 = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  meta_391_lru = _RAND_1175[0:0];
  _RAND_1176 = {1{`RANDOM}};
  meta_392_valid_0 = _RAND_1176[0:0];
  _RAND_1177 = {1{`RANDOM}};
  meta_392_valid_1 = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  meta_392_lru = _RAND_1178[0:0];
  _RAND_1179 = {1{`RANDOM}};
  meta_393_valid_0 = _RAND_1179[0:0];
  _RAND_1180 = {1{`RANDOM}};
  meta_393_valid_1 = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  meta_393_lru = _RAND_1181[0:0];
  _RAND_1182 = {1{`RANDOM}};
  meta_394_valid_0 = _RAND_1182[0:0];
  _RAND_1183 = {1{`RANDOM}};
  meta_394_valid_1 = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  meta_394_lru = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  meta_395_valid_0 = _RAND_1185[0:0];
  _RAND_1186 = {1{`RANDOM}};
  meta_395_valid_1 = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  meta_395_lru = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  meta_396_valid_0 = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  meta_396_valid_1 = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  meta_396_lru = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  meta_397_valid_0 = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  meta_397_valid_1 = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  meta_397_lru = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  meta_398_valid_0 = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  meta_398_valid_1 = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  meta_398_lru = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  meta_399_valid_0 = _RAND_1197[0:0];
  _RAND_1198 = {1{`RANDOM}};
  meta_399_valid_1 = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  meta_399_lru = _RAND_1199[0:0];
  _RAND_1200 = {1{`RANDOM}};
  meta_400_valid_0 = _RAND_1200[0:0];
  _RAND_1201 = {1{`RANDOM}};
  meta_400_valid_1 = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  meta_400_lru = _RAND_1202[0:0];
  _RAND_1203 = {1{`RANDOM}};
  meta_401_valid_0 = _RAND_1203[0:0];
  _RAND_1204 = {1{`RANDOM}};
  meta_401_valid_1 = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  meta_401_lru = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  meta_402_valid_0 = _RAND_1206[0:0];
  _RAND_1207 = {1{`RANDOM}};
  meta_402_valid_1 = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  meta_402_lru = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  meta_403_valid_0 = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  meta_403_valid_1 = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  meta_403_lru = _RAND_1211[0:0];
  _RAND_1212 = {1{`RANDOM}};
  meta_404_valid_0 = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  meta_404_valid_1 = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  meta_404_lru = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  meta_405_valid_0 = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  meta_405_valid_1 = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  meta_405_lru = _RAND_1217[0:0];
  _RAND_1218 = {1{`RANDOM}};
  meta_406_valid_0 = _RAND_1218[0:0];
  _RAND_1219 = {1{`RANDOM}};
  meta_406_valid_1 = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  meta_406_lru = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  meta_407_valid_0 = _RAND_1221[0:0];
  _RAND_1222 = {1{`RANDOM}};
  meta_407_valid_1 = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  meta_407_lru = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  meta_408_valid_0 = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  meta_408_valid_1 = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  meta_408_lru = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  meta_409_valid_0 = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  meta_409_valid_1 = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  meta_409_lru = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  meta_410_valid_0 = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  meta_410_valid_1 = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  meta_410_lru = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  meta_411_valid_0 = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  meta_411_valid_1 = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  meta_411_lru = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  meta_412_valid_0 = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  meta_412_valid_1 = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  meta_412_lru = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  meta_413_valid_0 = _RAND_1239[0:0];
  _RAND_1240 = {1{`RANDOM}};
  meta_413_valid_1 = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  meta_413_lru = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  meta_414_valid_0 = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  meta_414_valid_1 = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  meta_414_lru = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  meta_415_valid_0 = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  meta_415_valid_1 = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  meta_415_lru = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  meta_416_valid_0 = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  meta_416_valid_1 = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  meta_416_lru = _RAND_1250[0:0];
  _RAND_1251 = {1{`RANDOM}};
  meta_417_valid_0 = _RAND_1251[0:0];
  _RAND_1252 = {1{`RANDOM}};
  meta_417_valid_1 = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  meta_417_lru = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  meta_418_valid_0 = _RAND_1254[0:0];
  _RAND_1255 = {1{`RANDOM}};
  meta_418_valid_1 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  meta_418_lru = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  meta_419_valid_0 = _RAND_1257[0:0];
  _RAND_1258 = {1{`RANDOM}};
  meta_419_valid_1 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  meta_419_lru = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  meta_420_valid_0 = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  meta_420_valid_1 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  meta_420_lru = _RAND_1262[0:0];
  _RAND_1263 = {1{`RANDOM}};
  meta_421_valid_0 = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  meta_421_valid_1 = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  meta_421_lru = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  meta_422_valid_0 = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  meta_422_valid_1 = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  meta_422_lru = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  meta_423_valid_0 = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  meta_423_valid_1 = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  meta_423_lru = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  meta_424_valid_0 = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  meta_424_valid_1 = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  meta_424_lru = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  meta_425_valid_0 = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  meta_425_valid_1 = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  meta_425_lru = _RAND_1277[0:0];
  _RAND_1278 = {1{`RANDOM}};
  meta_426_valid_0 = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  meta_426_valid_1 = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  meta_426_lru = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  meta_427_valid_0 = _RAND_1281[0:0];
  _RAND_1282 = {1{`RANDOM}};
  meta_427_valid_1 = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  meta_427_lru = _RAND_1283[0:0];
  _RAND_1284 = {1{`RANDOM}};
  meta_428_valid_0 = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  meta_428_valid_1 = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  meta_428_lru = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  meta_429_valid_0 = _RAND_1287[0:0];
  _RAND_1288 = {1{`RANDOM}};
  meta_429_valid_1 = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  meta_429_lru = _RAND_1289[0:0];
  _RAND_1290 = {1{`RANDOM}};
  meta_430_valid_0 = _RAND_1290[0:0];
  _RAND_1291 = {1{`RANDOM}};
  meta_430_valid_1 = _RAND_1291[0:0];
  _RAND_1292 = {1{`RANDOM}};
  meta_430_lru = _RAND_1292[0:0];
  _RAND_1293 = {1{`RANDOM}};
  meta_431_valid_0 = _RAND_1293[0:0];
  _RAND_1294 = {1{`RANDOM}};
  meta_431_valid_1 = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  meta_431_lru = _RAND_1295[0:0];
  _RAND_1296 = {1{`RANDOM}};
  meta_432_valid_0 = _RAND_1296[0:0];
  _RAND_1297 = {1{`RANDOM}};
  meta_432_valid_1 = _RAND_1297[0:0];
  _RAND_1298 = {1{`RANDOM}};
  meta_432_lru = _RAND_1298[0:0];
  _RAND_1299 = {1{`RANDOM}};
  meta_433_valid_0 = _RAND_1299[0:0];
  _RAND_1300 = {1{`RANDOM}};
  meta_433_valid_1 = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  meta_433_lru = _RAND_1301[0:0];
  _RAND_1302 = {1{`RANDOM}};
  meta_434_valid_0 = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  meta_434_valid_1 = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  meta_434_lru = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  meta_435_valid_0 = _RAND_1305[0:0];
  _RAND_1306 = {1{`RANDOM}};
  meta_435_valid_1 = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  meta_435_lru = _RAND_1307[0:0];
  _RAND_1308 = {1{`RANDOM}};
  meta_436_valid_0 = _RAND_1308[0:0];
  _RAND_1309 = {1{`RANDOM}};
  meta_436_valid_1 = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  meta_436_lru = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  meta_437_valid_0 = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  meta_437_valid_1 = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  meta_437_lru = _RAND_1313[0:0];
  _RAND_1314 = {1{`RANDOM}};
  meta_438_valid_0 = _RAND_1314[0:0];
  _RAND_1315 = {1{`RANDOM}};
  meta_438_valid_1 = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  meta_438_lru = _RAND_1316[0:0];
  _RAND_1317 = {1{`RANDOM}};
  meta_439_valid_0 = _RAND_1317[0:0];
  _RAND_1318 = {1{`RANDOM}};
  meta_439_valid_1 = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  meta_439_lru = _RAND_1319[0:0];
  _RAND_1320 = {1{`RANDOM}};
  meta_440_valid_0 = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  meta_440_valid_1 = _RAND_1321[0:0];
  _RAND_1322 = {1{`RANDOM}};
  meta_440_lru = _RAND_1322[0:0];
  _RAND_1323 = {1{`RANDOM}};
  meta_441_valid_0 = _RAND_1323[0:0];
  _RAND_1324 = {1{`RANDOM}};
  meta_441_valid_1 = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  meta_441_lru = _RAND_1325[0:0];
  _RAND_1326 = {1{`RANDOM}};
  meta_442_valid_0 = _RAND_1326[0:0];
  _RAND_1327 = {1{`RANDOM}};
  meta_442_valid_1 = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  meta_442_lru = _RAND_1328[0:0];
  _RAND_1329 = {1{`RANDOM}};
  meta_443_valid_0 = _RAND_1329[0:0];
  _RAND_1330 = {1{`RANDOM}};
  meta_443_valid_1 = _RAND_1330[0:0];
  _RAND_1331 = {1{`RANDOM}};
  meta_443_lru = _RAND_1331[0:0];
  _RAND_1332 = {1{`RANDOM}};
  meta_444_valid_0 = _RAND_1332[0:0];
  _RAND_1333 = {1{`RANDOM}};
  meta_444_valid_1 = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  meta_444_lru = _RAND_1334[0:0];
  _RAND_1335 = {1{`RANDOM}};
  meta_445_valid_0 = _RAND_1335[0:0];
  _RAND_1336 = {1{`RANDOM}};
  meta_445_valid_1 = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  meta_445_lru = _RAND_1337[0:0];
  _RAND_1338 = {1{`RANDOM}};
  meta_446_valid_0 = _RAND_1338[0:0];
  _RAND_1339 = {1{`RANDOM}};
  meta_446_valid_1 = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  meta_446_lru = _RAND_1340[0:0];
  _RAND_1341 = {1{`RANDOM}};
  meta_447_valid_0 = _RAND_1341[0:0];
  _RAND_1342 = {1{`RANDOM}};
  meta_447_valid_1 = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  meta_447_lru = _RAND_1343[0:0];
  _RAND_1344 = {1{`RANDOM}};
  meta_448_valid_0 = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  meta_448_valid_1 = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  meta_448_lru = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  meta_449_valid_0 = _RAND_1347[0:0];
  _RAND_1348 = {1{`RANDOM}};
  meta_449_valid_1 = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  meta_449_lru = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  meta_450_valid_0 = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  meta_450_valid_1 = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  meta_450_lru = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  meta_451_valid_0 = _RAND_1353[0:0];
  _RAND_1354 = {1{`RANDOM}};
  meta_451_valid_1 = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  meta_451_lru = _RAND_1355[0:0];
  _RAND_1356 = {1{`RANDOM}};
  meta_452_valid_0 = _RAND_1356[0:0];
  _RAND_1357 = {1{`RANDOM}};
  meta_452_valid_1 = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  meta_452_lru = _RAND_1358[0:0];
  _RAND_1359 = {1{`RANDOM}};
  meta_453_valid_0 = _RAND_1359[0:0];
  _RAND_1360 = {1{`RANDOM}};
  meta_453_valid_1 = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  meta_453_lru = _RAND_1361[0:0];
  _RAND_1362 = {1{`RANDOM}};
  meta_454_valid_0 = _RAND_1362[0:0];
  _RAND_1363 = {1{`RANDOM}};
  meta_454_valid_1 = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  meta_454_lru = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  meta_455_valid_0 = _RAND_1365[0:0];
  _RAND_1366 = {1{`RANDOM}};
  meta_455_valid_1 = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  meta_455_lru = _RAND_1367[0:0];
  _RAND_1368 = {1{`RANDOM}};
  meta_456_valid_0 = _RAND_1368[0:0];
  _RAND_1369 = {1{`RANDOM}};
  meta_456_valid_1 = _RAND_1369[0:0];
  _RAND_1370 = {1{`RANDOM}};
  meta_456_lru = _RAND_1370[0:0];
  _RAND_1371 = {1{`RANDOM}};
  meta_457_valid_0 = _RAND_1371[0:0];
  _RAND_1372 = {1{`RANDOM}};
  meta_457_valid_1 = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  meta_457_lru = _RAND_1373[0:0];
  _RAND_1374 = {1{`RANDOM}};
  meta_458_valid_0 = _RAND_1374[0:0];
  _RAND_1375 = {1{`RANDOM}};
  meta_458_valid_1 = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  meta_458_lru = _RAND_1376[0:0];
  _RAND_1377 = {1{`RANDOM}};
  meta_459_valid_0 = _RAND_1377[0:0];
  _RAND_1378 = {1{`RANDOM}};
  meta_459_valid_1 = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  meta_459_lru = _RAND_1379[0:0];
  _RAND_1380 = {1{`RANDOM}};
  meta_460_valid_0 = _RAND_1380[0:0];
  _RAND_1381 = {1{`RANDOM}};
  meta_460_valid_1 = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  meta_460_lru = _RAND_1382[0:0];
  _RAND_1383 = {1{`RANDOM}};
  meta_461_valid_0 = _RAND_1383[0:0];
  _RAND_1384 = {1{`RANDOM}};
  meta_461_valid_1 = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  meta_461_lru = _RAND_1385[0:0];
  _RAND_1386 = {1{`RANDOM}};
  meta_462_valid_0 = _RAND_1386[0:0];
  _RAND_1387 = {1{`RANDOM}};
  meta_462_valid_1 = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  meta_462_lru = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  meta_463_valid_0 = _RAND_1389[0:0];
  _RAND_1390 = {1{`RANDOM}};
  meta_463_valid_1 = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  meta_463_lru = _RAND_1391[0:0];
  _RAND_1392 = {1{`RANDOM}};
  meta_464_valid_0 = _RAND_1392[0:0];
  _RAND_1393 = {1{`RANDOM}};
  meta_464_valid_1 = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  meta_464_lru = _RAND_1394[0:0];
  _RAND_1395 = {1{`RANDOM}};
  meta_465_valid_0 = _RAND_1395[0:0];
  _RAND_1396 = {1{`RANDOM}};
  meta_465_valid_1 = _RAND_1396[0:0];
  _RAND_1397 = {1{`RANDOM}};
  meta_465_lru = _RAND_1397[0:0];
  _RAND_1398 = {1{`RANDOM}};
  meta_466_valid_0 = _RAND_1398[0:0];
  _RAND_1399 = {1{`RANDOM}};
  meta_466_valid_1 = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  meta_466_lru = _RAND_1400[0:0];
  _RAND_1401 = {1{`RANDOM}};
  meta_467_valid_0 = _RAND_1401[0:0];
  _RAND_1402 = {1{`RANDOM}};
  meta_467_valid_1 = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  meta_467_lru = _RAND_1403[0:0];
  _RAND_1404 = {1{`RANDOM}};
  meta_468_valid_0 = _RAND_1404[0:0];
  _RAND_1405 = {1{`RANDOM}};
  meta_468_valid_1 = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  meta_468_lru = _RAND_1406[0:0];
  _RAND_1407 = {1{`RANDOM}};
  meta_469_valid_0 = _RAND_1407[0:0];
  _RAND_1408 = {1{`RANDOM}};
  meta_469_valid_1 = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  meta_469_lru = _RAND_1409[0:0];
  _RAND_1410 = {1{`RANDOM}};
  meta_470_valid_0 = _RAND_1410[0:0];
  _RAND_1411 = {1{`RANDOM}};
  meta_470_valid_1 = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  meta_470_lru = _RAND_1412[0:0];
  _RAND_1413 = {1{`RANDOM}};
  meta_471_valid_0 = _RAND_1413[0:0];
  _RAND_1414 = {1{`RANDOM}};
  meta_471_valid_1 = _RAND_1414[0:0];
  _RAND_1415 = {1{`RANDOM}};
  meta_471_lru = _RAND_1415[0:0];
  _RAND_1416 = {1{`RANDOM}};
  meta_472_valid_0 = _RAND_1416[0:0];
  _RAND_1417 = {1{`RANDOM}};
  meta_472_valid_1 = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  meta_472_lru = _RAND_1418[0:0];
  _RAND_1419 = {1{`RANDOM}};
  meta_473_valid_0 = _RAND_1419[0:0];
  _RAND_1420 = {1{`RANDOM}};
  meta_473_valid_1 = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  meta_473_lru = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  meta_474_valid_0 = _RAND_1422[0:0];
  _RAND_1423 = {1{`RANDOM}};
  meta_474_valid_1 = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  meta_474_lru = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  meta_475_valid_0 = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  meta_475_valid_1 = _RAND_1426[0:0];
  _RAND_1427 = {1{`RANDOM}};
  meta_475_lru = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  meta_476_valid_0 = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  meta_476_valid_1 = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  meta_476_lru = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  meta_477_valid_0 = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  meta_477_valid_1 = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  meta_477_lru = _RAND_1433[0:0];
  _RAND_1434 = {1{`RANDOM}};
  meta_478_valid_0 = _RAND_1434[0:0];
  _RAND_1435 = {1{`RANDOM}};
  meta_478_valid_1 = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  meta_478_lru = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  meta_479_valid_0 = _RAND_1437[0:0];
  _RAND_1438 = {1{`RANDOM}};
  meta_479_valid_1 = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  meta_479_lru = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  meta_480_valid_0 = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  meta_480_valid_1 = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  meta_480_lru = _RAND_1442[0:0];
  _RAND_1443 = {1{`RANDOM}};
  meta_481_valid_0 = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  meta_481_valid_1 = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  meta_481_lru = _RAND_1445[0:0];
  _RAND_1446 = {1{`RANDOM}};
  meta_482_valid_0 = _RAND_1446[0:0];
  _RAND_1447 = {1{`RANDOM}};
  meta_482_valid_1 = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  meta_482_lru = _RAND_1448[0:0];
  _RAND_1449 = {1{`RANDOM}};
  meta_483_valid_0 = _RAND_1449[0:0];
  _RAND_1450 = {1{`RANDOM}};
  meta_483_valid_1 = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  meta_483_lru = _RAND_1451[0:0];
  _RAND_1452 = {1{`RANDOM}};
  meta_484_valid_0 = _RAND_1452[0:0];
  _RAND_1453 = {1{`RANDOM}};
  meta_484_valid_1 = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  meta_484_lru = _RAND_1454[0:0];
  _RAND_1455 = {1{`RANDOM}};
  meta_485_valid_0 = _RAND_1455[0:0];
  _RAND_1456 = {1{`RANDOM}};
  meta_485_valid_1 = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  meta_485_lru = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  meta_486_valid_0 = _RAND_1458[0:0];
  _RAND_1459 = {1{`RANDOM}};
  meta_486_valid_1 = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  meta_486_lru = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  meta_487_valid_0 = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  meta_487_valid_1 = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  meta_487_lru = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  meta_488_valid_0 = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  meta_488_valid_1 = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  meta_488_lru = _RAND_1466[0:0];
  _RAND_1467 = {1{`RANDOM}};
  meta_489_valid_0 = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  meta_489_valid_1 = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  meta_489_lru = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  meta_490_valid_0 = _RAND_1470[0:0];
  _RAND_1471 = {1{`RANDOM}};
  meta_490_valid_1 = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  meta_490_lru = _RAND_1472[0:0];
  _RAND_1473 = {1{`RANDOM}};
  meta_491_valid_0 = _RAND_1473[0:0];
  _RAND_1474 = {1{`RANDOM}};
  meta_491_valid_1 = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  meta_491_lru = _RAND_1475[0:0];
  _RAND_1476 = {1{`RANDOM}};
  meta_492_valid_0 = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  meta_492_valid_1 = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  meta_492_lru = _RAND_1478[0:0];
  _RAND_1479 = {1{`RANDOM}};
  meta_493_valid_0 = _RAND_1479[0:0];
  _RAND_1480 = {1{`RANDOM}};
  meta_493_valid_1 = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  meta_493_lru = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  meta_494_valid_0 = _RAND_1482[0:0];
  _RAND_1483 = {1{`RANDOM}};
  meta_494_valid_1 = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  meta_494_lru = _RAND_1484[0:0];
  _RAND_1485 = {1{`RANDOM}};
  meta_495_valid_0 = _RAND_1485[0:0];
  _RAND_1486 = {1{`RANDOM}};
  meta_495_valid_1 = _RAND_1486[0:0];
  _RAND_1487 = {1{`RANDOM}};
  meta_495_lru = _RAND_1487[0:0];
  _RAND_1488 = {1{`RANDOM}};
  meta_496_valid_0 = _RAND_1488[0:0];
  _RAND_1489 = {1{`RANDOM}};
  meta_496_valid_1 = _RAND_1489[0:0];
  _RAND_1490 = {1{`RANDOM}};
  meta_496_lru = _RAND_1490[0:0];
  _RAND_1491 = {1{`RANDOM}};
  meta_497_valid_0 = _RAND_1491[0:0];
  _RAND_1492 = {1{`RANDOM}};
  meta_497_valid_1 = _RAND_1492[0:0];
  _RAND_1493 = {1{`RANDOM}};
  meta_497_lru = _RAND_1493[0:0];
  _RAND_1494 = {1{`RANDOM}};
  meta_498_valid_0 = _RAND_1494[0:0];
  _RAND_1495 = {1{`RANDOM}};
  meta_498_valid_1 = _RAND_1495[0:0];
  _RAND_1496 = {1{`RANDOM}};
  meta_498_lru = _RAND_1496[0:0];
  _RAND_1497 = {1{`RANDOM}};
  meta_499_valid_0 = _RAND_1497[0:0];
  _RAND_1498 = {1{`RANDOM}};
  meta_499_valid_1 = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  meta_499_lru = _RAND_1499[0:0];
  _RAND_1500 = {1{`RANDOM}};
  meta_500_valid_0 = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  meta_500_valid_1 = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  meta_500_lru = _RAND_1502[0:0];
  _RAND_1503 = {1{`RANDOM}};
  meta_501_valid_0 = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  meta_501_valid_1 = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  meta_501_lru = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  meta_502_valid_0 = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  meta_502_valid_1 = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  meta_502_lru = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  meta_503_valid_0 = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  meta_503_valid_1 = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  meta_503_lru = _RAND_1511[0:0];
  _RAND_1512 = {1{`RANDOM}};
  meta_504_valid_0 = _RAND_1512[0:0];
  _RAND_1513 = {1{`RANDOM}};
  meta_504_valid_1 = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  meta_504_lru = _RAND_1514[0:0];
  _RAND_1515 = {1{`RANDOM}};
  meta_505_valid_0 = _RAND_1515[0:0];
  _RAND_1516 = {1{`RANDOM}};
  meta_505_valid_1 = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  meta_505_lru = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  meta_506_valid_0 = _RAND_1518[0:0];
  _RAND_1519 = {1{`RANDOM}};
  meta_506_valid_1 = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  meta_506_lru = _RAND_1520[0:0];
  _RAND_1521 = {1{`RANDOM}};
  meta_507_valid_0 = _RAND_1521[0:0];
  _RAND_1522 = {1{`RANDOM}};
  meta_507_valid_1 = _RAND_1522[0:0];
  _RAND_1523 = {1{`RANDOM}};
  meta_507_lru = _RAND_1523[0:0];
  _RAND_1524 = {1{`RANDOM}};
  meta_508_valid_0 = _RAND_1524[0:0];
  _RAND_1525 = {1{`RANDOM}};
  meta_508_valid_1 = _RAND_1525[0:0];
  _RAND_1526 = {1{`RANDOM}};
  meta_508_lru = _RAND_1526[0:0];
  _RAND_1527 = {1{`RANDOM}};
  meta_509_valid_0 = _RAND_1527[0:0];
  _RAND_1528 = {1{`RANDOM}};
  meta_509_valid_1 = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  meta_509_lru = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  meta_510_valid_0 = _RAND_1530[0:0];
  _RAND_1531 = {1{`RANDOM}};
  meta_510_valid_1 = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  meta_510_lru = _RAND_1532[0:0];
  _RAND_1533 = {1{`RANDOM}};
  meta_511_valid_0 = _RAND_1533[0:0];
  _RAND_1534 = {1{`RANDOM}};
  meta_511_valid_1 = _RAND_1534[0:0];
  _RAND_1535 = {1{`RANDOM}};
  meta_511_lru = _RAND_1535[0:0];
  _RAND_1536 = {1{`RANDOM}};
  tlb_vpn = _RAND_1536[16:0];
  _RAND_1537 = {1{`RANDOM}};
  tlb_ppn = _RAND_1537[16:0];
  _RAND_1538 = {1{`RANDOM}};
  tlb_uncached = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  tlb_valid = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  state = _RAND_1540[2:0];
  _RAND_1541 = {1{`RANDOM}};
  replace_line_addr = _RAND_1541[5:0];
  _RAND_1542 = {1{`RANDOM}};
  data_wen_0 = _RAND_1542[7:0];
  _RAND_1543 = {1{`RANDOM}};
  data_wen_1 = _RAND_1543[7:0];
  _RAND_1544 = {1{`RANDOM}};
  tag_wen_0 = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  tag_wen_1 = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  tag_ram_wdata = _RAND_1546[16:0];
  _RAND_1547 = {1{`RANDOM}};
  saved_0_inst = _RAND_1547[31:0];
  _RAND_1548 = {1{`RANDOM}};
  saved_0_valid = _RAND_1548[0:0];
  _RAND_1549 = {1{`RANDOM}};
  saved_1_inst = _RAND_1549[31:0];
  _RAND_1550 = {1{`RANDOM}};
  saved_1_valid = _RAND_1550[0:0];
  _RAND_1551 = {1{`RANDOM}};
  axi_cnt = _RAND_1551[4:0];
  _RAND_1552 = {1{`RANDOM}};
  ar_addr = _RAND_1552[31:0];
  _RAND_1553 = {1{`RANDOM}};
  ar_len = _RAND_1553[7:0];
  _RAND_1554 = {1{`RANDOM}};
  ar_size = _RAND_1554[2:0];
  _RAND_1555 = {1{`RANDOM}};
  arvalid = _RAND_1555[0:0];
  _RAND_1556 = {1{`RANDOM}};
  rready = _RAND_1556[0:0];
  _RAND_1557 = {1{`RANDOM}};
  tlb1_invalid = _RAND_1557[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
