module Ctrl(
  input        io_cacheCtrl_iCache_stall,
  input        io_cacheCtrl_dCache_stall,
  output       io_fetchUnit_allow_to_go,
  output       io_instBuffer_delay_slot_do_flush,
  input        io_decoderUnit_inst0_src1_ren,
  input  [4:0] io_decoderUnit_inst0_src1_raddr,
  input        io_decoderUnit_inst0_src2_ren,
  input  [4:0] io_decoderUnit_inst0_src2_raddr,
  input        io_decoderUnit_branch_flag,
  output       io_decoderUnit_allow_to_go,
  output       io_decoderUnit_do_flush,
  input        io_executeUnit_inst_0_mem_ren,
  input  [4:0] io_executeUnit_inst_0_reg_waddr,
  input        io_executeUnit_inst_1_mem_ren,
  input  [4:0] io_executeUnit_inst_1_reg_waddr,
  input        io_executeUnit_fu_stall,
  input        io_executeUnit_branch_flag,
  output       io_executeUnit_allow_to_go,
  output       io_executeUnit_do_flush,
  output       io_executeUnit_fu_allow_to_go,
  output       io_executeUnit_fu_do_flush,
  input        io_memoryUnit_flush_req,
  output       io_memoryUnit_allow_to_go,
  output       io_memoryUnit_do_flush,
  output       io_writeBackUnit_allow_to_go
);
  wire  _inst0_lw_stall_T_5 = io_decoderUnit_inst0_src2_ren & io_decoderUnit_inst0_src2_raddr ==
    io_executeUnit_inst_0_reg_waddr; // @[Ctrl.scala 22:37]
  wire  _inst0_lw_stall_T_6 = io_decoderUnit_inst0_src1_ren & io_decoderUnit_inst0_src1_raddr ==
    io_executeUnit_inst_0_reg_waddr | _inst0_lw_stall_T_5; // @[Ctrl.scala 21:108]
  wire  inst0_lw_stall = io_executeUnit_inst_0_mem_ren & |io_executeUnit_inst_0_reg_waddr & _inst0_lw_stall_T_6; // @[Ctrl.scala 20:99]
  wire  _inst1_lw_stall_T_5 = io_decoderUnit_inst0_src2_ren & io_decoderUnit_inst0_src2_raddr ==
    io_executeUnit_inst_1_reg_waddr; // @[Ctrl.scala 25:37]
  wire  _inst1_lw_stall_T_6 = io_decoderUnit_inst0_src1_ren & io_decoderUnit_inst0_src1_raddr ==
    io_executeUnit_inst_1_reg_waddr | _inst1_lw_stall_T_5; // @[Ctrl.scala 24:108]
  wire  inst1_lw_stall = io_executeUnit_inst_1_mem_ren & |io_executeUnit_inst_1_reg_waddr & _inst1_lw_stall_T_6; // @[Ctrl.scala 23:99]
  wire  lw_stall = inst0_lw_stall | inst1_lw_stall; // @[Ctrl.scala 26:38]
  wire  longest_stall = io_executeUnit_fu_stall | io_cacheCtrl_iCache_stall | io_cacheCtrl_dCache_stall; // @[Ctrl.scala 27:76]
  wire  _io_executeUnit_allow_to_go_T = ~longest_stall; // @[Ctrl.scala 32:36]
  assign io_fetchUnit_allow_to_go = ~io_cacheCtrl_iCache_stall; // @[Ctrl.scala 30:36]
  assign io_instBuffer_delay_slot_do_flush = io_memoryUnit_flush_req; // @[Ctrl.scala 38:37]
  assign io_decoderUnit_allow_to_go = ~(lw_stall | longest_stall); // @[Ctrl.scala 31:36]
  assign io_decoderUnit_do_flush = io_memoryUnit_flush_req | io_executeUnit_branch_flag | io_decoderUnit_branch_flag; // @[Ctrl.scala 39:87]
  assign io_executeUnit_allow_to_go = ~longest_stall; // @[Ctrl.scala 32:36]
  assign io_executeUnit_do_flush = io_memoryUnit_flush_req | io_executeUnit_branch_flag; // @[Ctrl.scala 40:57]
  assign io_executeUnit_fu_allow_to_go = io_memoryUnit_allow_to_go; // @[Ctrl.scala 33:33]
  assign io_executeUnit_fu_do_flush = io_memoryUnit_do_flush; // @[Ctrl.scala 41:30]
  assign io_memoryUnit_allow_to_go = ~longest_stall; // @[Ctrl.scala 34:36]
  assign io_memoryUnit_do_flush = io_memoryUnit_flush_req; // @[Ctrl.scala 42:30]
  assign io_writeBackUnit_allow_to_go = _io_executeUnit_allow_to_go_T | io_memoryUnit_flush_req; // @[Ctrl.scala 35:51]
endmodule
module FetchStage(
  input         clock,
  input         reset,
  input         io_memory_ex,
  input  [31:0] io_memory_ex_pc,
  input         io_memory_flush,
  input  [31:0] io_memory_flush_pc,
  input         io_decoder_branch,
  input  [31:0] io_decoder_target,
  input         io_execute_branch,
  input  [31:0] io_execute_target,
  input         io_instBuffer_full,
  input         io_iCache_inst_valid_0,
  input         io_iCache_inst_valid_1,
  output [31:0] io_iCache_pc,
  output [31:0] io_iCache_pc_next
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[FetchStage.scala 32:19]
  wire [31:0] _io_iCache_pc_next_T_1 = pc + 32'h8; // @[FetchStage.scala 44:38]
  wire [31:0] _io_iCache_pc_next_T_3 = pc + 32'h4; // @[FetchStage.scala 45:38]
  wire [31:0] _io_iCache_pc_next_T_4 = io_iCache_inst_valid_0 ? _io_iCache_pc_next_T_3 : pc; // @[Mux.scala 101:16]
  wire [31:0] _io_iCache_pc_next_T_5 = io_iCache_inst_valid_1 ? _io_iCache_pc_next_T_1 : _io_iCache_pc_next_T_4; // @[Mux.scala 101:16]
  wire [31:0] _io_iCache_pc_next_T_6 = io_instBuffer_full ? pc : _io_iCache_pc_next_T_5; // @[Mux.scala 101:16]
  wire [31:0] _io_iCache_pc_next_T_7 = io_decoder_branch ? io_decoder_target : _io_iCache_pc_next_T_6; // @[Mux.scala 101:16]
  wire [31:0] _io_iCache_pc_next_T_8 = io_execute_branch ? io_execute_target : _io_iCache_pc_next_T_7; // @[Mux.scala 101:16]
  wire [31:0] _io_iCache_pc_next_T_9 = io_memory_flush ? io_memory_flush_pc : _io_iCache_pc_next_T_8; // @[Mux.scala 101:16]
  assign io_iCache_pc = pc; // @[FetchStage.scala 33:16]
  assign io_iCache_pc_next = io_memory_ex ? io_memory_ex_pc : _io_iCache_pc_next_T_9; // @[Mux.scala 101:16]
  always @(posedge clock) begin
    if (reset) begin // @[FetchStage.scala 32:19]
      pc <= 32'hbfc00000; // @[FetchStage.scala 32:19]
    end else begin
      pc <= io_iCache_pc_next; // @[FetchStage.scala 32:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU(
  input         clock,
  input         reset,
  input  [31:0] io_instrD,
  input         io_enaD,
  input  [31:0] io_pcD,
  input  [31:0] io_pc_plus4D,
  input  [31:0] io_pcE,
  input         io_branchE,
  input         io_actual_takeE,
  output        io_branchD,
  output        io_pred_takeD,
  output [31:0] io_branch_targetD
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
`endif // RANDOMIZE_REG_INIT
  wire [13:0] _io_branch_targetD_T_2 = io_instrD[15] ? 14'h3fff : 14'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_branch_targetD_T_4 = {_io_branch_targetD_T_2,io_instrD[15:0],2'h0}; // @[Cat.scala 33:92]
  reg [5:0] BHT_0; // @[BPU.scala 31:26]
  reg [5:0] BHT_1; // @[BPU.scala 31:26]
  reg [5:0] BHT_2; // @[BPU.scala 31:26]
  reg [5:0] BHT_3; // @[BPU.scala 31:26]
  reg [5:0] BHT_4; // @[BPU.scala 31:26]
  reg [5:0] BHT_5; // @[BPU.scala 31:26]
  reg [5:0] BHT_6; // @[BPU.scala 31:26]
  reg [5:0] BHT_7; // @[BPU.scala 31:26]
  reg [5:0] BHT_8; // @[BPU.scala 31:26]
  reg [5:0] BHT_9; // @[BPU.scala 31:26]
  reg [5:0] BHT_10; // @[BPU.scala 31:26]
  reg [5:0] BHT_11; // @[BPU.scala 31:26]
  reg [5:0] BHT_12; // @[BPU.scala 31:26]
  reg [5:0] BHT_13; // @[BPU.scala 31:26]
  reg [5:0] BHT_14; // @[BPU.scala 31:26]
  reg [5:0] BHT_15; // @[BPU.scala 31:26]
  reg [1:0] PHT_0; // @[BPU.scala 32:26]
  reg [1:0] PHT_1; // @[BPU.scala 32:26]
  reg [1:0] PHT_2; // @[BPU.scala 32:26]
  reg [1:0] PHT_3; // @[BPU.scala 32:26]
  reg [1:0] PHT_4; // @[BPU.scala 32:26]
  reg [1:0] PHT_5; // @[BPU.scala 32:26]
  reg [1:0] PHT_6; // @[BPU.scala 32:26]
  reg [1:0] PHT_7; // @[BPU.scala 32:26]
  reg [1:0] PHT_8; // @[BPU.scala 32:26]
  reg [1:0] PHT_9; // @[BPU.scala 32:26]
  reg [1:0] PHT_10; // @[BPU.scala 32:26]
  reg [1:0] PHT_11; // @[BPU.scala 32:26]
  reg [1:0] PHT_12; // @[BPU.scala 32:26]
  reg [1:0] PHT_13; // @[BPU.scala 32:26]
  reg [1:0] PHT_14; // @[BPU.scala 32:26]
  reg [1:0] PHT_15; // @[BPU.scala 32:26]
  reg [1:0] PHT_16; // @[BPU.scala 32:26]
  reg [1:0] PHT_17; // @[BPU.scala 32:26]
  reg [1:0] PHT_18; // @[BPU.scala 32:26]
  reg [1:0] PHT_19; // @[BPU.scala 32:26]
  reg [1:0] PHT_20; // @[BPU.scala 32:26]
  reg [1:0] PHT_21; // @[BPU.scala 32:26]
  reg [1:0] PHT_22; // @[BPU.scala 32:26]
  reg [1:0] PHT_23; // @[BPU.scala 32:26]
  reg [1:0] PHT_24; // @[BPU.scala 32:26]
  reg [1:0] PHT_25; // @[BPU.scala 32:26]
  reg [1:0] PHT_26; // @[BPU.scala 32:26]
  reg [1:0] PHT_27; // @[BPU.scala 32:26]
  reg [1:0] PHT_28; // @[BPU.scala 32:26]
  reg [1:0] PHT_29; // @[BPU.scala 32:26]
  reg [1:0] PHT_30; // @[BPU.scala 32:26]
  reg [1:0] PHT_31; // @[BPU.scala 32:26]
  reg [1:0] PHT_32; // @[BPU.scala 32:26]
  reg [1:0] PHT_33; // @[BPU.scala 32:26]
  reg [1:0] PHT_34; // @[BPU.scala 32:26]
  reg [1:0] PHT_35; // @[BPU.scala 32:26]
  reg [1:0] PHT_36; // @[BPU.scala 32:26]
  reg [1:0] PHT_37; // @[BPU.scala 32:26]
  reg [1:0] PHT_38; // @[BPU.scala 32:26]
  reg [1:0] PHT_39; // @[BPU.scala 32:26]
  reg [1:0] PHT_40; // @[BPU.scala 32:26]
  reg [1:0] PHT_41; // @[BPU.scala 32:26]
  reg [1:0] PHT_42; // @[BPU.scala 32:26]
  reg [1:0] PHT_43; // @[BPU.scala 32:26]
  reg [1:0] PHT_44; // @[BPU.scala 32:26]
  reg [1:0] PHT_45; // @[BPU.scala 32:26]
  reg [1:0] PHT_46; // @[BPU.scala 32:26]
  reg [1:0] PHT_47; // @[BPU.scala 32:26]
  reg [1:0] PHT_48; // @[BPU.scala 32:26]
  reg [1:0] PHT_49; // @[BPU.scala 32:26]
  reg [1:0] PHT_50; // @[BPU.scala 32:26]
  reg [1:0] PHT_51; // @[BPU.scala 32:26]
  reg [1:0] PHT_52; // @[BPU.scala 32:26]
  reg [1:0] PHT_53; // @[BPU.scala 32:26]
  reg [1:0] PHT_54; // @[BPU.scala 32:26]
  reg [1:0] PHT_55; // @[BPU.scala 32:26]
  reg [1:0] PHT_56; // @[BPU.scala 32:26]
  reg [1:0] PHT_57; // @[BPU.scala 32:26]
  reg [1:0] PHT_58; // @[BPU.scala 32:26]
  reg [1:0] PHT_59; // @[BPU.scala 32:26]
  reg [1:0] PHT_60; // @[BPU.scala 32:26]
  reg [1:0] PHT_61; // @[BPU.scala 32:26]
  reg [1:0] PHT_62; // @[BPU.scala 32:26]
  reg [1:0] PHT_63; // @[BPU.scala 32:26]
  wire [3:0] BHT_index = io_pcD[5:2]; // @[BPU.scala 33:25]
  wire [5:0] _GEN_1 = 4'h1 == BHT_index ? BHT_1 : BHT_0; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_2 = 4'h2 == BHT_index ? BHT_2 : _GEN_1; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_3 = 4'h3 == BHT_index ? BHT_3 : _GEN_2; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_4 = 4'h4 == BHT_index ? BHT_4 : _GEN_3; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_5 = 4'h5 == BHT_index ? BHT_5 : _GEN_4; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_6 = 4'h6 == BHT_index ? BHT_6 : _GEN_5; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_7 = 4'h7 == BHT_index ? BHT_7 : _GEN_6; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_8 = 4'h8 == BHT_index ? BHT_8 : _GEN_7; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_9 = 4'h9 == BHT_index ? BHT_9 : _GEN_8; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_10 = 4'ha == BHT_index ? BHT_10 : _GEN_9; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_11 = 4'hb == BHT_index ? BHT_11 : _GEN_10; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_12 = 4'hc == BHT_index ? BHT_12 : _GEN_11; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_13 = 4'hd == BHT_index ? BHT_13 : _GEN_12; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_14 = 4'he == BHT_index ? BHT_14 : _GEN_13; // @[BPU.scala 37:{61,61}]
  wire [5:0] _GEN_15 = 4'hf == BHT_index ? BHT_15 : _GEN_14; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_17 = 6'h1 == _GEN_15 ? PHT_1 : PHT_0; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_18 = 6'h2 == _GEN_15 ? PHT_2 : _GEN_17; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_19 = 6'h3 == _GEN_15 ? PHT_3 : _GEN_18; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_20 = 6'h4 == _GEN_15 ? PHT_4 : _GEN_19; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_21 = 6'h5 == _GEN_15 ? PHT_5 : _GEN_20; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_22 = 6'h6 == _GEN_15 ? PHT_6 : _GEN_21; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_23 = 6'h7 == _GEN_15 ? PHT_7 : _GEN_22; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_24 = 6'h8 == _GEN_15 ? PHT_8 : _GEN_23; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_25 = 6'h9 == _GEN_15 ? PHT_9 : _GEN_24; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_26 = 6'ha == _GEN_15 ? PHT_10 : _GEN_25; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_27 = 6'hb == _GEN_15 ? PHT_11 : _GEN_26; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_28 = 6'hc == _GEN_15 ? PHT_12 : _GEN_27; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_29 = 6'hd == _GEN_15 ? PHT_13 : _GEN_28; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_30 = 6'he == _GEN_15 ? PHT_14 : _GEN_29; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_31 = 6'hf == _GEN_15 ? PHT_15 : _GEN_30; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_32 = 6'h10 == _GEN_15 ? PHT_16 : _GEN_31; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_33 = 6'h11 == _GEN_15 ? PHT_17 : _GEN_32; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_34 = 6'h12 == _GEN_15 ? PHT_18 : _GEN_33; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_35 = 6'h13 == _GEN_15 ? PHT_19 : _GEN_34; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_36 = 6'h14 == _GEN_15 ? PHT_20 : _GEN_35; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_37 = 6'h15 == _GEN_15 ? PHT_21 : _GEN_36; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_38 = 6'h16 == _GEN_15 ? PHT_22 : _GEN_37; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_39 = 6'h17 == _GEN_15 ? PHT_23 : _GEN_38; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_40 = 6'h18 == _GEN_15 ? PHT_24 : _GEN_39; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_41 = 6'h19 == _GEN_15 ? PHT_25 : _GEN_40; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_42 = 6'h1a == _GEN_15 ? PHT_26 : _GEN_41; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_43 = 6'h1b == _GEN_15 ? PHT_27 : _GEN_42; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_44 = 6'h1c == _GEN_15 ? PHT_28 : _GEN_43; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_45 = 6'h1d == _GEN_15 ? PHT_29 : _GEN_44; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_46 = 6'h1e == _GEN_15 ? PHT_30 : _GEN_45; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_47 = 6'h1f == _GEN_15 ? PHT_31 : _GEN_46; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_48 = 6'h20 == _GEN_15 ? PHT_32 : _GEN_47; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_49 = 6'h21 == _GEN_15 ? PHT_33 : _GEN_48; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_50 = 6'h22 == _GEN_15 ? PHT_34 : _GEN_49; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_51 = 6'h23 == _GEN_15 ? PHT_35 : _GEN_50; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_52 = 6'h24 == _GEN_15 ? PHT_36 : _GEN_51; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_53 = 6'h25 == _GEN_15 ? PHT_37 : _GEN_52; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_54 = 6'h26 == _GEN_15 ? PHT_38 : _GEN_53; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_55 = 6'h27 == _GEN_15 ? PHT_39 : _GEN_54; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_56 = 6'h28 == _GEN_15 ? PHT_40 : _GEN_55; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_57 = 6'h29 == _GEN_15 ? PHT_41 : _GEN_56; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_58 = 6'h2a == _GEN_15 ? PHT_42 : _GEN_57; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_59 = 6'h2b == _GEN_15 ? PHT_43 : _GEN_58; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_60 = 6'h2c == _GEN_15 ? PHT_44 : _GEN_59; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_61 = 6'h2d == _GEN_15 ? PHT_45 : _GEN_60; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_62 = 6'h2e == _GEN_15 ? PHT_46 : _GEN_61; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_63 = 6'h2f == _GEN_15 ? PHT_47 : _GEN_62; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_64 = 6'h30 == _GEN_15 ? PHT_48 : _GEN_63; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_65 = 6'h31 == _GEN_15 ? PHT_49 : _GEN_64; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_66 = 6'h32 == _GEN_15 ? PHT_50 : _GEN_65; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_67 = 6'h33 == _GEN_15 ? PHT_51 : _GEN_66; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_68 = 6'h34 == _GEN_15 ? PHT_52 : _GEN_67; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_69 = 6'h35 == _GEN_15 ? PHT_53 : _GEN_68; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_70 = 6'h36 == _GEN_15 ? PHT_54 : _GEN_69; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_71 = 6'h37 == _GEN_15 ? PHT_55 : _GEN_70; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_72 = 6'h38 == _GEN_15 ? PHT_56 : _GEN_71; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_73 = 6'h39 == _GEN_15 ? PHT_57 : _GEN_72; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_74 = 6'h3a == _GEN_15 ? PHT_58 : _GEN_73; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_75 = 6'h3b == _GEN_15 ? PHT_59 : _GEN_74; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_76 = 6'h3c == _GEN_15 ? PHT_60 : _GEN_75; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_77 = 6'h3d == _GEN_15 ? PHT_61 : _GEN_76; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_78 = 6'h3e == _GEN_15 ? PHT_62 : _GEN_77; // @[BPU.scala 37:{61,61}]
  wire [1:0] _GEN_79 = 6'h3f == _GEN_15 ? PHT_63 : _GEN_78; // @[BPU.scala 37:{61,61}]
  wire [3:0] update_BHT_index = io_pcE[5:2]; // @[BPU.scala 39:32]
  wire [5:0] _GEN_145 = 4'h1 == update_BHT_index ? BHT_1 : BHT_0; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_146 = 4'h2 == update_BHT_index ? BHT_2 : _GEN_145; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_147 = 4'h3 == update_BHT_index ? BHT_3 : _GEN_146; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_148 = 4'h4 == update_BHT_index ? BHT_4 : _GEN_147; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_149 = 4'h5 == update_BHT_index ? BHT_5 : _GEN_148; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_150 = 4'h6 == update_BHT_index ? BHT_6 : _GEN_149; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_151 = 4'h7 == update_BHT_index ? BHT_7 : _GEN_150; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_152 = 4'h8 == update_BHT_index ? BHT_8 : _GEN_151; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_153 = 4'h9 == update_BHT_index ? BHT_9 : _GEN_152; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_154 = 4'ha == update_BHT_index ? BHT_10 : _GEN_153; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_155 = 4'hb == update_BHT_index ? BHT_11 : _GEN_154; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_156 = 4'hc == update_BHT_index ? BHT_12 : _GEN_155; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_157 = 4'hd == update_BHT_index ? BHT_13 : _GEN_156; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_158 = 4'he == update_BHT_index ? BHT_14 : _GEN_157; // @[BPU.scala 44:{55,55}]
  wire [5:0] _GEN_159 = 4'hf == update_BHT_index ? BHT_15 : _GEN_158; // @[BPU.scala 44:{55,55}]
  wire [5:0] _BHT_T_1 = {_GEN_159[5:1],io_actual_takeE}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_177 = 6'h1 == _GEN_159 ? PHT_1 : PHT_0; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_178 = 6'h2 == _GEN_159 ? PHT_2 : _GEN_177; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_179 = 6'h3 == _GEN_159 ? PHT_3 : _GEN_178; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_180 = 6'h4 == _GEN_159 ? PHT_4 : _GEN_179; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_181 = 6'h5 == _GEN_159 ? PHT_5 : _GEN_180; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_182 = 6'h6 == _GEN_159 ? PHT_6 : _GEN_181; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_183 = 6'h7 == _GEN_159 ? PHT_7 : _GEN_182; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_184 = 6'h8 == _GEN_159 ? PHT_8 : _GEN_183; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_185 = 6'h9 == _GEN_159 ? PHT_9 : _GEN_184; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_186 = 6'ha == _GEN_159 ? PHT_10 : _GEN_185; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_187 = 6'hb == _GEN_159 ? PHT_11 : _GEN_186; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_188 = 6'hc == _GEN_159 ? PHT_12 : _GEN_187; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_189 = 6'hd == _GEN_159 ? PHT_13 : _GEN_188; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_190 = 6'he == _GEN_159 ? PHT_14 : _GEN_189; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_191 = 6'hf == _GEN_159 ? PHT_15 : _GEN_190; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_192 = 6'h10 == _GEN_159 ? PHT_16 : _GEN_191; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_193 = 6'h11 == _GEN_159 ? PHT_17 : _GEN_192; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_194 = 6'h12 == _GEN_159 ? PHT_18 : _GEN_193; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_195 = 6'h13 == _GEN_159 ? PHT_19 : _GEN_194; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_196 = 6'h14 == _GEN_159 ? PHT_20 : _GEN_195; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_197 = 6'h15 == _GEN_159 ? PHT_21 : _GEN_196; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_198 = 6'h16 == _GEN_159 ? PHT_22 : _GEN_197; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_199 = 6'h17 == _GEN_159 ? PHT_23 : _GEN_198; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_200 = 6'h18 == _GEN_159 ? PHT_24 : _GEN_199; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_201 = 6'h19 == _GEN_159 ? PHT_25 : _GEN_200; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_202 = 6'h1a == _GEN_159 ? PHT_26 : _GEN_201; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_203 = 6'h1b == _GEN_159 ? PHT_27 : _GEN_202; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_204 = 6'h1c == _GEN_159 ? PHT_28 : _GEN_203; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_205 = 6'h1d == _GEN_159 ? PHT_29 : _GEN_204; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_206 = 6'h1e == _GEN_159 ? PHT_30 : _GEN_205; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_207 = 6'h1f == _GEN_159 ? PHT_31 : _GEN_206; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_208 = 6'h20 == _GEN_159 ? PHT_32 : _GEN_207; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_209 = 6'h21 == _GEN_159 ? PHT_33 : _GEN_208; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_210 = 6'h22 == _GEN_159 ? PHT_34 : _GEN_209; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_211 = 6'h23 == _GEN_159 ? PHT_35 : _GEN_210; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_212 = 6'h24 == _GEN_159 ? PHT_36 : _GEN_211; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_213 = 6'h25 == _GEN_159 ? PHT_37 : _GEN_212; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_214 = 6'h26 == _GEN_159 ? PHT_38 : _GEN_213; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_215 = 6'h27 == _GEN_159 ? PHT_39 : _GEN_214; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_216 = 6'h28 == _GEN_159 ? PHT_40 : _GEN_215; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_217 = 6'h29 == _GEN_159 ? PHT_41 : _GEN_216; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_218 = 6'h2a == _GEN_159 ? PHT_42 : _GEN_217; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_219 = 6'h2b == _GEN_159 ? PHT_43 : _GEN_218; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_220 = 6'h2c == _GEN_159 ? PHT_44 : _GEN_219; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_221 = 6'h2d == _GEN_159 ? PHT_45 : _GEN_220; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_222 = 6'h2e == _GEN_159 ? PHT_46 : _GEN_221; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_223 = 6'h2f == _GEN_159 ? PHT_47 : _GEN_222; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_224 = 6'h30 == _GEN_159 ? PHT_48 : _GEN_223; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_225 = 6'h31 == _GEN_159 ? PHT_49 : _GEN_224; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_226 = 6'h32 == _GEN_159 ? PHT_50 : _GEN_225; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_227 = 6'h33 == _GEN_159 ? PHT_51 : _GEN_226; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_228 = 6'h34 == _GEN_159 ? PHT_52 : _GEN_227; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_229 = 6'h35 == _GEN_159 ? PHT_53 : _GEN_228; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_230 = 6'h36 == _GEN_159 ? PHT_54 : _GEN_229; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_231 = 6'h37 == _GEN_159 ? PHT_55 : _GEN_230; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_232 = 6'h38 == _GEN_159 ? PHT_56 : _GEN_231; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_233 = 6'h39 == _GEN_159 ? PHT_57 : _GEN_232; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_234 = 6'h3a == _GEN_159 ? PHT_58 : _GEN_233; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_235 = 6'h3b == _GEN_159 ? PHT_59 : _GEN_234; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_236 = 6'h3c == _GEN_159 ? PHT_60 : _GEN_235; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_237 = 6'h3d == _GEN_159 ? PHT_61 : _GEN_236; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_238 = 6'h3e == _GEN_159 ? PHT_62 : _GEN_237; // @[BPU.scala 45:{35,35}]
  wire [1:0] _GEN_239 = 6'h3f == _GEN_159 ? PHT_63 : _GEN_238; // @[BPU.scala 45:{35,35}]
  wire [1:0] _PHT_T = io_actual_takeE ? 2'h1 : 2'h0; // @[BPU.scala 47:37]
  wire [1:0] _PHT_T_1 = io_actual_takeE ? 2'h2 : 2'h0; // @[BPU.scala 50:37]
  wire [1:0] _GEN_368 = 6'h0 == _GEN_159 ? _PHT_T_1 : PHT_0; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_369 = 6'h1 == _GEN_159 ? _PHT_T_1 : PHT_1; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_370 = 6'h2 == _GEN_159 ? _PHT_T_1 : PHT_2; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_371 = 6'h3 == _GEN_159 ? _PHT_T_1 : PHT_3; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_372 = 6'h4 == _GEN_159 ? _PHT_T_1 : PHT_4; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_373 = 6'h5 == _GEN_159 ? _PHT_T_1 : PHT_5; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_374 = 6'h6 == _GEN_159 ? _PHT_T_1 : PHT_6; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_375 = 6'h7 == _GEN_159 ? _PHT_T_1 : PHT_7; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_376 = 6'h8 == _GEN_159 ? _PHT_T_1 : PHT_8; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_377 = 6'h9 == _GEN_159 ? _PHT_T_1 : PHT_9; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_378 = 6'ha == _GEN_159 ? _PHT_T_1 : PHT_10; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_379 = 6'hb == _GEN_159 ? _PHT_T_1 : PHT_11; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_380 = 6'hc == _GEN_159 ? _PHT_T_1 : PHT_12; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_381 = 6'hd == _GEN_159 ? _PHT_T_1 : PHT_13; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_382 = 6'he == _GEN_159 ? _PHT_T_1 : PHT_14; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_383 = 6'hf == _GEN_159 ? _PHT_T_1 : PHT_15; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_384 = 6'h10 == _GEN_159 ? _PHT_T_1 : PHT_16; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_385 = 6'h11 == _GEN_159 ? _PHT_T_1 : PHT_17; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_386 = 6'h12 == _GEN_159 ? _PHT_T_1 : PHT_18; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_387 = 6'h13 == _GEN_159 ? _PHT_T_1 : PHT_19; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_388 = 6'h14 == _GEN_159 ? _PHT_T_1 : PHT_20; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_389 = 6'h15 == _GEN_159 ? _PHT_T_1 : PHT_21; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_390 = 6'h16 == _GEN_159 ? _PHT_T_1 : PHT_22; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_391 = 6'h17 == _GEN_159 ? _PHT_T_1 : PHT_23; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_392 = 6'h18 == _GEN_159 ? _PHT_T_1 : PHT_24; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_393 = 6'h19 == _GEN_159 ? _PHT_T_1 : PHT_25; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_394 = 6'h1a == _GEN_159 ? _PHT_T_1 : PHT_26; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_395 = 6'h1b == _GEN_159 ? _PHT_T_1 : PHT_27; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_396 = 6'h1c == _GEN_159 ? _PHT_T_1 : PHT_28; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_397 = 6'h1d == _GEN_159 ? _PHT_T_1 : PHT_29; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_398 = 6'h1e == _GEN_159 ? _PHT_T_1 : PHT_30; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_399 = 6'h1f == _GEN_159 ? _PHT_T_1 : PHT_31; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_400 = 6'h20 == _GEN_159 ? _PHT_T_1 : PHT_32; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_401 = 6'h21 == _GEN_159 ? _PHT_T_1 : PHT_33; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_402 = 6'h22 == _GEN_159 ? _PHT_T_1 : PHT_34; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_403 = 6'h23 == _GEN_159 ? _PHT_T_1 : PHT_35; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_404 = 6'h24 == _GEN_159 ? _PHT_T_1 : PHT_36; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_405 = 6'h25 == _GEN_159 ? _PHT_T_1 : PHT_37; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_406 = 6'h26 == _GEN_159 ? _PHT_T_1 : PHT_38; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_407 = 6'h27 == _GEN_159 ? _PHT_T_1 : PHT_39; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_408 = 6'h28 == _GEN_159 ? _PHT_T_1 : PHT_40; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_409 = 6'h29 == _GEN_159 ? _PHT_T_1 : PHT_41; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_410 = 6'h2a == _GEN_159 ? _PHT_T_1 : PHT_42; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_411 = 6'h2b == _GEN_159 ? _PHT_T_1 : PHT_43; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_412 = 6'h2c == _GEN_159 ? _PHT_T_1 : PHT_44; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_413 = 6'h2d == _GEN_159 ? _PHT_T_1 : PHT_45; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_414 = 6'h2e == _GEN_159 ? _PHT_T_1 : PHT_46; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_415 = 6'h2f == _GEN_159 ? _PHT_T_1 : PHT_47; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_416 = 6'h30 == _GEN_159 ? _PHT_T_1 : PHT_48; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_417 = 6'h31 == _GEN_159 ? _PHT_T_1 : PHT_49; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_418 = 6'h32 == _GEN_159 ? _PHT_T_1 : PHT_50; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_419 = 6'h33 == _GEN_159 ? _PHT_T_1 : PHT_51; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_420 = 6'h34 == _GEN_159 ? _PHT_T_1 : PHT_52; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_421 = 6'h35 == _GEN_159 ? _PHT_T_1 : PHT_53; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_422 = 6'h36 == _GEN_159 ? _PHT_T_1 : PHT_54; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_423 = 6'h37 == _GEN_159 ? _PHT_T_1 : PHT_55; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_424 = 6'h38 == _GEN_159 ? _PHT_T_1 : PHT_56; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_425 = 6'h39 == _GEN_159 ? _PHT_T_1 : PHT_57; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_426 = 6'h3a == _GEN_159 ? _PHT_T_1 : PHT_58; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_427 = 6'h3b == _GEN_159 ? _PHT_T_1 : PHT_59; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_428 = 6'h3c == _GEN_159 ? _PHT_T_1 : PHT_60; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_429 = 6'h3d == _GEN_159 ? _PHT_T_1 : PHT_61; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_430 = 6'h3e == _GEN_159 ? _PHT_T_1 : PHT_62; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _GEN_431 = 6'h3f == _GEN_159 ? _PHT_T_1 : PHT_63; // @[BPU.scala 32:26 50:{31,31}]
  wire [1:0] _PHT_T_2 = io_actual_takeE ? 2'h3 : 2'h1; // @[BPU.scala 53:37]
  wire [1:0] _GEN_496 = 6'h0 == _GEN_159 ? _PHT_T_2 : PHT_0; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_497 = 6'h1 == _GEN_159 ? _PHT_T_2 : PHT_1; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_498 = 6'h2 == _GEN_159 ? _PHT_T_2 : PHT_2; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_499 = 6'h3 == _GEN_159 ? _PHT_T_2 : PHT_3; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_500 = 6'h4 == _GEN_159 ? _PHT_T_2 : PHT_4; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_501 = 6'h5 == _GEN_159 ? _PHT_T_2 : PHT_5; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_502 = 6'h6 == _GEN_159 ? _PHT_T_2 : PHT_6; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_503 = 6'h7 == _GEN_159 ? _PHT_T_2 : PHT_7; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_504 = 6'h8 == _GEN_159 ? _PHT_T_2 : PHT_8; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_505 = 6'h9 == _GEN_159 ? _PHT_T_2 : PHT_9; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_506 = 6'ha == _GEN_159 ? _PHT_T_2 : PHT_10; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_507 = 6'hb == _GEN_159 ? _PHT_T_2 : PHT_11; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_508 = 6'hc == _GEN_159 ? _PHT_T_2 : PHT_12; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_509 = 6'hd == _GEN_159 ? _PHT_T_2 : PHT_13; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_510 = 6'he == _GEN_159 ? _PHT_T_2 : PHT_14; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_511 = 6'hf == _GEN_159 ? _PHT_T_2 : PHT_15; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_512 = 6'h10 == _GEN_159 ? _PHT_T_2 : PHT_16; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_513 = 6'h11 == _GEN_159 ? _PHT_T_2 : PHT_17; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_514 = 6'h12 == _GEN_159 ? _PHT_T_2 : PHT_18; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_515 = 6'h13 == _GEN_159 ? _PHT_T_2 : PHT_19; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_516 = 6'h14 == _GEN_159 ? _PHT_T_2 : PHT_20; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_517 = 6'h15 == _GEN_159 ? _PHT_T_2 : PHT_21; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_518 = 6'h16 == _GEN_159 ? _PHT_T_2 : PHT_22; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_519 = 6'h17 == _GEN_159 ? _PHT_T_2 : PHT_23; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_520 = 6'h18 == _GEN_159 ? _PHT_T_2 : PHT_24; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_521 = 6'h19 == _GEN_159 ? _PHT_T_2 : PHT_25; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_522 = 6'h1a == _GEN_159 ? _PHT_T_2 : PHT_26; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_523 = 6'h1b == _GEN_159 ? _PHT_T_2 : PHT_27; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_524 = 6'h1c == _GEN_159 ? _PHT_T_2 : PHT_28; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_525 = 6'h1d == _GEN_159 ? _PHT_T_2 : PHT_29; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_526 = 6'h1e == _GEN_159 ? _PHT_T_2 : PHT_30; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_527 = 6'h1f == _GEN_159 ? _PHT_T_2 : PHT_31; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_528 = 6'h20 == _GEN_159 ? _PHT_T_2 : PHT_32; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_529 = 6'h21 == _GEN_159 ? _PHT_T_2 : PHT_33; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_530 = 6'h22 == _GEN_159 ? _PHT_T_2 : PHT_34; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_531 = 6'h23 == _GEN_159 ? _PHT_T_2 : PHT_35; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_532 = 6'h24 == _GEN_159 ? _PHT_T_2 : PHT_36; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_533 = 6'h25 == _GEN_159 ? _PHT_T_2 : PHT_37; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_534 = 6'h26 == _GEN_159 ? _PHT_T_2 : PHT_38; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_535 = 6'h27 == _GEN_159 ? _PHT_T_2 : PHT_39; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_536 = 6'h28 == _GEN_159 ? _PHT_T_2 : PHT_40; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_537 = 6'h29 == _GEN_159 ? _PHT_T_2 : PHT_41; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_538 = 6'h2a == _GEN_159 ? _PHT_T_2 : PHT_42; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_539 = 6'h2b == _GEN_159 ? _PHT_T_2 : PHT_43; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_540 = 6'h2c == _GEN_159 ? _PHT_T_2 : PHT_44; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_541 = 6'h2d == _GEN_159 ? _PHT_T_2 : PHT_45; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_542 = 6'h2e == _GEN_159 ? _PHT_T_2 : PHT_46; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_543 = 6'h2f == _GEN_159 ? _PHT_T_2 : PHT_47; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_544 = 6'h30 == _GEN_159 ? _PHT_T_2 : PHT_48; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_545 = 6'h31 == _GEN_159 ? _PHT_T_2 : PHT_49; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_546 = 6'h32 == _GEN_159 ? _PHT_T_2 : PHT_50; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_547 = 6'h33 == _GEN_159 ? _PHT_T_2 : PHT_51; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_548 = 6'h34 == _GEN_159 ? _PHT_T_2 : PHT_52; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_549 = 6'h35 == _GEN_159 ? _PHT_T_2 : PHT_53; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_550 = 6'h36 == _GEN_159 ? _PHT_T_2 : PHT_54; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_551 = 6'h37 == _GEN_159 ? _PHT_T_2 : PHT_55; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_552 = 6'h38 == _GEN_159 ? _PHT_T_2 : PHT_56; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_553 = 6'h39 == _GEN_159 ? _PHT_T_2 : PHT_57; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_554 = 6'h3a == _GEN_159 ? _PHT_T_2 : PHT_58; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_555 = 6'h3b == _GEN_159 ? _PHT_T_2 : PHT_59; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_556 = 6'h3c == _GEN_159 ? _PHT_T_2 : PHT_60; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_557 = 6'h3d == _GEN_159 ? _PHT_T_2 : PHT_61; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_558 = 6'h3e == _GEN_159 ? _PHT_T_2 : PHT_62; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _GEN_559 = 6'h3f == _GEN_159 ? _PHT_T_2 : PHT_63; // @[BPU.scala 32:26 53:{31,31}]
  wire [1:0] _PHT_T_3 = io_actual_takeE ? 2'h3 : 2'h2; // @[BPU.scala 56:37]
  wire [1:0] _GEN_624 = 6'h0 == _GEN_159 ? _PHT_T_3 : PHT_0; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_625 = 6'h1 == _GEN_159 ? _PHT_T_3 : PHT_1; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_626 = 6'h2 == _GEN_159 ? _PHT_T_3 : PHT_2; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_627 = 6'h3 == _GEN_159 ? _PHT_T_3 : PHT_3; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_628 = 6'h4 == _GEN_159 ? _PHT_T_3 : PHT_4; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_629 = 6'h5 == _GEN_159 ? _PHT_T_3 : PHT_5; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_630 = 6'h6 == _GEN_159 ? _PHT_T_3 : PHT_6; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_631 = 6'h7 == _GEN_159 ? _PHT_T_3 : PHT_7; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_632 = 6'h8 == _GEN_159 ? _PHT_T_3 : PHT_8; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_633 = 6'h9 == _GEN_159 ? _PHT_T_3 : PHT_9; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_634 = 6'ha == _GEN_159 ? _PHT_T_3 : PHT_10; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_635 = 6'hb == _GEN_159 ? _PHT_T_3 : PHT_11; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_636 = 6'hc == _GEN_159 ? _PHT_T_3 : PHT_12; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_637 = 6'hd == _GEN_159 ? _PHT_T_3 : PHT_13; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_638 = 6'he == _GEN_159 ? _PHT_T_3 : PHT_14; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_639 = 6'hf == _GEN_159 ? _PHT_T_3 : PHT_15; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_640 = 6'h10 == _GEN_159 ? _PHT_T_3 : PHT_16; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_641 = 6'h11 == _GEN_159 ? _PHT_T_3 : PHT_17; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_642 = 6'h12 == _GEN_159 ? _PHT_T_3 : PHT_18; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_643 = 6'h13 == _GEN_159 ? _PHT_T_3 : PHT_19; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_644 = 6'h14 == _GEN_159 ? _PHT_T_3 : PHT_20; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_645 = 6'h15 == _GEN_159 ? _PHT_T_3 : PHT_21; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_646 = 6'h16 == _GEN_159 ? _PHT_T_3 : PHT_22; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_647 = 6'h17 == _GEN_159 ? _PHT_T_3 : PHT_23; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_648 = 6'h18 == _GEN_159 ? _PHT_T_3 : PHT_24; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_649 = 6'h19 == _GEN_159 ? _PHT_T_3 : PHT_25; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_650 = 6'h1a == _GEN_159 ? _PHT_T_3 : PHT_26; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_651 = 6'h1b == _GEN_159 ? _PHT_T_3 : PHT_27; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_652 = 6'h1c == _GEN_159 ? _PHT_T_3 : PHT_28; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_653 = 6'h1d == _GEN_159 ? _PHT_T_3 : PHT_29; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_654 = 6'h1e == _GEN_159 ? _PHT_T_3 : PHT_30; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_655 = 6'h1f == _GEN_159 ? _PHT_T_3 : PHT_31; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_656 = 6'h20 == _GEN_159 ? _PHT_T_3 : PHT_32; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_657 = 6'h21 == _GEN_159 ? _PHT_T_3 : PHT_33; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_658 = 6'h22 == _GEN_159 ? _PHT_T_3 : PHT_34; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_659 = 6'h23 == _GEN_159 ? _PHT_T_3 : PHT_35; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_660 = 6'h24 == _GEN_159 ? _PHT_T_3 : PHT_36; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_661 = 6'h25 == _GEN_159 ? _PHT_T_3 : PHT_37; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_662 = 6'h26 == _GEN_159 ? _PHT_T_3 : PHT_38; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_663 = 6'h27 == _GEN_159 ? _PHT_T_3 : PHT_39; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_664 = 6'h28 == _GEN_159 ? _PHT_T_3 : PHT_40; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_665 = 6'h29 == _GEN_159 ? _PHT_T_3 : PHT_41; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_666 = 6'h2a == _GEN_159 ? _PHT_T_3 : PHT_42; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_667 = 6'h2b == _GEN_159 ? _PHT_T_3 : PHT_43; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_668 = 6'h2c == _GEN_159 ? _PHT_T_3 : PHT_44; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_669 = 6'h2d == _GEN_159 ? _PHT_T_3 : PHT_45; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_670 = 6'h2e == _GEN_159 ? _PHT_T_3 : PHT_46; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_671 = 6'h2f == _GEN_159 ? _PHT_T_3 : PHT_47; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_672 = 6'h30 == _GEN_159 ? _PHT_T_3 : PHT_48; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_673 = 6'h31 == _GEN_159 ? _PHT_T_3 : PHT_49; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_674 = 6'h32 == _GEN_159 ? _PHT_T_3 : PHT_50; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_675 = 6'h33 == _GEN_159 ? _PHT_T_3 : PHT_51; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_676 = 6'h34 == _GEN_159 ? _PHT_T_3 : PHT_52; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_677 = 6'h35 == _GEN_159 ? _PHT_T_3 : PHT_53; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_678 = 6'h36 == _GEN_159 ? _PHT_T_3 : PHT_54; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_679 = 6'h37 == _GEN_159 ? _PHT_T_3 : PHT_55; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_680 = 6'h38 == _GEN_159 ? _PHT_T_3 : PHT_56; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_681 = 6'h39 == _GEN_159 ? _PHT_T_3 : PHT_57; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_682 = 6'h3a == _GEN_159 ? _PHT_T_3 : PHT_58; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_683 = 6'h3b == _GEN_159 ? _PHT_T_3 : PHT_59; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_684 = 6'h3c == _GEN_159 ? _PHT_T_3 : PHT_60; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_685 = 6'h3d == _GEN_159 ? _PHT_T_3 : PHT_61; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_686 = 6'h3e == _GEN_159 ? _PHT_T_3 : PHT_62; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_687 = 6'h3f == _GEN_159 ? _PHT_T_3 : PHT_63; // @[BPU.scala 32:26 56:{31,31}]
  wire [1:0] _GEN_688 = 2'h3 == _GEN_239 ? _GEN_624 : PHT_0; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_689 = 2'h3 == _GEN_239 ? _GEN_625 : PHT_1; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_690 = 2'h3 == _GEN_239 ? _GEN_626 : PHT_2; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_691 = 2'h3 == _GEN_239 ? _GEN_627 : PHT_3; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_692 = 2'h3 == _GEN_239 ? _GEN_628 : PHT_4; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_693 = 2'h3 == _GEN_239 ? _GEN_629 : PHT_5; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_694 = 2'h3 == _GEN_239 ? _GEN_630 : PHT_6; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_695 = 2'h3 == _GEN_239 ? _GEN_631 : PHT_7; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_696 = 2'h3 == _GEN_239 ? _GEN_632 : PHT_8; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_697 = 2'h3 == _GEN_239 ? _GEN_633 : PHT_9; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_698 = 2'h3 == _GEN_239 ? _GEN_634 : PHT_10; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_699 = 2'h3 == _GEN_239 ? _GEN_635 : PHT_11; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_700 = 2'h3 == _GEN_239 ? _GEN_636 : PHT_12; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_701 = 2'h3 == _GEN_239 ? _GEN_637 : PHT_13; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_702 = 2'h3 == _GEN_239 ? _GEN_638 : PHT_14; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_703 = 2'h3 == _GEN_239 ? _GEN_639 : PHT_15; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_704 = 2'h3 == _GEN_239 ? _GEN_640 : PHT_16; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_705 = 2'h3 == _GEN_239 ? _GEN_641 : PHT_17; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_706 = 2'h3 == _GEN_239 ? _GEN_642 : PHT_18; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_707 = 2'h3 == _GEN_239 ? _GEN_643 : PHT_19; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_708 = 2'h3 == _GEN_239 ? _GEN_644 : PHT_20; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_709 = 2'h3 == _GEN_239 ? _GEN_645 : PHT_21; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_710 = 2'h3 == _GEN_239 ? _GEN_646 : PHT_22; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_711 = 2'h3 == _GEN_239 ? _GEN_647 : PHT_23; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_712 = 2'h3 == _GEN_239 ? _GEN_648 : PHT_24; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_713 = 2'h3 == _GEN_239 ? _GEN_649 : PHT_25; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_714 = 2'h3 == _GEN_239 ? _GEN_650 : PHT_26; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_715 = 2'h3 == _GEN_239 ? _GEN_651 : PHT_27; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_716 = 2'h3 == _GEN_239 ? _GEN_652 : PHT_28; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_717 = 2'h3 == _GEN_239 ? _GEN_653 : PHT_29; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_718 = 2'h3 == _GEN_239 ? _GEN_654 : PHT_30; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_719 = 2'h3 == _GEN_239 ? _GEN_655 : PHT_31; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_720 = 2'h3 == _GEN_239 ? _GEN_656 : PHT_32; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_721 = 2'h3 == _GEN_239 ? _GEN_657 : PHT_33; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_722 = 2'h3 == _GEN_239 ? _GEN_658 : PHT_34; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_723 = 2'h3 == _GEN_239 ? _GEN_659 : PHT_35; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_724 = 2'h3 == _GEN_239 ? _GEN_660 : PHT_36; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_725 = 2'h3 == _GEN_239 ? _GEN_661 : PHT_37; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_726 = 2'h3 == _GEN_239 ? _GEN_662 : PHT_38; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_727 = 2'h3 == _GEN_239 ? _GEN_663 : PHT_39; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_728 = 2'h3 == _GEN_239 ? _GEN_664 : PHT_40; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_729 = 2'h3 == _GEN_239 ? _GEN_665 : PHT_41; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_730 = 2'h3 == _GEN_239 ? _GEN_666 : PHT_42; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_731 = 2'h3 == _GEN_239 ? _GEN_667 : PHT_43; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_732 = 2'h3 == _GEN_239 ? _GEN_668 : PHT_44; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_733 = 2'h3 == _GEN_239 ? _GEN_669 : PHT_45; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_734 = 2'h3 == _GEN_239 ? _GEN_670 : PHT_46; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_735 = 2'h3 == _GEN_239 ? _GEN_671 : PHT_47; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_736 = 2'h3 == _GEN_239 ? _GEN_672 : PHT_48; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_737 = 2'h3 == _GEN_239 ? _GEN_673 : PHT_49; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_738 = 2'h3 == _GEN_239 ? _GEN_674 : PHT_50; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_739 = 2'h3 == _GEN_239 ? _GEN_675 : PHT_51; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_740 = 2'h3 == _GEN_239 ? _GEN_676 : PHT_52; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_741 = 2'h3 == _GEN_239 ? _GEN_677 : PHT_53; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_742 = 2'h3 == _GEN_239 ? _GEN_678 : PHT_54; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_743 = 2'h3 == _GEN_239 ? _GEN_679 : PHT_55; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_744 = 2'h3 == _GEN_239 ? _GEN_680 : PHT_56; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_745 = 2'h3 == _GEN_239 ? _GEN_681 : PHT_57; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_746 = 2'h3 == _GEN_239 ? _GEN_682 : PHT_58; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_747 = 2'h3 == _GEN_239 ? _GEN_683 : PHT_59; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_748 = 2'h3 == _GEN_239 ? _GEN_684 : PHT_60; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_749 = 2'h3 == _GEN_239 ? _GEN_685 : PHT_61; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_750 = 2'h3 == _GEN_239 ? _GEN_686 : PHT_62; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_751 = 2'h3 == _GEN_239 ? _GEN_687 : PHT_63; // @[BPU.scala 32:26 45:35]
  wire [1:0] _GEN_752 = 2'h2 == _GEN_239 ? _GEN_496 : _GEN_688; // @[BPU.scala 45:35]
  wire [1:0] _GEN_753 = 2'h2 == _GEN_239 ? _GEN_497 : _GEN_689; // @[BPU.scala 45:35]
  wire [1:0] _GEN_754 = 2'h2 == _GEN_239 ? _GEN_498 : _GEN_690; // @[BPU.scala 45:35]
  wire [1:0] _GEN_755 = 2'h2 == _GEN_239 ? _GEN_499 : _GEN_691; // @[BPU.scala 45:35]
  wire [1:0] _GEN_756 = 2'h2 == _GEN_239 ? _GEN_500 : _GEN_692; // @[BPU.scala 45:35]
  wire [1:0] _GEN_757 = 2'h2 == _GEN_239 ? _GEN_501 : _GEN_693; // @[BPU.scala 45:35]
  wire [1:0] _GEN_758 = 2'h2 == _GEN_239 ? _GEN_502 : _GEN_694; // @[BPU.scala 45:35]
  wire [1:0] _GEN_759 = 2'h2 == _GEN_239 ? _GEN_503 : _GEN_695; // @[BPU.scala 45:35]
  wire [1:0] _GEN_760 = 2'h2 == _GEN_239 ? _GEN_504 : _GEN_696; // @[BPU.scala 45:35]
  wire [1:0] _GEN_761 = 2'h2 == _GEN_239 ? _GEN_505 : _GEN_697; // @[BPU.scala 45:35]
  wire [1:0] _GEN_762 = 2'h2 == _GEN_239 ? _GEN_506 : _GEN_698; // @[BPU.scala 45:35]
  wire [1:0] _GEN_763 = 2'h2 == _GEN_239 ? _GEN_507 : _GEN_699; // @[BPU.scala 45:35]
  wire [1:0] _GEN_764 = 2'h2 == _GEN_239 ? _GEN_508 : _GEN_700; // @[BPU.scala 45:35]
  wire [1:0] _GEN_765 = 2'h2 == _GEN_239 ? _GEN_509 : _GEN_701; // @[BPU.scala 45:35]
  wire [1:0] _GEN_766 = 2'h2 == _GEN_239 ? _GEN_510 : _GEN_702; // @[BPU.scala 45:35]
  wire [1:0] _GEN_767 = 2'h2 == _GEN_239 ? _GEN_511 : _GEN_703; // @[BPU.scala 45:35]
  wire [1:0] _GEN_768 = 2'h2 == _GEN_239 ? _GEN_512 : _GEN_704; // @[BPU.scala 45:35]
  wire [1:0] _GEN_769 = 2'h2 == _GEN_239 ? _GEN_513 : _GEN_705; // @[BPU.scala 45:35]
  wire [1:0] _GEN_770 = 2'h2 == _GEN_239 ? _GEN_514 : _GEN_706; // @[BPU.scala 45:35]
  wire [1:0] _GEN_771 = 2'h2 == _GEN_239 ? _GEN_515 : _GEN_707; // @[BPU.scala 45:35]
  wire [1:0] _GEN_772 = 2'h2 == _GEN_239 ? _GEN_516 : _GEN_708; // @[BPU.scala 45:35]
  wire [1:0] _GEN_773 = 2'h2 == _GEN_239 ? _GEN_517 : _GEN_709; // @[BPU.scala 45:35]
  wire [1:0] _GEN_774 = 2'h2 == _GEN_239 ? _GEN_518 : _GEN_710; // @[BPU.scala 45:35]
  wire [1:0] _GEN_775 = 2'h2 == _GEN_239 ? _GEN_519 : _GEN_711; // @[BPU.scala 45:35]
  wire [1:0] _GEN_776 = 2'h2 == _GEN_239 ? _GEN_520 : _GEN_712; // @[BPU.scala 45:35]
  wire [1:0] _GEN_777 = 2'h2 == _GEN_239 ? _GEN_521 : _GEN_713; // @[BPU.scala 45:35]
  wire [1:0] _GEN_778 = 2'h2 == _GEN_239 ? _GEN_522 : _GEN_714; // @[BPU.scala 45:35]
  wire [1:0] _GEN_779 = 2'h2 == _GEN_239 ? _GEN_523 : _GEN_715; // @[BPU.scala 45:35]
  wire [1:0] _GEN_780 = 2'h2 == _GEN_239 ? _GEN_524 : _GEN_716; // @[BPU.scala 45:35]
  wire [1:0] _GEN_781 = 2'h2 == _GEN_239 ? _GEN_525 : _GEN_717; // @[BPU.scala 45:35]
  wire [1:0] _GEN_782 = 2'h2 == _GEN_239 ? _GEN_526 : _GEN_718; // @[BPU.scala 45:35]
  wire [1:0] _GEN_783 = 2'h2 == _GEN_239 ? _GEN_527 : _GEN_719; // @[BPU.scala 45:35]
  wire [1:0] _GEN_784 = 2'h2 == _GEN_239 ? _GEN_528 : _GEN_720; // @[BPU.scala 45:35]
  wire [1:0] _GEN_785 = 2'h2 == _GEN_239 ? _GEN_529 : _GEN_721; // @[BPU.scala 45:35]
  wire [1:0] _GEN_786 = 2'h2 == _GEN_239 ? _GEN_530 : _GEN_722; // @[BPU.scala 45:35]
  wire [1:0] _GEN_787 = 2'h2 == _GEN_239 ? _GEN_531 : _GEN_723; // @[BPU.scala 45:35]
  wire [1:0] _GEN_788 = 2'h2 == _GEN_239 ? _GEN_532 : _GEN_724; // @[BPU.scala 45:35]
  wire [1:0] _GEN_789 = 2'h2 == _GEN_239 ? _GEN_533 : _GEN_725; // @[BPU.scala 45:35]
  wire [1:0] _GEN_790 = 2'h2 == _GEN_239 ? _GEN_534 : _GEN_726; // @[BPU.scala 45:35]
  wire [1:0] _GEN_791 = 2'h2 == _GEN_239 ? _GEN_535 : _GEN_727; // @[BPU.scala 45:35]
  wire [1:0] _GEN_792 = 2'h2 == _GEN_239 ? _GEN_536 : _GEN_728; // @[BPU.scala 45:35]
  wire [1:0] _GEN_793 = 2'h2 == _GEN_239 ? _GEN_537 : _GEN_729; // @[BPU.scala 45:35]
  wire [1:0] _GEN_794 = 2'h2 == _GEN_239 ? _GEN_538 : _GEN_730; // @[BPU.scala 45:35]
  wire [1:0] _GEN_795 = 2'h2 == _GEN_239 ? _GEN_539 : _GEN_731; // @[BPU.scala 45:35]
  wire [1:0] _GEN_796 = 2'h2 == _GEN_239 ? _GEN_540 : _GEN_732; // @[BPU.scala 45:35]
  wire [1:0] _GEN_797 = 2'h2 == _GEN_239 ? _GEN_541 : _GEN_733; // @[BPU.scala 45:35]
  wire [1:0] _GEN_798 = 2'h2 == _GEN_239 ? _GEN_542 : _GEN_734; // @[BPU.scala 45:35]
  wire [1:0] _GEN_799 = 2'h2 == _GEN_239 ? _GEN_543 : _GEN_735; // @[BPU.scala 45:35]
  wire [1:0] _GEN_800 = 2'h2 == _GEN_239 ? _GEN_544 : _GEN_736; // @[BPU.scala 45:35]
  wire [1:0] _GEN_801 = 2'h2 == _GEN_239 ? _GEN_545 : _GEN_737; // @[BPU.scala 45:35]
  wire [1:0] _GEN_802 = 2'h2 == _GEN_239 ? _GEN_546 : _GEN_738; // @[BPU.scala 45:35]
  wire [1:0] _GEN_803 = 2'h2 == _GEN_239 ? _GEN_547 : _GEN_739; // @[BPU.scala 45:35]
  wire [1:0] _GEN_804 = 2'h2 == _GEN_239 ? _GEN_548 : _GEN_740; // @[BPU.scala 45:35]
  wire [1:0] _GEN_805 = 2'h2 == _GEN_239 ? _GEN_549 : _GEN_741; // @[BPU.scala 45:35]
  wire [1:0] _GEN_806 = 2'h2 == _GEN_239 ? _GEN_550 : _GEN_742; // @[BPU.scala 45:35]
  wire [1:0] _GEN_807 = 2'h2 == _GEN_239 ? _GEN_551 : _GEN_743; // @[BPU.scala 45:35]
  wire [1:0] _GEN_808 = 2'h2 == _GEN_239 ? _GEN_552 : _GEN_744; // @[BPU.scala 45:35]
  wire [1:0] _GEN_809 = 2'h2 == _GEN_239 ? _GEN_553 : _GEN_745; // @[BPU.scala 45:35]
  wire [1:0] _GEN_810 = 2'h2 == _GEN_239 ? _GEN_554 : _GEN_746; // @[BPU.scala 45:35]
  wire [1:0] _GEN_811 = 2'h2 == _GEN_239 ? _GEN_555 : _GEN_747; // @[BPU.scala 45:35]
  wire [1:0] _GEN_812 = 2'h2 == _GEN_239 ? _GEN_556 : _GEN_748; // @[BPU.scala 45:35]
  wire [1:0] _GEN_813 = 2'h2 == _GEN_239 ? _GEN_557 : _GEN_749; // @[BPU.scala 45:35]
  wire [1:0] _GEN_814 = 2'h2 == _GEN_239 ? _GEN_558 : _GEN_750; // @[BPU.scala 45:35]
  wire [1:0] _GEN_815 = 2'h2 == _GEN_239 ? _GEN_559 : _GEN_751; // @[BPU.scala 45:35]
  assign io_branchD = io_instrD[31:26] == 6'h1 & io_instrD[19:17] == 3'h0 | io_instrD[31:28] == 4'h1; // @[BPU.scala 22:74]
  assign io_pred_takeD = io_enaD & io_branchD & (_GEN_79 == 2'h2 | _GEN_79 == 2'h3); // @[BPU.scala 37:42]
  assign io_branch_targetD = io_pc_plus4D + _io_branch_targetD_T_4; // @[BPU.scala 23:37]
  always @(posedge clock) begin
    if (reset) begin // @[BPU.scala 31:26]
      BHT_0 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h0 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_0 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_1 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h1 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_1 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_2 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h2 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_2 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_3 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h3 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_3 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_4 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h4 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_4 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_5 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h5 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_5 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_6 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h6 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_6 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_7 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h7 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_7 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_8 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h8 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_8 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_9 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'h9 == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_9 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_10 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'ha == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_10 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_11 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'hb == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_11 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_12 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'hc == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_12 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_13 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'hd == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_13 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_14 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'he == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_14 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 31:26]
      BHT_15 <= 6'h0; // @[BPU.scala 31:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (4'hf == update_BHT_index) begin // @[BPU.scala 44:27]
        BHT_15 <= _BHT_T_1; // @[BPU.scala 44:27]
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_0 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h0 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_0 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_0 <= _GEN_368;
      end else begin
        PHT_0 <= _GEN_752;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_1 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h1 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_1 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_1 <= _GEN_369;
      end else begin
        PHT_1 <= _GEN_753;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_2 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h2 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_2 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_2 <= _GEN_370;
      end else begin
        PHT_2 <= _GEN_754;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_3 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h3 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_3 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_3 <= _GEN_371;
      end else begin
        PHT_3 <= _GEN_755;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_4 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h4 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_4 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_4 <= _GEN_372;
      end else begin
        PHT_4 <= _GEN_756;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_5 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h5 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_5 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_5 <= _GEN_373;
      end else begin
        PHT_5 <= _GEN_757;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_6 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h6 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_6 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_6 <= _GEN_374;
      end else begin
        PHT_6 <= _GEN_758;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_7 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h7 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_7 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_7 <= _GEN_375;
      end else begin
        PHT_7 <= _GEN_759;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_8 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h8 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_8 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_8 <= _GEN_376;
      end else begin
        PHT_8 <= _GEN_760;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_9 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h9 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_9 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_9 <= _GEN_377;
      end else begin
        PHT_9 <= _GEN_761;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_10 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'ha == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_10 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_10 <= _GEN_378;
      end else begin
        PHT_10 <= _GEN_762;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_11 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'hb == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_11 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_11 <= _GEN_379;
      end else begin
        PHT_11 <= _GEN_763;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_12 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'hc == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_12 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_12 <= _GEN_380;
      end else begin
        PHT_12 <= _GEN_764;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_13 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'hd == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_13 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_13 <= _GEN_381;
      end else begin
        PHT_13 <= _GEN_765;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_14 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'he == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_14 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_14 <= _GEN_382;
      end else begin
        PHT_14 <= _GEN_766;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_15 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'hf == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_15 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_15 <= _GEN_383;
      end else begin
        PHT_15 <= _GEN_767;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_16 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h10 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_16 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_16 <= _GEN_384;
      end else begin
        PHT_16 <= _GEN_768;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_17 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h11 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_17 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_17 <= _GEN_385;
      end else begin
        PHT_17 <= _GEN_769;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_18 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h12 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_18 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_18 <= _GEN_386;
      end else begin
        PHT_18 <= _GEN_770;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_19 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h13 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_19 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_19 <= _GEN_387;
      end else begin
        PHT_19 <= _GEN_771;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_20 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h14 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_20 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_20 <= _GEN_388;
      end else begin
        PHT_20 <= _GEN_772;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_21 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h15 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_21 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_21 <= _GEN_389;
      end else begin
        PHT_21 <= _GEN_773;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_22 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h16 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_22 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_22 <= _GEN_390;
      end else begin
        PHT_22 <= _GEN_774;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_23 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h17 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_23 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_23 <= _GEN_391;
      end else begin
        PHT_23 <= _GEN_775;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_24 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h18 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_24 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_24 <= _GEN_392;
      end else begin
        PHT_24 <= _GEN_776;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_25 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h19 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_25 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_25 <= _GEN_393;
      end else begin
        PHT_25 <= _GEN_777;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_26 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h1a == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_26 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_26 <= _GEN_394;
      end else begin
        PHT_26 <= _GEN_778;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_27 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h1b == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_27 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_27 <= _GEN_395;
      end else begin
        PHT_27 <= _GEN_779;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_28 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h1c == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_28 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_28 <= _GEN_396;
      end else begin
        PHT_28 <= _GEN_780;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_29 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h1d == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_29 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_29 <= _GEN_397;
      end else begin
        PHT_29 <= _GEN_781;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_30 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h1e == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_30 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_30 <= _GEN_398;
      end else begin
        PHT_30 <= _GEN_782;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_31 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h1f == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_31 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_31 <= _GEN_399;
      end else begin
        PHT_31 <= _GEN_783;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_32 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h20 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_32 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_32 <= _GEN_400;
      end else begin
        PHT_32 <= _GEN_784;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_33 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h21 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_33 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_33 <= _GEN_401;
      end else begin
        PHT_33 <= _GEN_785;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_34 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h22 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_34 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_34 <= _GEN_402;
      end else begin
        PHT_34 <= _GEN_786;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_35 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h23 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_35 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_35 <= _GEN_403;
      end else begin
        PHT_35 <= _GEN_787;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_36 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h24 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_36 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_36 <= _GEN_404;
      end else begin
        PHT_36 <= _GEN_788;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_37 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h25 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_37 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_37 <= _GEN_405;
      end else begin
        PHT_37 <= _GEN_789;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_38 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h26 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_38 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_38 <= _GEN_406;
      end else begin
        PHT_38 <= _GEN_790;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_39 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h27 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_39 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_39 <= _GEN_407;
      end else begin
        PHT_39 <= _GEN_791;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_40 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h28 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_40 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_40 <= _GEN_408;
      end else begin
        PHT_40 <= _GEN_792;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_41 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h29 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_41 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_41 <= _GEN_409;
      end else begin
        PHT_41 <= _GEN_793;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_42 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h2a == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_42 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_42 <= _GEN_410;
      end else begin
        PHT_42 <= _GEN_794;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_43 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h2b == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_43 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_43 <= _GEN_411;
      end else begin
        PHT_43 <= _GEN_795;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_44 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h2c == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_44 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_44 <= _GEN_412;
      end else begin
        PHT_44 <= _GEN_796;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_45 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h2d == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_45 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_45 <= _GEN_413;
      end else begin
        PHT_45 <= _GEN_797;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_46 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h2e == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_46 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_46 <= _GEN_414;
      end else begin
        PHT_46 <= _GEN_798;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_47 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h2f == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_47 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_47 <= _GEN_415;
      end else begin
        PHT_47 <= _GEN_799;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_48 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h30 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_48 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_48 <= _GEN_416;
      end else begin
        PHT_48 <= _GEN_800;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_49 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h31 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_49 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_49 <= _GEN_417;
      end else begin
        PHT_49 <= _GEN_801;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_50 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h32 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_50 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_50 <= _GEN_418;
      end else begin
        PHT_50 <= _GEN_802;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_51 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h33 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_51 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_51 <= _GEN_419;
      end else begin
        PHT_51 <= _GEN_803;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_52 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h34 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_52 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_52 <= _GEN_420;
      end else begin
        PHT_52 <= _GEN_804;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_53 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h35 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_53 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_53 <= _GEN_421;
      end else begin
        PHT_53 <= _GEN_805;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_54 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h36 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_54 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_54 <= _GEN_422;
      end else begin
        PHT_54 <= _GEN_806;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_55 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h37 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_55 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_55 <= _GEN_423;
      end else begin
        PHT_55 <= _GEN_807;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_56 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h38 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_56 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_56 <= _GEN_424;
      end else begin
        PHT_56 <= _GEN_808;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_57 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h39 == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_57 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_57 <= _GEN_425;
      end else begin
        PHT_57 <= _GEN_809;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_58 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h3a == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_58 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_58 <= _GEN_426;
      end else begin
        PHT_58 <= _GEN_810;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_59 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h3b == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_59 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_59 <= _GEN_427;
      end else begin
        PHT_59 <= _GEN_811;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_60 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h3c == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_60 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_60 <= _GEN_428;
      end else begin
        PHT_60 <= _GEN_812;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_61 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h3d == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_61 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_61 <= _GEN_429;
      end else begin
        PHT_61 <= _GEN_813;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_62 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h3e == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_62 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_62 <= _GEN_430;
      end else begin
        PHT_62 <= _GEN_814;
      end
    end
    if (reset) begin // @[BPU.scala 32:26]
      PHT_63 <= 2'h0; // @[BPU.scala 32:26]
    end else if (io_branchE) begin // @[BPU.scala 43:20]
      if (2'h0 == _GEN_239) begin // @[BPU.scala 45:35]
        if (6'h3f == _GEN_159) begin // @[BPU.scala 47:31]
          PHT_63 <= _PHT_T; // @[BPU.scala 47:31]
        end
      end else if (2'h1 == _GEN_239) begin // @[BPU.scala 45:35]
        PHT_63 <= _GEN_431;
      end else begin
        PHT_63 <= _GEN_815;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  BHT_0 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  BHT_1 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  BHT_2 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  BHT_3 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  BHT_4 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  BHT_5 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  BHT_6 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  BHT_7 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  BHT_8 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  BHT_9 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  BHT_10 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  BHT_11 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  BHT_12 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  BHT_13 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  BHT_14 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  BHT_15 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  PHT_0 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  PHT_1 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  PHT_2 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  PHT_3 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  PHT_4 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  PHT_5 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  PHT_6 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  PHT_7 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  PHT_8 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  PHT_9 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  PHT_10 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  PHT_11 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  PHT_12 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  PHT_13 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  PHT_14 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  PHT_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  PHT_16 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  PHT_17 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  PHT_18 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  PHT_19 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  PHT_20 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  PHT_21 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  PHT_22 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  PHT_23 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  PHT_24 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  PHT_25 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  PHT_26 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  PHT_27 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  PHT_28 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  PHT_29 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  PHT_30 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  PHT_31 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  PHT_32 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  PHT_33 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  PHT_34 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  PHT_35 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  PHT_36 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  PHT_37 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  PHT_38 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  PHT_39 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  PHT_40 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  PHT_41 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  PHT_42 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  PHT_43 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  PHT_44 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  PHT_45 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  PHT_46 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  PHT_47 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  PHT_48 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  PHT_49 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  PHT_50 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  PHT_51 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  PHT_52 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  PHT_53 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  PHT_54 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  PHT_55 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  PHT_56 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  PHT_57 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  PHT_58 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  PHT_59 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  PHT_60 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  PHT_61 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  PHT_62 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  PHT_63 = _RAND_79[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstBuffer(
  input         clock,
  input         reset,
  input         io_fifo_rst,
  input         io_flush_delay_slot,
  input         io_delay_sel_rst,
  input         io_D_delay_rst,
  input         io_E_delay_rst,
  input         io_i_stall,
  input         io_master_is_branch,
  output        io_master_is_in_delayslot_o,
  input         io_read_en_0,
  input         io_read_en_1,
  output        io_read_0_tlb_invalid,
  output [31:0] io_read_0_data,
  output [31:0] io_read_0_addr,
  output        io_read_1_tlb_invalid,
  output [31:0] io_read_1_data,
  output [31:0] io_read_1_addr,
  input         io_write_en_0,
  input         io_write_en_1,
  input         io_write_0_tlb_invalid,
  input  [31:0] io_write_0_data,
  input  [31:0] io_write_0_addr,
  input         io_write_1_tlb_invalid,
  input  [31:0] io_write_1_data,
  input  [31:0] io_write_1_addr,
  output        io_empty,
  output        io_almost_empty,
  output        io_full
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
`endif // RANDOMIZE_REG_INIT
  reg  buffer_0_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_0_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_0_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_1_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_1_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_1_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_2_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_2_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_2_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_3_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_3_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_3_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_4_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_4_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_4_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_5_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_5_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_5_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_6_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_6_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_6_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_7_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_7_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_7_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_8_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_8_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_8_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_9_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_9_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_9_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_10_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_10_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_10_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_11_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_11_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_11_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_12_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_12_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_12_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_13_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_13_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_13_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_14_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_14_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_14_addr; // @[InstBuffer.scala 41:23]
  reg  buffer_15_tlb_invalid; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_15_data; // @[InstBuffer.scala 41:23]
  reg [31:0] buffer_15_addr; // @[InstBuffer.scala 41:23]
  reg [3:0] enq_ptr; // @[InstBuffer.scala 44:24]
  reg [3:0] deq_ptr; // @[InstBuffer.scala 45:24]
  wire [3:0] _count_T_1 = enq_ptr - deq_ptr; // @[InstBuffer.scala 46:29]
  wire [4:0] _GEN_477 = {{1'd0}, _count_T_1}; // @[InstBuffer.scala 46:64]
  reg  master_is_in_delayslot; // @[InstBuffer.scala 54:39]
  wire  _master_is_in_delayslot_T = ~io_read_en_0; // @[InstBuffer.scala 60:7]
  wire  _master_is_in_delayslot_T_2 = io_master_is_branch & ~io_read_en_1; // @[InstBuffer.scala 61:28]
  reg  delayslot_stall; // @[InstBuffer.scala 65:33]
  reg  delayslot_enable; // @[InstBuffer.scala 66:33]
  reg  delayslot_line_tlb_invalid; // @[InstBuffer.scala 67:33]
  reg [31:0] delayslot_line_data; // @[InstBuffer.scala 67:33]
  reg [31:0] delayslot_line_addr; // @[InstBuffer.scala 67:33]
  wire  _T_1 = ~io_flush_delay_slot; // @[InstBuffer.scala 69:40]
  wire [3:0] _T_5 = deq_ptr + 4'h1; // @[InstBuffer.scala 69:87]
  wire  _T_6 = _T_5 == enq_ptr; // @[InstBuffer.scala 69:93]
  wire  _T_7 = deq_ptr == enq_ptr; // @[InstBuffer.scala 69:116]
  wire  _T_9 = io_fifo_rst & io_delay_sel_rst & ~io_flush_delay_slot & io_i_stall & (_T_5 == enq_ptr | deq_ptr ==
    enq_ptr); // @[InstBuffer.scala 69:75]
  wire  _GEN_0 = delayslot_stall & io_write_en_0 ? 1'h0 : delayslot_stall; // @[InstBuffer.scala 72:49 73:21 65:33]
  wire  _GEN_1 = _T_9 | _GEN_0; // @[InstBuffer.scala 70:5 71:21]
  wire  _GEN_7 = 4'h1 == deq_ptr ? buffer_1_tlb_invalid : buffer_0_tlb_invalid; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_8 = 4'h1 == deq_ptr ? buffer_1_data : buffer_0_data; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_9 = 4'h1 == deq_ptr ? buffer_1_addr : buffer_0_addr; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_11 = 4'h2 == deq_ptr ? buffer_2_tlb_invalid : _GEN_7; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_12 = 4'h2 == deq_ptr ? buffer_2_data : _GEN_8; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_13 = 4'h2 == deq_ptr ? buffer_2_addr : _GEN_9; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_15 = 4'h3 == deq_ptr ? buffer_3_tlb_invalid : _GEN_11; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_16 = 4'h3 == deq_ptr ? buffer_3_data : _GEN_12; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_17 = 4'h3 == deq_ptr ? buffer_3_addr : _GEN_13; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_19 = 4'h4 == deq_ptr ? buffer_4_tlb_invalid : _GEN_15; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_20 = 4'h4 == deq_ptr ? buffer_4_data : _GEN_16; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_21 = 4'h4 == deq_ptr ? buffer_4_addr : _GEN_17; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_23 = 4'h5 == deq_ptr ? buffer_5_tlb_invalid : _GEN_19; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_24 = 4'h5 == deq_ptr ? buffer_5_data : _GEN_20; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_25 = 4'h5 == deq_ptr ? buffer_5_addr : _GEN_21; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_27 = 4'h6 == deq_ptr ? buffer_6_tlb_invalid : _GEN_23; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_28 = 4'h6 == deq_ptr ? buffer_6_data : _GEN_24; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_29 = 4'h6 == deq_ptr ? buffer_6_addr : _GEN_25; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_31 = 4'h7 == deq_ptr ? buffer_7_tlb_invalid : _GEN_27; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_32 = 4'h7 == deq_ptr ? buffer_7_data : _GEN_28; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_33 = 4'h7 == deq_ptr ? buffer_7_addr : _GEN_29; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_35 = 4'h8 == deq_ptr ? buffer_8_tlb_invalid : _GEN_31; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_36 = 4'h8 == deq_ptr ? buffer_8_data : _GEN_32; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_37 = 4'h8 == deq_ptr ? buffer_8_addr : _GEN_33; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_39 = 4'h9 == deq_ptr ? buffer_9_tlb_invalid : _GEN_35; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_40 = 4'h9 == deq_ptr ? buffer_9_data : _GEN_36; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_41 = 4'h9 == deq_ptr ? buffer_9_addr : _GEN_37; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_43 = 4'ha == deq_ptr ? buffer_10_tlb_invalid : _GEN_39; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_44 = 4'ha == deq_ptr ? buffer_10_data : _GEN_40; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_45 = 4'ha == deq_ptr ? buffer_10_addr : _GEN_41; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_47 = 4'hb == deq_ptr ? buffer_11_tlb_invalid : _GEN_43; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_48 = 4'hb == deq_ptr ? buffer_11_data : _GEN_44; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_49 = 4'hb == deq_ptr ? buffer_11_addr : _GEN_45; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_51 = 4'hc == deq_ptr ? buffer_12_tlb_invalid : _GEN_47; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_52 = 4'hc == deq_ptr ? buffer_12_data : _GEN_48; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_53 = 4'hc == deq_ptr ? buffer_12_addr : _GEN_49; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_55 = 4'hd == deq_ptr ? buffer_13_tlb_invalid : _GEN_51; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_56 = 4'hd == deq_ptr ? buffer_13_data : _GEN_52; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_57 = 4'hd == deq_ptr ? buffer_13_addr : _GEN_53; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_59 = 4'he == deq_ptr ? buffer_14_tlb_invalid : _GEN_55; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_60 = 4'he == deq_ptr ? buffer_14_data : _GEN_56; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_61 = 4'he == deq_ptr ? buffer_14_addr : _GEN_57; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_63 = 4'hf == deq_ptr ? buffer_15_tlb_invalid : _GEN_59; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_64 = 4'hf == deq_ptr ? buffer_15_data : _GEN_60; // @[InstBuffer.scala 79:{30,30}]
  wire [31:0] _GEN_65 = 4'hf == deq_ptr ? buffer_15_addr : _GEN_61; // @[InstBuffer.scala 79:{30,30}]
  wire  _GEN_71 = 4'h1 == _T_5 ? buffer_1_tlb_invalid : buffer_0_tlb_invalid; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_72 = 4'h1 == _T_5 ? buffer_1_data : buffer_0_data; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_73 = 4'h1 == _T_5 ? buffer_1_addr : buffer_0_addr; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_75 = 4'h2 == _T_5 ? buffer_2_tlb_invalid : _GEN_71; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_76 = 4'h2 == _T_5 ? buffer_2_data : _GEN_72; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_77 = 4'h2 == _T_5 ? buffer_2_addr : _GEN_73; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_79 = 4'h3 == _T_5 ? buffer_3_tlb_invalid : _GEN_75; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_80 = 4'h3 == _T_5 ? buffer_3_data : _GEN_76; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_81 = 4'h3 == _T_5 ? buffer_3_addr : _GEN_77; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_83 = 4'h4 == _T_5 ? buffer_4_tlb_invalid : _GEN_79; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_84 = 4'h4 == _T_5 ? buffer_4_data : _GEN_80; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_85 = 4'h4 == _T_5 ? buffer_4_addr : _GEN_81; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_87 = 4'h5 == _T_5 ? buffer_5_tlb_invalid : _GEN_83; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_88 = 4'h5 == _T_5 ? buffer_5_data : _GEN_84; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_89 = 4'h5 == _T_5 ? buffer_5_addr : _GEN_85; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_91 = 4'h6 == _T_5 ? buffer_6_tlb_invalid : _GEN_87; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_92 = 4'h6 == _T_5 ? buffer_6_data : _GEN_88; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_93 = 4'h6 == _T_5 ? buffer_6_addr : _GEN_89; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_95 = 4'h7 == _T_5 ? buffer_7_tlb_invalid : _GEN_91; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_96 = 4'h7 == _T_5 ? buffer_7_data : _GEN_92; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_97 = 4'h7 == _T_5 ? buffer_7_addr : _GEN_93; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_99 = 4'h8 == _T_5 ? buffer_8_tlb_invalid : _GEN_95; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_100 = 4'h8 == _T_5 ? buffer_8_data : _GEN_96; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_101 = 4'h8 == _T_5 ? buffer_8_addr : _GEN_97; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_103 = 4'h9 == _T_5 ? buffer_9_tlb_invalid : _GEN_99; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_104 = 4'h9 == _T_5 ? buffer_9_data : _GEN_100; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_105 = 4'h9 == _T_5 ? buffer_9_addr : _GEN_101; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_107 = 4'ha == _T_5 ? buffer_10_tlb_invalid : _GEN_103; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_108 = 4'ha == _T_5 ? buffer_10_data : _GEN_104; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_109 = 4'ha == _T_5 ? buffer_10_addr : _GEN_105; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_111 = 4'hb == _T_5 ? buffer_11_tlb_invalid : _GEN_107; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_112 = 4'hb == _T_5 ? buffer_11_data : _GEN_108; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_113 = 4'hb == _T_5 ? buffer_11_addr : _GEN_109; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_115 = 4'hc == _T_5 ? buffer_12_tlb_invalid : _GEN_111; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_116 = 4'hc == _T_5 ? buffer_12_data : _GEN_112; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_117 = 4'hc == _T_5 ? buffer_12_addr : _GEN_113; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_119 = 4'hd == _T_5 ? buffer_13_tlb_invalid : _GEN_115; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_120 = 4'hd == _T_5 ? buffer_13_data : _GEN_116; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_121 = 4'hd == _T_5 ? buffer_13_addr : _GEN_117; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_123 = 4'he == _T_5 ? buffer_14_tlb_invalid : _GEN_119; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_124 = 4'he == _T_5 ? buffer_14_data : _GEN_120; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_125 = 4'he == _T_5 ? buffer_14_addr : _GEN_121; // @[InstBuffer.scala 82:{28,28}]
  wire  _GEN_127 = 4'hf == _T_5 ? buffer_15_tlb_invalid : _GEN_123; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_128 = 4'hf == _T_5 ? buffer_15_data : _GEN_124; // @[InstBuffer.scala 82:{28,28}]
  wire [31:0] _GEN_129 = 4'hf == _T_5 ? buffer_15_addr : _GEN_125; // @[InstBuffer.scala 82:{28,28}]
  wire  _delayslot_line_T_7_tlb_invalid = _T_6 ? io_write_0_tlb_invalid : _GEN_127; // @[InstBuffer.scala 82:28]
  wire [31:0] _delayslot_line_T_7_data = _T_6 ? io_write_0_data : _GEN_128; // @[InstBuffer.scala 82:28]
  wire [31:0] _delayslot_line_T_7_addr = _T_6 ? io_write_0_addr : _GEN_129; // @[InstBuffer.scala 82:28]
  wire  _GEN_132 = io_D_delay_rst & _delayslot_line_T_7_tlb_invalid; // @[InstBuffer.scala 80:32 82:22 89:24]
  wire  _GEN_135 = io_E_delay_rst | io_D_delay_rst; // @[InstBuffer.scala 77:26 78:24]
  wire  _io_read_0_T_1_tlb_invalid = io_empty ? 1'h0 : _GEN_63; // @[Mux.scala 101:16]
  wire [31:0] _io_read_0_T_1_data = io_empty ? 32'h0 : _GEN_64; // @[Mux.scala 101:16]
  wire [31:0] _io_read_0_T_1_addr = io_empty ? 32'h0 : _GEN_65; // @[Mux.scala 101:16]
  wire  _io_read_1_T_2_tlb_invalid = io_almost_empty ? 1'h0 : _GEN_127; // @[Mux.scala 101:16]
  wire [31:0] _io_read_1_T_2_data = io_almost_empty ? 32'h0 : _GEN_128; // @[Mux.scala 101:16]
  wire [31:0] _io_read_1_T_2_addr = io_almost_empty ? 32'h0 : _GEN_129; // @[Mux.scala 101:16]
  wire  _io_read_1_T_3_tlb_invalid = io_empty ? 1'h0 : _io_read_1_T_2_tlb_invalid; // @[Mux.scala 101:16]
  wire [31:0] _io_read_1_T_3_data = io_empty ? 32'h0 : _io_read_1_T_2_data; // @[Mux.scala 101:16]
  wire [31:0] _io_read_1_T_3_addr = io_empty ? 32'h0 : _io_read_1_T_2_addr; // @[Mux.scala 101:16]
  wire [3:0] _deq_ptr_T_1 = deq_ptr + 4'h2; // @[InstBuffer.scala 118:24]
  wire [3:0] _GEN_214 = io_read_en_0 ? _T_5 : deq_ptr; // @[InstBuffer.scala 119:29 120:13 45:24]
  wire [4:0] _T_18 = {{1'd0}, enq_ptr}; // @[InstBuffer.scala 124:70]
  wire  _GEN_234 = 4'h0 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_0_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_235 = 4'h1 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_1_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_236 = 4'h2 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_2_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_237 = 4'h3 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_3_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_238 = 4'h4 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_4_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_239 = 4'h5 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_5_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_240 = 4'h6 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_6_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_241 = 4'h7 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_7_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_242 = 4'h8 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_8_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_243 = 4'h9 == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_9_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_244 = 4'ha == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_10_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_245 = 4'hb == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_11_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_246 = 4'hc == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_12_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_247 = 4'hd == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_13_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_248 = 4'he == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_14_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_249 = 4'hf == _T_18[3:0] ? io_write_0_tlb_invalid : buffer_15_tlb_invalid; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_250 = 4'h0 == _T_18[3:0] ? io_write_0_data : buffer_0_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_251 = 4'h1 == _T_18[3:0] ? io_write_0_data : buffer_1_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_252 = 4'h2 == _T_18[3:0] ? io_write_0_data : buffer_2_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_253 = 4'h3 == _T_18[3:0] ? io_write_0_data : buffer_3_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_254 = 4'h4 == _T_18[3:0] ? io_write_0_data : buffer_4_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_255 = 4'h5 == _T_18[3:0] ? io_write_0_data : buffer_5_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_256 = 4'h6 == _T_18[3:0] ? io_write_0_data : buffer_6_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_257 = 4'h7 == _T_18[3:0] ? io_write_0_data : buffer_7_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_258 = 4'h8 == _T_18[3:0] ? io_write_0_data : buffer_8_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_259 = 4'h9 == _T_18[3:0] ? io_write_0_data : buffer_9_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_260 = 4'ha == _T_18[3:0] ? io_write_0_data : buffer_10_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_261 = 4'hb == _T_18[3:0] ? io_write_0_data : buffer_11_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_262 = 4'hc == _T_18[3:0] ? io_write_0_data : buffer_12_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_263 = 4'hd == _T_18[3:0] ? io_write_0_data : buffer_13_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_264 = 4'he == _T_18[3:0] ? io_write_0_data : buffer_14_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_265 = 4'hf == _T_18[3:0] ? io_write_0_data : buffer_15_data; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_266 = 4'h0 == _T_18[3:0] ? io_write_0_addr : buffer_0_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_267 = 4'h1 == _T_18[3:0] ? io_write_0_addr : buffer_1_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_268 = 4'h2 == _T_18[3:0] ? io_write_0_addr : buffer_2_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_269 = 4'h3 == _T_18[3:0] ? io_write_0_addr : buffer_3_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_270 = 4'h4 == _T_18[3:0] ? io_write_0_addr : buffer_4_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_271 = 4'h5 == _T_18[3:0] ? io_write_0_addr : buffer_5_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_272 = 4'h6 == _T_18[3:0] ? io_write_0_addr : buffer_6_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_273 = 4'h7 == _T_18[3:0] ? io_write_0_addr : buffer_7_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_274 = 4'h8 == _T_18[3:0] ? io_write_0_addr : buffer_8_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_275 = 4'h9 == _T_18[3:0] ? io_write_0_addr : buffer_9_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_276 = 4'ha == _T_18[3:0] ? io_write_0_addr : buffer_10_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_277 = 4'hb == _T_18[3:0] ? io_write_0_addr : buffer_11_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_278 = 4'hc == _T_18[3:0] ? io_write_0_addr : buffer_12_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_279 = 4'hd == _T_18[3:0] ? io_write_0_addr : buffer_13_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_280 = 4'he == _T_18[3:0] ? io_write_0_addr : buffer_14_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire [31:0] _GEN_281 = 4'hf == _T_18[3:0] ? io_write_0_addr : buffer_15_addr; // @[InstBuffer.scala 124:{77,77} 41:23]
  wire  _GEN_298 = io_write_en_0 ? _GEN_234 : buffer_0_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_299 = io_write_en_0 ? _GEN_235 : buffer_1_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_300 = io_write_en_0 ? _GEN_236 : buffer_2_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_301 = io_write_en_0 ? _GEN_237 : buffer_3_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_302 = io_write_en_0 ? _GEN_238 : buffer_4_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_303 = io_write_en_0 ? _GEN_239 : buffer_5_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_304 = io_write_en_0 ? _GEN_240 : buffer_6_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_305 = io_write_en_0 ? _GEN_241 : buffer_7_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_306 = io_write_en_0 ? _GEN_242 : buffer_8_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_307 = io_write_en_0 ? _GEN_243 : buffer_9_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_308 = io_write_en_0 ? _GEN_244 : buffer_10_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_309 = io_write_en_0 ? _GEN_245 : buffer_11_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_310 = io_write_en_0 ? _GEN_246 : buffer_12_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_311 = io_write_en_0 ? _GEN_247 : buffer_13_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_312 = io_write_en_0 ? _GEN_248 : buffer_14_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire  _GEN_313 = io_write_en_0 ? _GEN_249 : buffer_15_tlb_invalid; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_314 = io_write_en_0 ? _GEN_250 : buffer_0_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_315 = io_write_en_0 ? _GEN_251 : buffer_1_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_316 = io_write_en_0 ? _GEN_252 : buffer_2_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_317 = io_write_en_0 ? _GEN_253 : buffer_3_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_318 = io_write_en_0 ? _GEN_254 : buffer_4_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_319 = io_write_en_0 ? _GEN_255 : buffer_5_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_320 = io_write_en_0 ? _GEN_256 : buffer_6_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_321 = io_write_en_0 ? _GEN_257 : buffer_7_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_322 = io_write_en_0 ? _GEN_258 : buffer_8_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_323 = io_write_en_0 ? _GEN_259 : buffer_9_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_324 = io_write_en_0 ? _GEN_260 : buffer_10_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_325 = io_write_en_0 ? _GEN_261 : buffer_11_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_326 = io_write_en_0 ? _GEN_262 : buffer_12_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_327 = io_write_en_0 ? _GEN_263 : buffer_13_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_328 = io_write_en_0 ? _GEN_264 : buffer_14_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_329 = io_write_en_0 ? _GEN_265 : buffer_15_data; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_330 = io_write_en_0 ? _GEN_266 : buffer_0_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_331 = io_write_en_0 ? _GEN_267 : buffer_1_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_332 = io_write_en_0 ? _GEN_268 : buffer_2_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_333 = io_write_en_0 ? _GEN_269 : buffer_3_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_334 = io_write_en_0 ? _GEN_270 : buffer_4_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_335 = io_write_en_0 ? _GEN_271 : buffer_5_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_336 = io_write_en_0 ? _GEN_272 : buffer_6_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_337 = io_write_en_0 ? _GEN_273 : buffer_7_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_338 = io_write_en_0 ? _GEN_274 : buffer_8_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_339 = io_write_en_0 ? _GEN_275 : buffer_9_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_340 = io_write_en_0 ? _GEN_276 : buffer_10_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_341 = io_write_en_0 ? _GEN_277 : buffer_11_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_342 = io_write_en_0 ? _GEN_278 : buffer_12_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_343 = io_write_en_0 ? _GEN_279 : buffer_13_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_344 = io_write_en_0 ? _GEN_280 : buffer_14_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [31:0] _GEN_345 = io_write_en_0 ? _GEN_281 : buffer_15_addr; // @[InstBuffer.scala 124:53 41:23]
  wire [3:0] _T_21 = enq_ptr + 4'h1; // @[InstBuffer.scala 124:70]
  wire [3:0] _enq_ptr_T_1 = enq_ptr + 4'h2; // @[InstBuffer.scala 129:24]
  assign io_master_is_in_delayslot_o = master_is_in_delayslot; // @[InstBuffer.scala 55:31]
  assign io_read_0_tlb_invalid = delayslot_enable ? delayslot_line_tlb_invalid : _io_read_0_T_1_tlb_invalid; // @[Mux.scala 101:16]
  assign io_read_0_data = delayslot_enable ? delayslot_line_data : _io_read_0_T_1_data; // @[Mux.scala 101:16]
  assign io_read_0_addr = delayslot_enable ? delayslot_line_addr : _io_read_0_T_1_addr; // @[Mux.scala 101:16]
  assign io_read_1_tlb_invalid = delayslot_enable ? 1'h0 : _io_read_1_T_3_tlb_invalid; // @[Mux.scala 101:16]
  assign io_read_1_data = delayslot_enable ? 32'h0 : _io_read_1_T_3_data; // @[Mux.scala 101:16]
  assign io_read_1_addr = delayslot_enable ? 32'h0 : _io_read_1_T_3_addr; // @[Mux.scala 101:16]
  assign io_empty = _GEN_477 == 5'h0; // @[InstBuffer.scala 51:28]
  assign io_almost_empty = _GEN_477 == 5'h1; // @[InstBuffer.scala 52:28]
  assign io_full = _GEN_477 >= 5'he; // @[InstBuffer.scala 50:28]
  always @(posedge clock) begin
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_0_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h0 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_0_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_0_tlb_invalid <= _GEN_298;
      end
    end else begin
      buffer_0_tlb_invalid <= _GEN_298;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_0_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h0 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_0_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_0_data <= _GEN_314;
      end
    end else begin
      buffer_0_data <= _GEN_314;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_0_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h0 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_0_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_0_addr <= _GEN_330;
      end
    end else begin
      buffer_0_addr <= _GEN_330;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_1_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h1 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_1_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_1_tlb_invalid <= _GEN_299;
      end
    end else begin
      buffer_1_tlb_invalid <= _GEN_299;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_1_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h1 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_1_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_1_data <= _GEN_315;
      end
    end else begin
      buffer_1_data <= _GEN_315;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_1_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h1 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_1_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_1_addr <= _GEN_331;
      end
    end else begin
      buffer_1_addr <= _GEN_331;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_2_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h2 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_2_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_2_tlb_invalid <= _GEN_300;
      end
    end else begin
      buffer_2_tlb_invalid <= _GEN_300;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_2_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h2 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_2_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_2_data <= _GEN_316;
      end
    end else begin
      buffer_2_data <= _GEN_316;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_2_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h2 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_2_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_2_addr <= _GEN_332;
      end
    end else begin
      buffer_2_addr <= _GEN_332;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_3_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h3 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_3_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_3_tlb_invalid <= _GEN_301;
      end
    end else begin
      buffer_3_tlb_invalid <= _GEN_301;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_3_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h3 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_3_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_3_data <= _GEN_317;
      end
    end else begin
      buffer_3_data <= _GEN_317;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_3_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h3 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_3_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_3_addr <= _GEN_333;
      end
    end else begin
      buffer_3_addr <= _GEN_333;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_4_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h4 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_4_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_4_tlb_invalid <= _GEN_302;
      end
    end else begin
      buffer_4_tlb_invalid <= _GEN_302;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_4_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h4 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_4_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_4_data <= _GEN_318;
      end
    end else begin
      buffer_4_data <= _GEN_318;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_4_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h4 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_4_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_4_addr <= _GEN_334;
      end
    end else begin
      buffer_4_addr <= _GEN_334;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_5_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h5 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_5_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_5_tlb_invalid <= _GEN_303;
      end
    end else begin
      buffer_5_tlb_invalid <= _GEN_303;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_5_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h5 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_5_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_5_data <= _GEN_319;
      end
    end else begin
      buffer_5_data <= _GEN_319;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_5_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h5 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_5_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_5_addr <= _GEN_335;
      end
    end else begin
      buffer_5_addr <= _GEN_335;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_6_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h6 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_6_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_6_tlb_invalid <= _GEN_304;
      end
    end else begin
      buffer_6_tlb_invalid <= _GEN_304;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_6_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h6 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_6_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_6_data <= _GEN_320;
      end
    end else begin
      buffer_6_data <= _GEN_320;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_6_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h6 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_6_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_6_addr <= _GEN_336;
      end
    end else begin
      buffer_6_addr <= _GEN_336;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_7_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h7 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_7_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_7_tlb_invalid <= _GEN_305;
      end
    end else begin
      buffer_7_tlb_invalid <= _GEN_305;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_7_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h7 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_7_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_7_data <= _GEN_321;
      end
    end else begin
      buffer_7_data <= _GEN_321;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_7_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h7 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_7_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_7_addr <= _GEN_337;
      end
    end else begin
      buffer_7_addr <= _GEN_337;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_8_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h8 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_8_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_8_tlb_invalid <= _GEN_306;
      end
    end else begin
      buffer_8_tlb_invalid <= _GEN_306;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_8_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h8 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_8_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_8_data <= _GEN_322;
      end
    end else begin
      buffer_8_data <= _GEN_322;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_8_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h8 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_8_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_8_addr <= _GEN_338;
      end
    end else begin
      buffer_8_addr <= _GEN_338;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_9_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h9 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_9_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_9_tlb_invalid <= _GEN_307;
      end
    end else begin
      buffer_9_tlb_invalid <= _GEN_307;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_9_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h9 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_9_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_9_data <= _GEN_323;
      end
    end else begin
      buffer_9_data <= _GEN_323;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_9_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'h9 == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_9_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_9_addr <= _GEN_339;
      end
    end else begin
      buffer_9_addr <= _GEN_339;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_10_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'ha == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_10_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_10_tlb_invalid <= _GEN_308;
      end
    end else begin
      buffer_10_tlb_invalid <= _GEN_308;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_10_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'ha == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_10_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_10_data <= _GEN_324;
      end
    end else begin
      buffer_10_data <= _GEN_324;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_10_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'ha == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_10_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_10_addr <= _GEN_340;
      end
    end else begin
      buffer_10_addr <= _GEN_340;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_11_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hb == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_11_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_11_tlb_invalid <= _GEN_309;
      end
    end else begin
      buffer_11_tlb_invalid <= _GEN_309;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_11_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hb == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_11_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_11_data <= _GEN_325;
      end
    end else begin
      buffer_11_data <= _GEN_325;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_11_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hb == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_11_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_11_addr <= _GEN_341;
      end
    end else begin
      buffer_11_addr <= _GEN_341;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_12_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hc == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_12_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_12_tlb_invalid <= _GEN_310;
      end
    end else begin
      buffer_12_tlb_invalid <= _GEN_310;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_12_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hc == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_12_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_12_data <= _GEN_326;
      end
    end else begin
      buffer_12_data <= _GEN_326;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_12_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hc == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_12_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_12_addr <= _GEN_342;
      end
    end else begin
      buffer_12_addr <= _GEN_342;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_13_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hd == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_13_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_13_tlb_invalid <= _GEN_311;
      end
    end else begin
      buffer_13_tlb_invalid <= _GEN_311;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_13_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hd == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_13_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_13_data <= _GEN_327;
      end
    end else begin
      buffer_13_data <= _GEN_327;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_13_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hd == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_13_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_13_addr <= _GEN_343;
      end
    end else begin
      buffer_13_addr <= _GEN_343;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_14_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'he == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_14_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_14_tlb_invalid <= _GEN_312;
      end
    end else begin
      buffer_14_tlb_invalid <= _GEN_312;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_14_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'he == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_14_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_14_data <= _GEN_328;
      end
    end else begin
      buffer_14_data <= _GEN_328;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_14_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'he == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_14_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_14_addr <= _GEN_344;
      end
    end else begin
      buffer_14_addr <= _GEN_344;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_15_tlb_invalid <= 1'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hf == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_15_tlb_invalid <= io_write_1_tlb_invalid; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_15_tlb_invalid <= _GEN_313;
      end
    end else begin
      buffer_15_tlb_invalid <= _GEN_313;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_15_data <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hf == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_15_data <= io_write_1_data; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_15_data <= _GEN_329;
      end
    end else begin
      buffer_15_data <= _GEN_329;
    end
    if (reset) begin // @[InstBuffer.scala 41:23]
      buffer_15_addr <= 32'h0; // @[InstBuffer.scala 41:23]
    end else if (io_write_en_1) begin // @[InstBuffer.scala 124:53]
      if (4'hf == _T_21) begin // @[InstBuffer.scala 124:77]
        buffer_15_addr <= io_write_1_addr; // @[InstBuffer.scala 124:77]
      end else begin
        buffer_15_addr <= _GEN_345;
      end
    end else begin
      buffer_15_addr <= _GEN_345;
    end
    if (reset) begin // @[InstBuffer.scala 44:24]
      enq_ptr <= 4'h0; // @[InstBuffer.scala 44:24]
    end else if (io_fifo_rst) begin // @[InstBuffer.scala 126:21]
      enq_ptr <= 4'h0; // @[InstBuffer.scala 127:13]
    end else if (io_write_en_0 & io_write_en_1) begin // @[InstBuffer.scala 128:48]
      enq_ptr <= _enq_ptr_T_1; // @[InstBuffer.scala 129:13]
    end else if (io_write_en_0) begin // @[InstBuffer.scala 130:30]
      enq_ptr <= _T_21; // @[InstBuffer.scala 131:13]
    end
    if (reset) begin // @[InstBuffer.scala 45:24]
      deq_ptr <= 4'h0; // @[InstBuffer.scala 45:24]
    end else if (io_fifo_rst) begin // @[InstBuffer.scala 113:21]
      deq_ptr <= 4'h0; // @[InstBuffer.scala 114:13]
    end else if (!(io_empty | delayslot_enable)) begin // @[InstBuffer.scala 115:44]
      if (io_read_en_0 & io_read_en_1) begin // @[InstBuffer.scala 117:46]
        deq_ptr <= _deq_ptr_T_1; // @[InstBuffer.scala 118:13]
      end else begin
        deq_ptr <= _GEN_214;
      end
    end
    if (reset) begin // @[InstBuffer.scala 54:39]
      master_is_in_delayslot <= 1'h0; // @[InstBuffer.scala 54:39]
    end else if (io_flush_delay_slot) begin // @[Mux.scala 101:16]
      master_is_in_delayslot <= 1'h0;
    end else if (!(_master_is_in_delayslot_T)) begin // @[Mux.scala 101:16]
      master_is_in_delayslot <= _master_is_in_delayslot_T_2;
    end
    if (reset) begin // @[InstBuffer.scala 65:33]
      delayslot_stall <= 1'h0; // @[InstBuffer.scala 65:33]
    end else begin
      delayslot_stall <= _GEN_1;
    end
    if (reset) begin // @[InstBuffer.scala 66:33]
      delayslot_enable <= 1'h0; // @[InstBuffer.scala 66:33]
    end else if (io_fifo_rst & _T_1 & io_delay_sel_rst) begin // @[InstBuffer.scala 76:65]
      delayslot_enable <= _GEN_135;
    end else if (~delayslot_stall & io_read_en_0) begin // @[InstBuffer.scala 91:49]
      delayslot_enable <= 1'h0; // @[InstBuffer.scala 92:22]
    end
    if (reset) begin // @[InstBuffer.scala 67:33]
      delayslot_line_tlb_invalid <= 1'h0; // @[InstBuffer.scala 67:33]
    end else if (io_fifo_rst & _T_1 & io_delay_sel_rst) begin // @[InstBuffer.scala 76:65]
      if (io_E_delay_rst) begin // @[InstBuffer.scala 77:26]
        if (_T_7) begin // @[InstBuffer.scala 79:30]
          delayslot_line_tlb_invalid <= io_write_0_tlb_invalid;
        end else begin
          delayslot_line_tlb_invalid <= _GEN_63;
        end
      end else begin
        delayslot_line_tlb_invalid <= _GEN_132;
      end
    end else if (~delayslot_stall & io_read_en_0) begin // @[InstBuffer.scala 91:49]
      delayslot_line_tlb_invalid <= 1'h0; // @[InstBuffer.scala 93:22]
    end
    if (reset) begin // @[InstBuffer.scala 67:33]
      delayslot_line_data <= 32'h0; // @[InstBuffer.scala 67:33]
    end else if (io_fifo_rst & _T_1 & io_delay_sel_rst) begin // @[InstBuffer.scala 76:65]
      if (io_E_delay_rst) begin // @[InstBuffer.scala 77:26]
        if (_T_7) begin // @[InstBuffer.scala 79:30]
          delayslot_line_data <= io_write_0_data;
        end else begin
          delayslot_line_data <= _GEN_64;
        end
      end else if (io_D_delay_rst) begin // @[InstBuffer.scala 80:32]
        delayslot_line_data <= _delayslot_line_T_7_data; // @[InstBuffer.scala 82:22]
      end else begin
        delayslot_line_data <= 32'h0; // @[InstBuffer.scala 89:24]
      end
    end else if (~delayslot_stall & io_read_en_0) begin // @[InstBuffer.scala 91:49]
      delayslot_line_data <= 32'h0; // @[InstBuffer.scala 93:22]
    end
    if (reset) begin // @[InstBuffer.scala 67:33]
      delayslot_line_addr <= 32'h0; // @[InstBuffer.scala 67:33]
    end else if (io_fifo_rst & _T_1 & io_delay_sel_rst) begin // @[InstBuffer.scala 76:65]
      if (io_E_delay_rst) begin // @[InstBuffer.scala 77:26]
        if (_T_7) begin // @[InstBuffer.scala 79:30]
          delayslot_line_addr <= io_write_0_addr;
        end else begin
          delayslot_line_addr <= _GEN_65;
        end
      end else if (io_D_delay_rst) begin // @[InstBuffer.scala 80:32]
        delayslot_line_addr <= _delayslot_line_T_7_addr; // @[InstBuffer.scala 82:22]
      end else begin
        delayslot_line_addr <= 32'h0; // @[InstBuffer.scala 89:24]
      end
    end else if (~delayslot_stall & io_read_en_0) begin // @[InstBuffer.scala 91:49]
      delayslot_line_addr <= 32'h0; // @[InstBuffer.scala 93:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buffer_0_tlb_invalid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  buffer_0_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_0_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_1_tlb_invalid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_1_data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_1_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_2_tlb_invalid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_2_data = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_2_addr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_3_tlb_invalid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_3_data = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_3_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_4_tlb_invalid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_4_data = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_4_addr = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_5_tlb_invalid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_5_data = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_5_addr = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_6_tlb_invalid = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  buffer_6_data = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_6_addr = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_7_tlb_invalid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  buffer_7_data = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  buffer_7_addr = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  buffer_8_tlb_invalid = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_8_data = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  buffer_8_addr = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_9_tlb_invalid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_9_data = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  buffer_9_addr = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  buffer_10_tlb_invalid = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_10_data = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_10_addr = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_11_tlb_invalid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  buffer_11_data = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  buffer_11_addr = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  buffer_12_tlb_invalid = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_12_data = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_12_addr = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  buffer_13_tlb_invalid = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_13_data = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  buffer_13_addr = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  buffer_14_tlb_invalid = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_14_data = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  buffer_14_addr = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_15_tlb_invalid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_15_data = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  buffer_15_addr = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  enq_ptr = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  deq_ptr = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  master_is_in_delayslot = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  delayslot_stall = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  delayslot_enable = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  delayslot_line_tlb_invalid = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  delayslot_line_data = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  delayslot_line_addr = _RAND_55[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Issue(
  input        io_allow_to_go,
  input        io_instBuffer_empty,
  input        io_instBuffer_almost_empty,
  input  [3:0] io_decodeInst_0_fusel,
  input        io_decodeInst_0_reg_wen,
  input  [4:0] io_decodeInst_0_reg_waddr,
  input        io_decodeInst_0_dual_issue,
  input        io_decodeInst_1_reg1_ren,
  input  [4:0] io_decodeInst_1_reg1_raddr,
  input        io_decodeInst_1_reg2_ren,
  input  [4:0] io_decodeInst_1_reg2_raddr,
  input  [3:0] io_decodeInst_1_fusel,
  input        io_decodeInst_1_dual_issue,
  input        io_execute_0_mem_ren,
  input  [4:0] io_execute_0_reg_waddr,
  input        io_execute_1_mem_ren,
  input  [4:0] io_execute_1_reg_waddr,
  output       io_inst1_is_in_delayslot,
  output       io_inst1_allow_to_go
);
  wire  instBuffer_invalid = io_instBuffer_empty | io_instBuffer_almost_empty; // @[Issue.scala 30:48]
  wire  mem_conflict = io_decodeInst_0_fusel == 4'h4 & io_decodeInst_1_fusel == 4'h4; // @[Issue.scala 33:48]
  wire  mul_conflict = io_decodeInst_0_fusel == 4'hb & io_decodeInst_1_fusel == 4'hb; // @[Issue.scala 34:48]
  wire  div_conflict = io_decodeInst_0_fusel == 4'hc & io_decodeInst_1_fusel == 4'hc; // @[Issue.scala 35:48]
  wire  struct_conflict = mem_conflict | mul_conflict | div_conflict; // @[Issue.scala 36:54]
  wire  _load_stall_T_3 = io_decodeInst_1_reg2_ren & io_decodeInst_1_reg2_raddr == io_execute_0_reg_waddr; // @[Issue.scala 41:22]
  wire  _load_stall_T_5 = io_execute_0_mem_ren & (io_decodeInst_1_reg1_ren & io_decodeInst_1_reg1_raddr ==
    io_execute_0_reg_waddr | _load_stall_T_3); // @[Issue.scala 40:27]
  wire  _load_stall_T_9 = io_decodeInst_1_reg2_ren & io_decodeInst_1_reg2_raddr == io_execute_1_reg_waddr; // @[Issue.scala 43:24]
  wire  _load_stall_T_11 = io_execute_1_mem_ren & (io_decodeInst_1_reg1_ren & io_decodeInst_1_reg1_raddr ==
    io_execute_1_reg_waddr | _load_stall_T_9); // @[Issue.scala 42:29]
  wire  load_stall = _load_stall_T_5 | _load_stall_T_11; // @[Issue.scala 41:71]
  wire  raw_reg = io_decodeInst_0_reg_wen & (io_decodeInst_0_reg_waddr == io_decodeInst_1_reg1_raddr &
    io_decodeInst_1_reg1_ren | io_decodeInst_0_reg_waddr == io_decodeInst_1_reg2_raddr & io_decodeInst_1_reg2_ren); // @[Issue.scala 45:19]
  wire  _raw_hilo_T_13 = 4'hc == io_decodeInst_1_fusel | 4'hb == io_decodeInst_1_fusel | 4'h9 == io_decodeInst_1_fusel
     | 4'ha == io_decodeInst_1_fusel; // @[Issue.scala 47:59]
  wire  raw_hilo = (4'hc == io_decodeInst_0_fusel | 4'hb == io_decodeInst_0_fusel | 4'h9 == io_decodeInst_0_fusel) &
    _raw_hilo_T_13; // @[Issue.scala 46:75]
  wire  raw_cp0 = io_decodeInst_0_fusel == 4'h2 & io_decodeInst_1_fusel == 4'h3; // @[Issue.scala 49:29]
  wire  data_conflict = raw_reg | raw_hilo | raw_cp0 | load_stall; // @[Issue.scala 50:54]
  wire  _io_inst1_allow_to_go_T = ~instBuffer_invalid; // @[Issue.scala 56:5]
  wire  _io_inst1_allow_to_go_T_1 = io_allow_to_go & _io_inst1_allow_to_go_T; // @[Issue.scala 55:42]
  wire  _io_inst1_allow_to_go_T_2 = _io_inst1_allow_to_go_T_1 & io_decodeInst_0_dual_issue; // @[Issue.scala 56:25]
  wire  _io_inst1_allow_to_go_T_3 = _io_inst1_allow_to_go_T_2 & io_decodeInst_1_dual_issue; // @[Issue.scala 57:22]
  wire  _io_inst1_allow_to_go_T_4 = ~struct_conflict; // @[Issue.scala 59:5]
  wire  _io_inst1_allow_to_go_T_5 = _io_inst1_allow_to_go_T_3 & _io_inst1_allow_to_go_T_4; // @[Issue.scala 58:22]
  wire  _io_inst1_allow_to_go_T_6 = ~data_conflict; // @[Issue.scala 60:5]
  wire  _io_inst1_allow_to_go_T_7 = _io_inst1_allow_to_go_T_5 & _io_inst1_allow_to_go_T_6; // @[Issue.scala 59:22]
  wire  _io_inst1_allow_to_go_T_14 = ~(4'h5 == io_decodeInst_1_fusel | 4'h8 == io_decodeInst_1_fusel | 4'h7 ==
    io_decodeInst_1_fusel); // @[Issue.scala 61:5]
  assign io_inst1_is_in_delayslot = io_decodeInst_0_fusel == 4'h5 & io_inst1_allow_to_go; // @[Issue.scala 53:53]
  assign io_inst1_allow_to_go = _io_inst1_allow_to_go_T_7 & _io_inst1_allow_to_go_T_14; // @[Issue.scala 60:20]
endmodule
module Decoder(
  input  [31:0] io_in_inst,
  output        io_out_inst_valid,
  output        io_out_reg1_ren,
  output [4:0]  io_out_reg1_raddr,
  output        io_out_reg2_ren,
  output [4:0]  io_out_reg2_raddr,
  output [3:0]  io_out_fusel,
  output [6:0]  io_out_op,
  output        io_out_reg_wen,
  output [4:0]  io_out_reg_waddr,
  output [31:0] io_out_imm32,
  output [7:0]  io_out_cp0_addr,
  output        io_out_dual_issue,
  output [31:0] io_out_inst
);
  wire  _signals_T_1 = 32'h0 == io_in_inst; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_2 = io_in_inst & 32'hfc0007ff; // @[Lookup.scala 31:38]
  wire  _signals_T_3 = 32'h25 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_5 = 32'h24 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_7 = 32'h26 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_9 = 32'h27 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_11 = 32'h4 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_13 = 32'h6 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_15 = 32'h7 == _signals_T_2; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_16 = io_in_inst & 32'hffe0003f; // @[Lookup.scala 31:38]
  wire  _signals_T_17 = 32'h0 == _signals_T_16; // @[Lookup.scala 31:38]
  wire  _signals_T_19 = 32'h2 == _signals_T_16; // @[Lookup.scala 31:38]
  wire  _signals_T_21 = 32'h3 == _signals_T_16; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_22 = io_in_inst & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _signals_T_23 = 32'h34000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_25 = 32'h30000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_27 = 32'h38000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_28 = io_in_inst & 32'hffe00000; // @[Lookup.scala 31:38]
  wire  _signals_T_29 = 32'h3c000000 == _signals_T_28; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_30 = io_in_inst & 32'hffff07ff; // @[Lookup.scala 31:38]
  wire  _signals_T_31 = 32'h10 == _signals_T_30; // @[Lookup.scala 31:38]
  wire  _signals_T_33 = 32'h12 == _signals_T_30; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_34 = io_in_inst & 32'hfc1fffff; // @[Lookup.scala 31:38]
  wire  _signals_T_35 = 32'h11 == _signals_T_34; // @[Lookup.scala 31:38]
  wire  _signals_T_37 = 32'h13 == _signals_T_34; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_38 = io_in_inst & 32'hffe007f8; // @[Lookup.scala 31:38]
  wire  _signals_T_39 = 32'h40000000 == _signals_T_38; // @[Lookup.scala 31:38]
  wire  _signals_T_41 = 32'h40800000 == _signals_T_38; // @[Lookup.scala 31:38]
  wire  _signals_T_43 = 32'h2a == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_45 = 32'h2b == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_47 = 32'h28000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_49 = 32'h2c000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_51 = 32'h20 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_53 = 32'h21 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_55 = 32'h22 == _signals_T_2; // @[Lookup.scala 31:38]
  wire  _signals_T_57 = 32'h23 == _signals_T_2; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_58 = io_in_inst & 32'hfc00ffff; // @[Lookup.scala 31:38]
  wire  _signals_T_59 = 32'h18 == _signals_T_58; // @[Lookup.scala 31:38]
  wire  _signals_T_61 = 32'h19 == _signals_T_58; // @[Lookup.scala 31:38]
  wire  _signals_T_63 = 32'h1a == _signals_T_58; // @[Lookup.scala 31:38]
  wire  _signals_T_65 = 32'h1b == _signals_T_58; // @[Lookup.scala 31:38]
  wire  _signals_T_67 = 32'h20000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_69 = 32'h24000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_71 = 32'h8000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_73 = 32'hc000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_74 = io_in_inst & 32'hfc1ff83f; // @[Lookup.scala 31:38]
  wire  _signals_T_75 = 32'h8 == _signals_T_74; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_76 = io_in_inst & 32'hfc1f003f; // @[Lookup.scala 31:38]
  wire  _signals_T_77 = 32'h9 == _signals_T_76; // @[Lookup.scala 31:38]
  wire  _signals_T_79 = 32'h10000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_81 = 32'h14000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_82 = io_in_inst & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _signals_T_83 = 32'h1c000000 == _signals_T_82; // @[Lookup.scala 31:38]
  wire  _signals_T_85 = 32'h18000000 == _signals_T_82; // @[Lookup.scala 31:38]
  wire  _signals_T_87 = 32'h4010000 == _signals_T_82; // @[Lookup.scala 31:38]
  wire  _signals_T_89 = 32'h4110000 == _signals_T_82; // @[Lookup.scala 31:38]
  wire  _signals_T_91 = 32'h4000000 == _signals_T_82; // @[Lookup.scala 31:38]
  wire  _signals_T_93 = 32'h4100000 == _signals_T_82; // @[Lookup.scala 31:38]
  wire  _signals_T_95 = 32'h42000008 == io_in_inst; // @[Lookup.scala 31:38]
  wire  _signals_T_97 = 32'h42000001 == io_in_inst; // @[Lookup.scala 31:38]
  wire  _signals_T_99 = 32'h42000002 == io_in_inst; // @[Lookup.scala 31:38]
  wire  _signals_T_101 = 32'h42000006 == io_in_inst; // @[Lookup.scala 31:38]
  wire [31:0] _signals_T_102 = io_in_inst & 32'hfc00003f; // @[Lookup.scala 31:38]
  wire  _signals_T_103 = 32'hc == _signals_T_102; // @[Lookup.scala 31:38]
  wire  _signals_T_105 = 32'hd == _signals_T_102; // @[Lookup.scala 31:38]
  wire  _signals_T_107 = 32'h42000018 == io_in_inst; // @[Lookup.scala 31:38]
  wire  _signals_T_109 = 32'h80000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_111 = 32'h90000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_113 = 32'h84000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_115 = 32'h94000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_117 = 32'h8c000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_119 = 32'ha0000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_121 = 32'ha4000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_123 = 32'hac000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_125 = 32'h88000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_127 = 32'h98000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_129 = 32'ha8000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_131 = 32'hb8000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_133 = 32'hbc000000 == _signals_T_22; // @[Lookup.scala 31:38]
  wire  _signals_T_134 = _signals_T_133 ? 1'h0 : 1'h1; // @[Lookup.scala 34:39]
  wire  _signals_T_135 = _signals_T_131 ? 1'h0 : _signals_T_134; // @[Lookup.scala 34:39]
  wire  _signals_T_136 = _signals_T_129 ? 1'h0 : _signals_T_135; // @[Lookup.scala 34:39]
  wire  _signals_T_137 = _signals_T_127 ? 1'h0 : _signals_T_136; // @[Lookup.scala 34:39]
  wire  _signals_T_138 = _signals_T_125 ? 1'h0 : _signals_T_137; // @[Lookup.scala 34:39]
  wire  _signals_T_139 = _signals_T_123 ? 1'h0 : _signals_T_138; // @[Lookup.scala 34:39]
  wire  _signals_T_140 = _signals_T_121 ? 1'h0 : _signals_T_139; // @[Lookup.scala 34:39]
  wire  _signals_T_141 = _signals_T_119 ? 1'h0 : _signals_T_140; // @[Lookup.scala 34:39]
  wire  _signals_T_142 = _signals_T_117 ? 1'h0 : _signals_T_141; // @[Lookup.scala 34:39]
  wire  _signals_T_143 = _signals_T_115 ? 1'h0 : _signals_T_142; // @[Lookup.scala 34:39]
  wire  _signals_T_144 = _signals_T_113 ? 1'h0 : _signals_T_143; // @[Lookup.scala 34:39]
  wire  _signals_T_145 = _signals_T_111 ? 1'h0 : _signals_T_144; // @[Lookup.scala 34:39]
  wire  _signals_T_146 = _signals_T_109 ? 1'h0 : _signals_T_145; // @[Lookup.scala 34:39]
  wire  _signals_T_147 = _signals_T_107 ? 1'h0 : _signals_T_146; // @[Lookup.scala 34:39]
  wire  _signals_T_148 = _signals_T_105 ? 1'h0 : _signals_T_147; // @[Lookup.scala 34:39]
  wire  _signals_T_149 = _signals_T_103 ? 1'h0 : _signals_T_148; // @[Lookup.scala 34:39]
  wire  _signals_T_150 = _signals_T_101 ? 1'h0 : _signals_T_149; // @[Lookup.scala 34:39]
  wire  _signals_T_151 = _signals_T_99 ? 1'h0 : _signals_T_150; // @[Lookup.scala 34:39]
  wire  _signals_T_152 = _signals_T_97 ? 1'h0 : _signals_T_151; // @[Lookup.scala 34:39]
  wire  _signals_T_153 = _signals_T_95 ? 1'h0 : _signals_T_152; // @[Lookup.scala 34:39]
  wire  _signals_T_154 = _signals_T_93 ? 1'h0 : _signals_T_153; // @[Lookup.scala 34:39]
  wire  _signals_T_155 = _signals_T_91 ? 1'h0 : _signals_T_154; // @[Lookup.scala 34:39]
  wire  _signals_T_156 = _signals_T_89 ? 1'h0 : _signals_T_155; // @[Lookup.scala 34:39]
  wire  _signals_T_157 = _signals_T_87 ? 1'h0 : _signals_T_156; // @[Lookup.scala 34:39]
  wire  _signals_T_158 = _signals_T_85 ? 1'h0 : _signals_T_157; // @[Lookup.scala 34:39]
  wire  _signals_T_159 = _signals_T_83 ? 1'h0 : _signals_T_158; // @[Lookup.scala 34:39]
  wire  _signals_T_160 = _signals_T_81 ? 1'h0 : _signals_T_159; // @[Lookup.scala 34:39]
  wire  _signals_T_161 = _signals_T_79 ? 1'h0 : _signals_T_160; // @[Lookup.scala 34:39]
  wire  _signals_T_162 = _signals_T_77 ? 1'h0 : _signals_T_161; // @[Lookup.scala 34:39]
  wire  _signals_T_163 = _signals_T_75 ? 1'h0 : _signals_T_162; // @[Lookup.scala 34:39]
  wire  _signals_T_164 = _signals_T_73 ? 1'h0 : _signals_T_163; // @[Lookup.scala 34:39]
  wire  _signals_T_165 = _signals_T_71 ? 1'h0 : _signals_T_164; // @[Lookup.scala 34:39]
  wire  _signals_T_166 = _signals_T_69 ? 1'h0 : _signals_T_165; // @[Lookup.scala 34:39]
  wire  _signals_T_167 = _signals_T_67 ? 1'h0 : _signals_T_166; // @[Lookup.scala 34:39]
  wire  _signals_T_168 = _signals_T_65 ? 1'h0 : _signals_T_167; // @[Lookup.scala 34:39]
  wire  _signals_T_169 = _signals_T_63 ? 1'h0 : _signals_T_168; // @[Lookup.scala 34:39]
  wire  _signals_T_170 = _signals_T_61 ? 1'h0 : _signals_T_169; // @[Lookup.scala 34:39]
  wire  _signals_T_171 = _signals_T_59 ? 1'h0 : _signals_T_170; // @[Lookup.scala 34:39]
  wire  _signals_T_172 = _signals_T_57 ? 1'h0 : _signals_T_171; // @[Lookup.scala 34:39]
  wire  _signals_T_173 = _signals_T_55 ? 1'h0 : _signals_T_172; // @[Lookup.scala 34:39]
  wire  _signals_T_174 = _signals_T_53 ? 1'h0 : _signals_T_173; // @[Lookup.scala 34:39]
  wire  _signals_T_175 = _signals_T_51 ? 1'h0 : _signals_T_174; // @[Lookup.scala 34:39]
  wire  _signals_T_176 = _signals_T_49 ? 1'h0 : _signals_T_175; // @[Lookup.scala 34:39]
  wire  _signals_T_177 = _signals_T_47 ? 1'h0 : _signals_T_176; // @[Lookup.scala 34:39]
  wire  _signals_T_178 = _signals_T_45 ? 1'h0 : _signals_T_177; // @[Lookup.scala 34:39]
  wire  _signals_T_179 = _signals_T_43 ? 1'h0 : _signals_T_178; // @[Lookup.scala 34:39]
  wire  _signals_T_180 = _signals_T_41 ? 1'h0 : _signals_T_179; // @[Lookup.scala 34:39]
  wire  _signals_T_181 = _signals_T_39 ? 1'h0 : _signals_T_180; // @[Lookup.scala 34:39]
  wire  _signals_T_182 = _signals_T_37 ? 1'h0 : _signals_T_181; // @[Lookup.scala 34:39]
  wire  _signals_T_183 = _signals_T_35 ? 1'h0 : _signals_T_182; // @[Lookup.scala 34:39]
  wire  _signals_T_184 = _signals_T_33 ? 1'h0 : _signals_T_183; // @[Lookup.scala 34:39]
  wire  _signals_T_185 = _signals_T_31 ? 1'h0 : _signals_T_184; // @[Lookup.scala 34:39]
  wire  _signals_T_186 = _signals_T_29 ? 1'h0 : _signals_T_185; // @[Lookup.scala 34:39]
  wire  _signals_T_187 = _signals_T_27 ? 1'h0 : _signals_T_186; // @[Lookup.scala 34:39]
  wire  _signals_T_188 = _signals_T_25 ? 1'h0 : _signals_T_187; // @[Lookup.scala 34:39]
  wire  _signals_T_189 = _signals_T_23 ? 1'h0 : _signals_T_188; // @[Lookup.scala 34:39]
  wire  _signals_T_190 = _signals_T_21 ? 1'h0 : _signals_T_189; // @[Lookup.scala 34:39]
  wire  _signals_T_191 = _signals_T_19 ? 1'h0 : _signals_T_190; // @[Lookup.scala 34:39]
  wire  _signals_T_192 = _signals_T_17 ? 1'h0 : _signals_T_191; // @[Lookup.scala 34:39]
  wire  _signals_T_193 = _signals_T_15 ? 1'h0 : _signals_T_192; // @[Lookup.scala 34:39]
  wire  _signals_T_194 = _signals_T_13 ? 1'h0 : _signals_T_193; // @[Lookup.scala 34:39]
  wire  _signals_T_195 = _signals_T_11 ? 1'h0 : _signals_T_194; // @[Lookup.scala 34:39]
  wire  _signals_T_196 = _signals_T_9 ? 1'h0 : _signals_T_195; // @[Lookup.scala 34:39]
  wire  _signals_T_197 = _signals_T_7 ? 1'h0 : _signals_T_196; // @[Lookup.scala 34:39]
  wire  _signals_T_198 = _signals_T_5 ? 1'h0 : _signals_T_197; // @[Lookup.scala 34:39]
  wire  _signals_T_199 = _signals_T_3 ? 1'h0 : _signals_T_198; // @[Lookup.scala 34:39]
  wire  _signals_T_213 = _signals_T_107 ? 1'h0 : _signals_T_109 | (_signals_T_111 | (_signals_T_113 | (_signals_T_115 |
    (_signals_T_117 | (_signals_T_119 | (_signals_T_121 | (_signals_T_123 | (_signals_T_125 | (_signals_T_127 | (
    _signals_T_129 | (_signals_T_131 | _signals_T_133))))))))))); // @[Lookup.scala 34:39]
  wire  _signals_T_214 = _signals_T_105 ? 1'h0 : _signals_T_213; // @[Lookup.scala 34:39]
  wire  _signals_T_215 = _signals_T_103 ? 1'h0 : _signals_T_214; // @[Lookup.scala 34:39]
  wire  _signals_T_216 = _signals_T_101 ? 1'h0 : _signals_T_215; // @[Lookup.scala 34:39]
  wire  _signals_T_217 = _signals_T_99 ? 1'h0 : _signals_T_216; // @[Lookup.scala 34:39]
  wire  _signals_T_218 = _signals_T_97 ? 1'h0 : _signals_T_217; // @[Lookup.scala 34:39]
  wire  _signals_T_219 = _signals_T_95 ? 1'h0 : _signals_T_218; // @[Lookup.scala 34:39]
  wire  _signals_T_230 = _signals_T_73 ? 1'h0 : _signals_T_75 | (_signals_T_77 | (_signals_T_79 | (_signals_T_81 | (
    _signals_T_83 | (_signals_T_85 | (_signals_T_87 | (_signals_T_89 | (_signals_T_91 | (_signals_T_93 | _signals_T_219)
    )))))))); // @[Lookup.scala 34:39]
  wire  _signals_T_231 = _signals_T_71 ? 1'h0 : _signals_T_230; // @[Lookup.scala 34:39]
  wire  _signals_T_246 = _signals_T_41 ? 1'h0 : _signals_T_43 | (_signals_T_45 | (_signals_T_47 | (_signals_T_49 | (
    _signals_T_51 | (_signals_T_53 | (_signals_T_55 | (_signals_T_57 | (_signals_T_59 | (_signals_T_61 | (_signals_T_63
     | (_signals_T_65 | (_signals_T_67 | (_signals_T_69 | _signals_T_231))))))))))))); // @[Lookup.scala 34:39]
  wire  _signals_T_247 = _signals_T_39 ? 1'h0 : _signals_T_246; // @[Lookup.scala 34:39]
  wire  _signals_T_250 = _signals_T_33 ? 1'h0 : _signals_T_35 | (_signals_T_37 | _signals_T_247); // @[Lookup.scala 34:39]
  wire  _signals_T_251 = _signals_T_31 ? 1'h0 : _signals_T_250; // @[Lookup.scala 34:39]
  wire  _signals_T_256 = _signals_T_21 ? 1'h0 : _signals_T_23 | (_signals_T_25 | (_signals_T_27 | (_signals_T_29 |
    _signals_T_251))); // @[Lookup.scala 34:39]
  wire  _signals_T_257 = _signals_T_19 ? 1'h0 : _signals_T_256; // @[Lookup.scala 34:39]
  wire  _signals_T_258 = _signals_T_17 ? 1'h0 : _signals_T_257; // @[Lookup.scala 34:39]
  wire  _signals_T_274 = _signals_T_117 ? 1'h0 : _signals_T_119 | (_signals_T_121 | (_signals_T_123 | (_signals_T_125 |
    (_signals_T_127 | (_signals_T_129 | _signals_T_131))))); // @[Lookup.scala 34:39]
  wire  _signals_T_275 = _signals_T_115 ? 1'h0 : _signals_T_274; // @[Lookup.scala 34:39]
  wire  _signals_T_276 = _signals_T_113 ? 1'h0 : _signals_T_275; // @[Lookup.scala 34:39]
  wire  _signals_T_277 = _signals_T_111 ? 1'h0 : _signals_T_276; // @[Lookup.scala 34:39]
  wire  _signals_T_278 = _signals_T_109 ? 1'h0 : _signals_T_277; // @[Lookup.scala 34:39]
  wire  _signals_T_279 = _signals_T_107 ? 1'h0 : _signals_T_278; // @[Lookup.scala 34:39]
  wire  _signals_T_280 = _signals_T_105 ? 1'h0 : _signals_T_279; // @[Lookup.scala 34:39]
  wire  _signals_T_281 = _signals_T_103 ? 1'h0 : _signals_T_280; // @[Lookup.scala 34:39]
  wire  _signals_T_282 = _signals_T_101 ? 1'h0 : _signals_T_281; // @[Lookup.scala 34:39]
  wire  _signals_T_283 = _signals_T_99 ? 1'h0 : _signals_T_282; // @[Lookup.scala 34:39]
  wire  _signals_T_284 = _signals_T_97 ? 1'h0 : _signals_T_283; // @[Lookup.scala 34:39]
  wire  _signals_T_285 = _signals_T_95 ? 1'h0 : _signals_T_284; // @[Lookup.scala 34:39]
  wire  _signals_T_286 = _signals_T_93 ? 1'h0 : _signals_T_285; // @[Lookup.scala 34:39]
  wire  _signals_T_287 = _signals_T_91 ? 1'h0 : _signals_T_286; // @[Lookup.scala 34:39]
  wire  _signals_T_288 = _signals_T_89 ? 1'h0 : _signals_T_287; // @[Lookup.scala 34:39]
  wire  _signals_T_289 = _signals_T_87 ? 1'h0 : _signals_T_288; // @[Lookup.scala 34:39]
  wire  _signals_T_290 = _signals_T_85 ? 1'h0 : _signals_T_289; // @[Lookup.scala 34:39]
  wire  _signals_T_291 = _signals_T_83 ? 1'h0 : _signals_T_290; // @[Lookup.scala 34:39]
  wire  _signals_T_294 = _signals_T_77 ? 1'h0 : _signals_T_79 | (_signals_T_81 | _signals_T_291); // @[Lookup.scala 34:39]
  wire  _signals_T_295 = _signals_T_75 ? 1'h0 : _signals_T_294; // @[Lookup.scala 34:39]
  wire  _signals_T_296 = _signals_T_73 ? 1'h0 : _signals_T_295; // @[Lookup.scala 34:39]
  wire  _signals_T_297 = _signals_T_71 ? 1'h0 : _signals_T_296; // @[Lookup.scala 34:39]
  wire  _signals_T_298 = _signals_T_69 ? 1'h0 : _signals_T_297; // @[Lookup.scala 34:39]
  wire  _signals_T_299 = _signals_T_67 ? 1'h0 : _signals_T_298; // @[Lookup.scala 34:39]
  wire  _signals_T_308 = _signals_T_49 ? 1'h0 : _signals_T_51 | (_signals_T_53 | (_signals_T_55 | (_signals_T_57 | (
    _signals_T_59 | (_signals_T_61 | (_signals_T_63 | (_signals_T_65 | _signals_T_299))))))); // @[Lookup.scala 34:39]
  wire  _signals_T_309 = _signals_T_47 ? 1'h0 : _signals_T_308; // @[Lookup.scala 34:39]
  wire  _signals_T_313 = _signals_T_39 ? 1'h0 : _signals_T_41 | (_signals_T_43 | (_signals_T_45 | _signals_T_309)); // @[Lookup.scala 34:39]
  wire  _signals_T_314 = _signals_T_37 ? 1'h0 : _signals_T_313; // @[Lookup.scala 34:39]
  wire  _signals_T_315 = _signals_T_35 ? 1'h0 : _signals_T_314; // @[Lookup.scala 34:39]
  wire  _signals_T_316 = _signals_T_33 ? 1'h0 : _signals_T_315; // @[Lookup.scala 34:39]
  wire  _signals_T_317 = _signals_T_31 ? 1'h0 : _signals_T_316; // @[Lookup.scala 34:39]
  wire  _signals_T_318 = _signals_T_29 ? 1'h0 : _signals_T_317; // @[Lookup.scala 34:39]
  wire  _signals_T_319 = _signals_T_27 ? 1'h0 : _signals_T_318; // @[Lookup.scala 34:39]
  wire  _signals_T_320 = _signals_T_25 ? 1'h0 : _signals_T_319; // @[Lookup.scala 34:39]
  wire  _signals_T_321 = _signals_T_23 ? 1'h0 : _signals_T_320; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_332 = _signals_T_133 ? 4'h1 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_333 = _signals_T_131 ? 4'h4 : _signals_T_332; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_334 = _signals_T_129 ? 4'h4 : _signals_T_333; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_335 = _signals_T_127 ? 4'h4 : _signals_T_334; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_336 = _signals_T_125 ? 4'h4 : _signals_T_335; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_337 = _signals_T_123 ? 4'h4 : _signals_T_336; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_338 = _signals_T_121 ? 4'h4 : _signals_T_337; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_339 = _signals_T_119 ? 4'h4 : _signals_T_338; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_340 = _signals_T_117 ? 4'h4 : _signals_T_339; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_341 = _signals_T_115 ? 4'h4 : _signals_T_340; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_342 = _signals_T_113 ? 4'h4 : _signals_T_341; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_343 = _signals_T_111 ? 4'h4 : _signals_T_342; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_344 = _signals_T_109 ? 4'h4 : _signals_T_343; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_345 = _signals_T_107 ? 4'h7 : _signals_T_344; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_346 = _signals_T_105 ? 4'h7 : _signals_T_345; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_347 = _signals_T_103 ? 4'h7 : _signals_T_346; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_348 = _signals_T_101 ? 4'h6 : _signals_T_347; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_349 = _signals_T_99 ? 4'h6 : _signals_T_348; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_350 = _signals_T_97 ? 4'h6 : _signals_T_349; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_351 = _signals_T_95 ? 4'h6 : _signals_T_350; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_352 = _signals_T_93 ? 4'h5 : _signals_T_351; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_353 = _signals_T_91 ? 4'h5 : _signals_T_352; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_354 = _signals_T_89 ? 4'h5 : _signals_T_353; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_355 = _signals_T_87 ? 4'h5 : _signals_T_354; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_356 = _signals_T_85 ? 4'h5 : _signals_T_355; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_357 = _signals_T_83 ? 4'h5 : _signals_T_356; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_358 = _signals_T_81 ? 4'h5 : _signals_T_357; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_359 = _signals_T_79 ? 4'h5 : _signals_T_358; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_360 = _signals_T_77 ? 4'h5 : _signals_T_359; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_361 = _signals_T_75 ? 4'h5 : _signals_T_360; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_362 = _signals_T_73 ? 4'h5 : _signals_T_361; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_363 = _signals_T_71 ? 4'h5 : _signals_T_362; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_364 = _signals_T_69 ? 4'h1 : _signals_T_363; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_365 = _signals_T_67 ? 4'h1 : _signals_T_364; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_366 = _signals_T_65 ? 4'hc : _signals_T_365; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_367 = _signals_T_63 ? 4'hc : _signals_T_366; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_368 = _signals_T_61 ? 4'hb : _signals_T_367; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_369 = _signals_T_59 ? 4'hb : _signals_T_368; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_370 = _signals_T_57 ? 4'h1 : _signals_T_369; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_371 = _signals_T_55 ? 4'h1 : _signals_T_370; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_372 = _signals_T_53 ? 4'h1 : _signals_T_371; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_373 = _signals_T_51 ? 4'h1 : _signals_T_372; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_374 = _signals_T_49 ? 4'h1 : _signals_T_373; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_375 = _signals_T_47 ? 4'h1 : _signals_T_374; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_376 = _signals_T_45 ? 4'h1 : _signals_T_375; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_377 = _signals_T_43 ? 4'h1 : _signals_T_376; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_378 = _signals_T_41 ? 4'h2 : _signals_T_377; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_379 = _signals_T_39 ? 4'h3 : _signals_T_378; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_380 = _signals_T_37 ? 4'h9 : _signals_T_379; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_381 = _signals_T_35 ? 4'h9 : _signals_T_380; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_382 = _signals_T_33 ? 4'ha : _signals_T_381; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_383 = _signals_T_31 ? 4'ha : _signals_T_382; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_384 = _signals_T_29 ? 4'h1 : _signals_T_383; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_385 = _signals_T_27 ? 4'h1 : _signals_T_384; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_386 = _signals_T_25 ? 4'h1 : _signals_T_385; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_387 = _signals_T_23 ? 4'h1 : _signals_T_386; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_388 = _signals_T_21 ? 4'h1 : _signals_T_387; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_389 = _signals_T_19 ? 4'h1 : _signals_T_388; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_390 = _signals_T_17 ? 4'h1 : _signals_T_389; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_391 = _signals_T_15 ? 4'h1 : _signals_T_390; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_392 = _signals_T_13 ? 4'h1 : _signals_T_391; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_393 = _signals_T_11 ? 4'h1 : _signals_T_392; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_394 = _signals_T_9 ? 4'h1 : _signals_T_393; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_395 = _signals_T_7 ? 4'h1 : _signals_T_394; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_396 = _signals_T_5 ? 4'h1 : _signals_T_395; // @[Lookup.scala 34:39]
  wire [3:0] _signals_T_397 = _signals_T_3 ? 4'h1 : _signals_T_396; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_398 = _signals_T_133 ? 7'h4c : 7'h0; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_399 = _signals_T_131 ? 7'h3d : _signals_T_398; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_400 = _signals_T_129 ? 7'h3c : _signals_T_399; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_401 = _signals_T_127 ? 7'h37 : _signals_T_400; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_402 = _signals_T_125 ? 7'h36 : _signals_T_401; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_403 = _signals_T_123 ? 7'h3b : _signals_T_402; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_404 = _signals_T_121 ? 7'h3a : _signals_T_403; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_405 = _signals_T_119 ? 7'h38 : _signals_T_404; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_406 = _signals_T_117 ? 7'h35 : _signals_T_405; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_407 = _signals_T_115 ? 7'h33 : _signals_T_406; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_408 = _signals_T_113 ? 7'h32 : _signals_T_407; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_409 = _signals_T_111 ? 7'h31 : _signals_T_408; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_410 = _signals_T_109 ? 7'h30 : _signals_T_409; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_411 = _signals_T_107 ? 7'h46 : _signals_T_410; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_412 = _signals_T_105 ? 7'h45 : _signals_T_411; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_413 = _signals_T_103 ? 7'h44 : _signals_T_412; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_414 = _signals_T_101 ? 7'h4b : _signals_T_413; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_415 = _signals_T_99 ? 7'h4a : _signals_T_414; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_416 = _signals_T_97 ? 7'h49 : _signals_T_415; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_417 = _signals_T_95 ? 7'h48 : _signals_T_416; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_418 = _signals_T_93 ? 7'h2e : _signals_T_417; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_419 = _signals_T_91 ? 7'h2d : _signals_T_418; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_420 = _signals_T_89 ? 7'h2a : _signals_T_419; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_421 = _signals_T_87 ? 7'h29 : _signals_T_420; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_422 = _signals_T_85 ? 7'h2c : _signals_T_421; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_423 = _signals_T_83 ? 7'h2b : _signals_T_422; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_424 = _signals_T_81 ? 7'h2f : _signals_T_423; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_425 = _signals_T_79 ? 7'h28 : _signals_T_424; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_426 = _signals_T_77 ? 7'h26 : _signals_T_425; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_427 = _signals_T_75 ? 7'h27 : _signals_T_426; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_428 = _signals_T_73 ? 7'h25 : _signals_T_427; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_429 = _signals_T_71 ? 7'h24 : _signals_T_428; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_430 = _signals_T_69 ? 7'h16 : _signals_T_429; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_431 = _signals_T_67 ? 7'h15 : _signals_T_430; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_432 = _signals_T_65 ? 7'h23 : _signals_T_431; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_433 = _signals_T_63 ? 7'h22 : _signals_T_432; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_434 = _signals_T_61 ? 7'h1c : _signals_T_433; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_435 = _signals_T_59 ? 7'h1b : _signals_T_434; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_436 = _signals_T_57 ? 7'h18 : _signals_T_435; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_437 = _signals_T_55 ? 7'h17 : _signals_T_436; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_438 = _signals_T_53 ? 7'h16 : _signals_T_437; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_439 = _signals_T_51 ? 7'h15 : _signals_T_438; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_440 = _signals_T_49 ? 7'h14 : _signals_T_439; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_441 = _signals_T_47 ? 7'h13 : _signals_T_440; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_442 = _signals_T_45 ? 7'h14 : _signals_T_441; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_443 = _signals_T_43 ? 7'h13 : _signals_T_442; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_444 = _signals_T_41 ? 7'h12 : _signals_T_443; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_445 = _signals_T_39 ? 7'h11 : _signals_T_444; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_446 = _signals_T_37 ? 7'h10 : _signals_T_445; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_447 = _signals_T_35 ? 7'he : _signals_T_446; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_448 = _signals_T_33 ? 7'hf : _signals_T_447; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_449 = _signals_T_31 ? 7'hd : _signals_T_448; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_450 = _signals_T_29 ? 7'h2 : _signals_T_449; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_451 = _signals_T_27 ? 7'h3 : _signals_T_450; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_452 = _signals_T_25 ? 7'h1 : _signals_T_451; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_453 = _signals_T_23 ? 7'h2 : _signals_T_452; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_454 = _signals_T_21 ? 7'h9 : _signals_T_453; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_455 = _signals_T_19 ? 7'h7 : _signals_T_454; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_456 = _signals_T_17 ? 7'h5 : _signals_T_455; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_457 = _signals_T_15 ? 7'h9 : _signals_T_456; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_458 = _signals_T_13 ? 7'h7 : _signals_T_457; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_459 = _signals_T_11 ? 7'h5 : _signals_T_458; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_460 = _signals_T_9 ? 7'h4 : _signals_T_459; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_461 = _signals_T_7 ? 7'h3 : _signals_T_460; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_462 = _signals_T_5 ? 7'h1 : _signals_T_461; // @[Lookup.scala 34:39]
  wire [6:0] _signals_T_463 = _signals_T_3 ? 7'h2 : _signals_T_462; // @[Lookup.scala 34:39]
  wire  _signals_T_469 = _signals_T_123 ? 1'h0 : _signals_T_125 | _signals_T_127; // @[Lookup.scala 34:39]
  wire  _signals_T_470 = _signals_T_121 ? 1'h0 : _signals_T_469; // @[Lookup.scala 34:39]
  wire  _signals_T_471 = _signals_T_119 ? 1'h0 : _signals_T_470; // @[Lookup.scala 34:39]
  wire  _signals_T_477 = _signals_T_107 ? 1'h0 : _signals_T_109 | (_signals_T_111 | (_signals_T_113 | (_signals_T_115 |
    (_signals_T_117 | _signals_T_471)))); // @[Lookup.scala 34:39]
  wire  _signals_T_478 = _signals_T_105 ? 1'h0 : _signals_T_477; // @[Lookup.scala 34:39]
  wire  _signals_T_479 = _signals_T_103 ? 1'h0 : _signals_T_478; // @[Lookup.scala 34:39]
  wire  _signals_T_480 = _signals_T_101 ? 1'h0 : _signals_T_479; // @[Lookup.scala 34:39]
  wire  _signals_T_481 = _signals_T_99 ? 1'h0 : _signals_T_480; // @[Lookup.scala 34:39]
  wire  _signals_T_482 = _signals_T_97 ? 1'h0 : _signals_T_481; // @[Lookup.scala 34:39]
  wire  _signals_T_483 = _signals_T_95 ? 1'h0 : _signals_T_482; // @[Lookup.scala 34:39]
  wire  _signals_T_485 = _signals_T_91 ? 1'h0 : _signals_T_93 | _signals_T_483; // @[Lookup.scala 34:39]
  wire  _signals_T_487 = _signals_T_87 ? 1'h0 : _signals_T_89 | _signals_T_485; // @[Lookup.scala 34:39]
  wire  _signals_T_488 = _signals_T_85 ? 1'h0 : _signals_T_487; // @[Lookup.scala 34:39]
  wire  _signals_T_489 = _signals_T_83 ? 1'h0 : _signals_T_488; // @[Lookup.scala 34:39]
  wire  _signals_T_490 = _signals_T_81 ? 1'h0 : _signals_T_489; // @[Lookup.scala 34:39]
  wire  _signals_T_491 = _signals_T_79 ? 1'h0 : _signals_T_490; // @[Lookup.scala 34:39]
  wire  _signals_T_493 = _signals_T_75 ? 1'h0 : _signals_T_77 | _signals_T_491; // @[Lookup.scala 34:39]
  wire  _signals_T_495 = _signals_T_71 ? 1'h0 : _signals_T_73 | _signals_T_493; // @[Lookup.scala 34:39]
  wire  _signals_T_498 = _signals_T_65 ? 1'h0 : _signals_T_67 | (_signals_T_69 | _signals_T_495); // @[Lookup.scala 34:39]
  wire  _signals_T_499 = _signals_T_63 ? 1'h0 : _signals_T_498; // @[Lookup.scala 34:39]
  wire  _signals_T_500 = _signals_T_61 ? 1'h0 : _signals_T_499; // @[Lookup.scala 34:39]
  wire  _signals_T_501 = _signals_T_59 ? 1'h0 : _signals_T_500; // @[Lookup.scala 34:39]
  wire  _signals_T_510 = _signals_T_41 ? 1'h0 : _signals_T_43 | (_signals_T_45 | (_signals_T_47 | (_signals_T_49 | (
    _signals_T_51 | (_signals_T_53 | (_signals_T_55 | (_signals_T_57 | _signals_T_501))))))); // @[Lookup.scala 34:39]
  wire  _signals_T_512 = _signals_T_37 ? 1'h0 : _signals_T_39 | _signals_T_510; // @[Lookup.scala 34:39]
  wire  _signals_T_513 = _signals_T_35 ? 1'h0 : _signals_T_512; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_533 = _signals_T_127 ? 2'h1 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_534 = _signals_T_125 ? 2'h1 : _signals_T_533; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_535 = _signals_T_123 ? 2'h0 : _signals_T_534; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_536 = _signals_T_121 ? 2'h0 : _signals_T_535; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_537 = _signals_T_119 ? 2'h0 : _signals_T_536; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_538 = _signals_T_117 ? 2'h1 : _signals_T_537; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_539 = _signals_T_115 ? 2'h1 : _signals_T_538; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_540 = _signals_T_113 ? 2'h1 : _signals_T_539; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_541 = _signals_T_111 ? 2'h1 : _signals_T_540; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_542 = _signals_T_109 ? 2'h1 : _signals_T_541; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_543 = _signals_T_107 ? 2'h0 : _signals_T_542; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_544 = _signals_T_105 ? 2'h0 : _signals_T_543; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_545 = _signals_T_103 ? 2'h0 : _signals_T_544; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_546 = _signals_T_101 ? 2'h0 : _signals_T_545; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_547 = _signals_T_99 ? 2'h0 : _signals_T_546; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_548 = _signals_T_97 ? 2'h0 : _signals_T_547; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_549 = _signals_T_95 ? 2'h0 : _signals_T_548; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_550 = _signals_T_93 ? 2'h2 : _signals_T_549; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_551 = _signals_T_91 ? 2'h0 : _signals_T_550; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_552 = _signals_T_89 ? 2'h2 : _signals_T_551; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_553 = _signals_T_87 ? 2'h0 : _signals_T_552; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_554 = _signals_T_85 ? 2'h0 : _signals_T_553; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_555 = _signals_T_83 ? 2'h0 : _signals_T_554; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_556 = _signals_T_81 ? 2'h0 : _signals_T_555; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_557 = _signals_T_79 ? 2'h0 : _signals_T_556; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_558 = _signals_T_77 ? 2'h0 : _signals_T_557; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_559 = _signals_T_75 ? 2'h0 : _signals_T_558; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_560 = _signals_T_73 ? 2'h2 : _signals_T_559; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_561 = _signals_T_71 ? 2'h0 : _signals_T_560; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_562 = _signals_T_69 ? 2'h1 : _signals_T_561; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_563 = _signals_T_67 ? 2'h1 : _signals_T_562; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_564 = _signals_T_65 ? 2'h0 : _signals_T_563; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_565 = _signals_T_63 ? 2'h0 : _signals_T_564; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_566 = _signals_T_61 ? 2'h0 : _signals_T_565; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_567 = _signals_T_59 ? 2'h0 : _signals_T_566; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_568 = _signals_T_57 ? 2'h0 : _signals_T_567; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_569 = _signals_T_55 ? 2'h0 : _signals_T_568; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_570 = _signals_T_53 ? 2'h0 : _signals_T_569; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_571 = _signals_T_51 ? 2'h0 : _signals_T_570; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_572 = _signals_T_49 ? 2'h1 : _signals_T_571; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_573 = _signals_T_47 ? 2'h1 : _signals_T_572; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_574 = _signals_T_45 ? 2'h0 : _signals_T_573; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_575 = _signals_T_43 ? 2'h0 : _signals_T_574; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_576 = _signals_T_41 ? 2'h0 : _signals_T_575; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_577 = _signals_T_39 ? 2'h1 : _signals_T_576; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_578 = _signals_T_37 ? 2'h0 : _signals_T_577; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_579 = _signals_T_35 ? 2'h0 : _signals_T_578; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_580 = _signals_T_33 ? 2'h0 : _signals_T_579; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_581 = _signals_T_31 ? 2'h0 : _signals_T_580; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_582 = _signals_T_29 ? 2'h1 : _signals_T_581; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_583 = _signals_T_27 ? 2'h1 : _signals_T_582; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_584 = _signals_T_25 ? 2'h1 : _signals_T_583; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_585 = _signals_T_23 ? 2'h1 : _signals_T_584; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_586 = _signals_T_21 ? 2'h0 : _signals_T_585; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_587 = _signals_T_19 ? 2'h0 : _signals_T_586; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_588 = _signals_T_17 ? 2'h0 : _signals_T_587; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_589 = _signals_T_15 ? 2'h0 : _signals_T_588; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_590 = _signals_T_13 ? 2'h0 : _signals_T_589; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_591 = _signals_T_11 ? 2'h0 : _signals_T_590; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_592 = _signals_T_9 ? 2'h0 : _signals_T_591; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_593 = _signals_T_7 ? 2'h0 : _signals_T_592; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_594 = _signals_T_5 ? 2'h0 : _signals_T_593; // @[Lookup.scala 34:39]
  wire [1:0] _signals_T_595 = _signals_T_3 ? 2'h0 : _signals_T_594; // @[Lookup.scala 34:39]
  wire [1:0] reg_waddr_type = _signals_T_1 ? 2'h0 : _signals_T_595; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_628 = _signals_T_69 ? 3'h1 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_629 = _signals_T_67 ? 3'h1 : _signals_T_628; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_630 = _signals_T_65 ? 3'h0 : _signals_T_629; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_631 = _signals_T_63 ? 3'h0 : _signals_T_630; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_632 = _signals_T_61 ? 3'h0 : _signals_T_631; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_633 = _signals_T_59 ? 3'h0 : _signals_T_632; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_634 = _signals_T_57 ? 3'h0 : _signals_T_633; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_635 = _signals_T_55 ? 3'h0 : _signals_T_634; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_636 = _signals_T_53 ? 3'h0 : _signals_T_635; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_637 = _signals_T_51 ? 3'h0 : _signals_T_636; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_638 = _signals_T_49 ? 3'h1 : _signals_T_637; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_639 = _signals_T_47 ? 3'h1 : _signals_T_638; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_640 = _signals_T_45 ? 3'h0 : _signals_T_639; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_641 = _signals_T_43 ? 3'h0 : _signals_T_640; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_642 = _signals_T_41 ? 3'h0 : _signals_T_641; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_643 = _signals_T_39 ? 3'h0 : _signals_T_642; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_644 = _signals_T_37 ? 3'h0 : _signals_T_643; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_645 = _signals_T_35 ? 3'h0 : _signals_T_644; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_646 = _signals_T_33 ? 3'h0 : _signals_T_645; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_647 = _signals_T_31 ? 3'h0 : _signals_T_646; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_648 = _signals_T_29 ? 3'h3 : _signals_T_647; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_649 = _signals_T_27 ? 3'h2 : _signals_T_648; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_650 = _signals_T_25 ? 3'h2 : _signals_T_649; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_651 = _signals_T_23 ? 3'h2 : _signals_T_650; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_652 = _signals_T_21 ? 3'h4 : _signals_T_651; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_653 = _signals_T_19 ? 3'h4 : _signals_T_652; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_654 = _signals_T_17 ? 3'h4 : _signals_T_653; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_655 = _signals_T_15 ? 3'h0 : _signals_T_654; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_656 = _signals_T_13 ? 3'h0 : _signals_T_655; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_657 = _signals_T_11 ? 3'h0 : _signals_T_656; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_658 = _signals_T_9 ? 3'h0 : _signals_T_657; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_659 = _signals_T_7 ? 3'h0 : _signals_T_658; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_660 = _signals_T_5 ? 3'h0 : _signals_T_659; // @[Lookup.scala 34:39]
  wire [2:0] _signals_T_661 = _signals_T_3 ? 3'h0 : _signals_T_660; // @[Lookup.scala 34:39]
  wire [2:0] imm_type = _signals_T_1 ? 3'h0 : _signals_T_661; // @[Lookup.scala 34:39]
  wire  _signals_T_675 = _signals_T_107 ? 1'h0 : _signals_T_109 | (_signals_T_111 | (_signals_T_113 | (_signals_T_115 |
    (_signals_T_117 | (_signals_T_119 | (_signals_T_121 | (_signals_T_123 | (_signals_T_125 | (_signals_T_127 | (
    _signals_T_129 | (_signals_T_131 | _signals_T_134))))))))))); // @[Lookup.scala 34:39]
  wire  _signals_T_676 = _signals_T_105 ? 1'h0 : _signals_T_675; // @[Lookup.scala 34:39]
  wire  _signals_T_677 = _signals_T_103 ? 1'h0 : _signals_T_676; // @[Lookup.scala 34:39]
  wire  _signals_T_678 = _signals_T_101 ? 1'h0 : _signals_T_677; // @[Lookup.scala 34:39]
  wire  _signals_T_679 = _signals_T_99 ? 1'h0 : _signals_T_678; // @[Lookup.scala 34:39]
  wire  _signals_T_680 = _signals_T_97 ? 1'h0 : _signals_T_679; // @[Lookup.scala 34:39]
  wire  _signals_T_681 = _signals_T_95 ? 1'h0 : _signals_T_680; // @[Lookup.scala 34:39]
  wire  _signals_T_708 = _signals_T_41 ? 1'h0 : _signals_T_43 | (_signals_T_45 | (_signals_T_47 | (_signals_T_49 | (
    _signals_T_51 | (_signals_T_53 | (_signals_T_55 | (_signals_T_57 | (_signals_T_59 | (_signals_T_61 | (_signals_T_63
     | (_signals_T_65 | (_signals_T_67 | (_signals_T_69 | (_signals_T_71 | (_signals_T_73 | (_signals_T_75 | (
    _signals_T_77 | (_signals_T_79 | (_signals_T_81 | (_signals_T_83 | (_signals_T_85 | (_signals_T_87 | (_signals_T_89
     | (_signals_T_91 | (_signals_T_93 | _signals_T_681))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _signals_T_709 = _signals_T_39 ? 1'h0 : _signals_T_708; // @[Lookup.scala 34:39]
  wire [4:0] rt = io_in_inst[20:16]; // @[Decoder.scala 152:19]
  wire [4:0] rd = io_in_inst[15:11]; // @[Decoder.scala 153:19]
  wire [4:0] sa = io_in_inst[10:6]; // @[Decoder.scala 154:19]
  wire [15:0] imm16 = io_in_inst[15:0]; // @[Decoder.scala 156:19]
  wire [4:0] _io_out_reg_waddr_T_1 = 2'h0 == reg_waddr_type ? rd : 5'h1f; // @[Mux.scala 81:58]
  wire [31:0] _io_out_imm32_T_1 = {27'h0,sa}; // @[Cat.scala 33:92]
  wire [15:0] _io_out_imm32_T_4 = imm16[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_out_imm32_T_5 = {_io_out_imm32_T_4,imm16}; // @[Cat.scala 33:92]
  wire [31:0] _io_out_imm32_T_7 = {16'h0,imm16}; // @[Cat.scala 33:92]
  wire [31:0] _io_out_imm32_T_9 = {imm16,16'h0}; // @[Cat.scala 33:92]
  wire [31:0] _io_out_imm32_T_11 = 3'h1 == imm_type ? _io_out_imm32_T_5 : _io_out_imm32_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_out_imm32_T_13 = 3'h2 == imm_type ? _io_out_imm32_T_7 : _io_out_imm32_T_11; // @[Mux.scala 81:58]
  assign io_out_inst_valid = _signals_T_1 ? 1'h0 : _signals_T_199; // @[Lookup.scala 34:39]
  assign io_out_reg1_ren = _signals_T_1 ? 1'h0 : _signals_T_3 | (_signals_T_5 | (_signals_T_7 | (_signals_T_9 | (
    _signals_T_11 | (_signals_T_13 | (_signals_T_15 | _signals_T_258)))))); // @[Lookup.scala 34:39]
  assign io_out_reg1_raddr = io_in_inst[25:21]; // @[Decoder.scala 155:19]
  assign io_out_reg2_ren = _signals_T_1 ? 1'h0 : _signals_T_3 | (_signals_T_5 | (_signals_T_7 | (_signals_T_9 | (
    _signals_T_11 | (_signals_T_13 | (_signals_T_15 | (_signals_T_17 | (_signals_T_19 | (_signals_T_21 | _signals_T_321)
    )))))))); // @[Lookup.scala 34:39]
  assign io_out_reg2_raddr = io_in_inst[20:16]; // @[Decoder.scala 152:19]
  assign io_out_fusel = _signals_T_1 ? 4'h0 : _signals_T_397; // @[Lookup.scala 34:39]
  assign io_out_op = _signals_T_1 ? 7'h0 : _signals_T_463; // @[Lookup.scala 34:39]
  assign io_out_reg_wen = _signals_T_1 ? 1'h0 : _signals_T_3 | (_signals_T_5 | (_signals_T_7 | (_signals_T_9 | (
    _signals_T_11 | (_signals_T_13 | (_signals_T_15 | (_signals_T_17 | (_signals_T_19 | (_signals_T_21 | (_signals_T_23
     | (_signals_T_25 | (_signals_T_27 | (_signals_T_29 | (_signals_T_31 | (_signals_T_33 | _signals_T_513))))))))))))))
    ); // @[Lookup.scala 34:39]
  assign io_out_reg_waddr = 2'h1 == reg_waddr_type ? rt : _io_out_reg_waddr_T_1; // @[Mux.scala 81:58]
  assign io_out_imm32 = 3'h3 == imm_type ? _io_out_imm32_T_9 : _io_out_imm32_T_13; // @[Mux.scala 81:58]
  assign io_out_cp0_addr = {rd,io_in_inst[2:0]}; // @[Cat.scala 33:92]
  assign io_out_dual_issue = _signals_T_1 | (_signals_T_3 | (_signals_T_5 | (_signals_T_7 | (_signals_T_9 | (
    _signals_T_11 | (_signals_T_13 | (_signals_T_15 | (_signals_T_17 | (_signals_T_19 | (_signals_T_21 | (_signals_T_23
     | (_signals_T_25 | (_signals_T_27 | (_signals_T_29 | (_signals_T_31 | (_signals_T_33 | (_signals_T_35 | (
    _signals_T_37 | _signals_T_709)))))))))))))))))); // @[Lookup.scala 34:39]
  assign io_out_inst = io_in_inst; // @[Decoder.scala 185:21]
endmodule
module JumpCtrl(
  input         io_in_allow_to_go,
  input  [31:0] io_in_pc,
  input  [4:0]  io_in_decoded_inst0_reg1_raddr,
  input  [6:0]  io_in_decoded_inst0_op,
  input  [31:0] io_in_decoded_inst0_inst,
  input  [31:0] io_in_reg1_data,
  input         io_in_forward_0_exe_wen,
  input  [4:0]  io_in_forward_0_exe_waddr,
  input         io_in_forward_0_mem_wen,
  input  [4:0]  io_in_forward_0_mem_waddr,
  input         io_in_forward_1_exe_wen,
  input  [4:0]  io_in_forward_1_exe_waddr,
  input         io_in_forward_1_mem_wen,
  input  [4:0]  io_in_forward_1_mem_waddr,
  output        io_out_inst_is_jump,
  output        io_out_jump_register,
  output        io_out_jump_flag,
  output [31:0] io_out_jump_target
);
  wire  inst_is_j = 7'h24 == io_in_decoded_inst0_op | 7'h25 == io_in_decoded_inst0_op; // @[JumpCtrl.scala 28:52]
  wire  inst_is_jr = 7'h27 == io_in_decoded_inst0_op | 7'h26 == io_in_decoded_inst0_op; // @[JumpCtrl.scala 29:54]
  wire  _io_out_jump_register_T_3 = io_in_forward_1_exe_wen & io_in_decoded_inst0_reg1_raddr ==
    io_in_forward_1_exe_waddr; // @[JumpCtrl.scala 34:33]
  wire  _io_out_jump_register_T_4 = io_in_forward_0_exe_wen & io_in_decoded_inst0_reg1_raddr ==
    io_in_forward_0_exe_waddr | _io_out_jump_register_T_3; // @[JumpCtrl.scala 33:98]
  wire  _io_out_jump_register_T_6 = io_in_forward_0_mem_wen & io_in_decoded_inst0_reg1_raddr ==
    io_in_forward_0_mem_waddr; // @[JumpCtrl.scala 35:33]
  wire  _io_out_jump_register_T_7 = _io_out_jump_register_T_4 | _io_out_jump_register_T_6; // @[JumpCtrl.scala 34:99]
  wire  _io_out_jump_register_T_9 = io_in_forward_1_mem_wen & io_in_decoded_inst0_reg1_raddr ==
    io_in_forward_1_mem_waddr; // @[JumpCtrl.scala 36:33]
  wire  _io_out_jump_register_T_10 = _io_out_jump_register_T_7 | _io_out_jump_register_T_9; // @[JumpCtrl.scala 35:99]
  wire [31:0] pc_plus_4 = io_in_pc + 32'h4; // @[JumpCtrl.scala 37:28]
  wire [31:0] _io_out_jump_target_T_2 = {pc_plus_4[31:28],io_in_decoded_inst0_inst[25:0],2'h0}; // @[Cat.scala 33:92]
  assign io_out_inst_is_jump = inst_is_j | inst_is_jr; // @[JumpCtrl.scala 30:36]
  assign io_out_jump_register = inst_is_jr & _io_out_jump_register_T_10; // @[JumpCtrl.scala 32:38]
  assign io_out_jump_flag = io_in_allow_to_go & (inst_is_j | inst_is_jr & ~io_out_jump_register); // @[JumpCtrl.scala 31:44]
  assign io_out_jump_target = inst_is_j ? _io_out_jump_target_T_2 : io_in_reg1_data; // @[JumpCtrl.scala 38:28]
endmodule
module ForwardCtrl(
  input         io_in_forward_0_exe_wen,
  input  [4:0]  io_in_forward_0_exe_waddr,
  input  [31:0] io_in_forward_0_exe_wdata,
  input         io_in_forward_0_exe_mem_ren,
  input         io_in_forward_0_mem_wen,
  input  [4:0]  io_in_forward_0_mem_waddr,
  input  [31:0] io_in_forward_0_mem_wdata,
  input         io_in_forward_1_exe_wen,
  input  [4:0]  io_in_forward_1_exe_waddr,
  input  [31:0] io_in_forward_1_exe_wdata,
  input         io_in_forward_1_exe_mem_ren,
  input         io_in_forward_1_mem_wen,
  input  [4:0]  io_in_forward_1_mem_waddr,
  input  [31:0] io_in_forward_1_mem_wdata,
  input  [4:0]  io_in_regfile_0_src1_raddr,
  input  [31:0] io_in_regfile_0_src1_rdata,
  input  [4:0]  io_in_regfile_0_src2_raddr,
  input  [31:0] io_in_regfile_0_src2_rdata,
  input  [4:0]  io_in_regfile_1_src1_raddr,
  input  [31:0] io_in_regfile_1_src1_rdata,
  input  [4:0]  io_in_regfile_1_src2_raddr,
  input  [31:0] io_in_regfile_1_src2_rdata,
  output [31:0] io_out_inst_0_src1_rdata,
  output [31:0] io_out_inst_0_src2_rdata,
  output [31:0] io_out_inst_1_src1_rdata,
  output [31:0] io_out_inst_1_src2_rdata
);
  wire  _T = io_in_forward_0_mem_waddr == io_in_regfile_0_src1_raddr; // @[ForwardCtrl.scala 34:38]
  wire  _T_1 = io_in_forward_0_mem_wen & _T; // @[ForwardCtrl.scala 33:34]
  wire [31:0] _GEN_0 = _T_1 ? io_in_forward_0_mem_wdata : io_in_regfile_0_src1_rdata; // @[ForwardCtrl.scala 25:31 35:9 36:35]
  wire  _T_2 = io_in_forward_0_mem_waddr == io_in_regfile_0_src2_raddr; // @[ForwardCtrl.scala 40:38]
  wire  _T_3 = io_in_forward_0_mem_wen & _T_2; // @[ForwardCtrl.scala 39:34]
  wire [31:0] _GEN_1 = _T_3 ? io_in_forward_0_mem_wdata : io_in_regfile_0_src2_rdata; // @[ForwardCtrl.scala 26:31 41:9 42:35]
  wire  _T_4 = io_in_forward_1_mem_waddr == io_in_regfile_0_src1_raddr; // @[ForwardCtrl.scala 34:38]
  wire  _T_5 = io_in_forward_1_mem_wen & _T_4; // @[ForwardCtrl.scala 33:34]
  wire [31:0] _GEN_2 = _T_5 ? io_in_forward_1_mem_wdata : _GEN_0; // @[ForwardCtrl.scala 35:9 36:35]
  wire  _T_6 = io_in_forward_1_mem_waddr == io_in_regfile_0_src2_raddr; // @[ForwardCtrl.scala 40:38]
  wire  _T_7 = io_in_forward_1_mem_wen & _T_6; // @[ForwardCtrl.scala 39:34]
  wire [31:0] _GEN_3 = _T_7 ? io_in_forward_1_mem_wdata : _GEN_1; // @[ForwardCtrl.scala 41:9 42:35]
  wire  _T_8 = io_in_forward_0_mem_waddr == io_in_regfile_1_src1_raddr; // @[ForwardCtrl.scala 34:38]
  wire  _T_9 = io_in_forward_0_mem_wen & _T_8; // @[ForwardCtrl.scala 33:34]
  wire [31:0] _GEN_4 = _T_9 ? io_in_forward_0_mem_wdata : io_in_regfile_1_src1_rdata; // @[ForwardCtrl.scala 25:31 35:9 36:35]
  wire  _T_10 = io_in_forward_0_mem_waddr == io_in_regfile_1_src2_raddr; // @[ForwardCtrl.scala 40:38]
  wire  _T_11 = io_in_forward_0_mem_wen & _T_10; // @[ForwardCtrl.scala 39:34]
  wire [31:0] _GEN_5 = _T_11 ? io_in_forward_0_mem_wdata : io_in_regfile_1_src2_rdata; // @[ForwardCtrl.scala 26:31 41:9 42:35]
  wire  _T_12 = io_in_forward_1_mem_waddr == io_in_regfile_1_src1_raddr; // @[ForwardCtrl.scala 34:38]
  wire  _T_13 = io_in_forward_1_mem_wen & _T_12; // @[ForwardCtrl.scala 33:34]
  wire [31:0] _GEN_6 = _T_13 ? io_in_forward_1_mem_wdata : _GEN_4; // @[ForwardCtrl.scala 35:9 36:35]
  wire  _T_14 = io_in_forward_1_mem_waddr == io_in_regfile_1_src2_raddr; // @[ForwardCtrl.scala 40:38]
  wire  _T_15 = io_in_forward_1_mem_wen & _T_14; // @[ForwardCtrl.scala 39:34]
  wire [31:0] _GEN_7 = _T_15 ? io_in_forward_1_mem_wdata : _GEN_5; // @[ForwardCtrl.scala 41:9 42:35]
  wire  _T_17 = io_in_forward_0_exe_wen & ~io_in_forward_0_exe_mem_ren; // @[ForwardCtrl.scala 51:34]
  wire  _T_18 = io_in_forward_0_exe_waddr == io_in_regfile_0_src1_raddr; // @[ForwardCtrl.scala 52:38]
  wire  _T_19 = io_in_forward_0_exe_wen & ~io_in_forward_0_exe_mem_ren & _T_18; // @[ForwardCtrl.scala 51:67]
  wire [31:0] _GEN_8 = _T_19 ? io_in_forward_0_exe_wdata : _GEN_2; // @[ForwardCtrl.scala 53:9 54:35]
  wire  _T_22 = io_in_forward_0_exe_waddr == io_in_regfile_0_src2_raddr; // @[ForwardCtrl.scala 58:38]
  wire  _T_23 = _T_17 & _T_22; // @[ForwardCtrl.scala 57:67]
  wire [31:0] _GEN_9 = _T_23 ? io_in_forward_0_exe_wdata : _GEN_3; // @[ForwardCtrl.scala 59:9 60:35]
  wire  _T_25 = io_in_forward_1_exe_wen & ~io_in_forward_1_exe_mem_ren; // @[ForwardCtrl.scala 51:34]
  wire  _T_26 = io_in_forward_1_exe_waddr == io_in_regfile_0_src1_raddr; // @[ForwardCtrl.scala 52:38]
  wire  _T_27 = io_in_forward_1_exe_wen & ~io_in_forward_1_exe_mem_ren & _T_26; // @[ForwardCtrl.scala 51:67]
  wire  _T_30 = io_in_forward_1_exe_waddr == io_in_regfile_0_src2_raddr; // @[ForwardCtrl.scala 58:38]
  wire  _T_31 = _T_25 & _T_30; // @[ForwardCtrl.scala 57:67]
  wire  _T_34 = io_in_forward_0_exe_waddr == io_in_regfile_1_src1_raddr; // @[ForwardCtrl.scala 52:38]
  wire  _T_35 = io_in_forward_0_exe_wen & ~io_in_forward_0_exe_mem_ren & _T_34; // @[ForwardCtrl.scala 51:67]
  wire [31:0] _GEN_12 = _T_35 ? io_in_forward_0_exe_wdata : _GEN_6; // @[ForwardCtrl.scala 53:9 54:35]
  wire  _T_38 = io_in_forward_0_exe_waddr == io_in_regfile_1_src2_raddr; // @[ForwardCtrl.scala 58:38]
  wire  _T_39 = _T_17 & _T_38; // @[ForwardCtrl.scala 57:67]
  wire [31:0] _GEN_13 = _T_39 ? io_in_forward_0_exe_wdata : _GEN_7; // @[ForwardCtrl.scala 59:9 60:35]
  wire  _T_42 = io_in_forward_1_exe_waddr == io_in_regfile_1_src1_raddr; // @[ForwardCtrl.scala 52:38]
  wire  _T_43 = io_in_forward_1_exe_wen & ~io_in_forward_1_exe_mem_ren & _T_42; // @[ForwardCtrl.scala 51:67]
  wire  _T_46 = io_in_forward_1_exe_waddr == io_in_regfile_1_src2_raddr; // @[ForwardCtrl.scala 58:38]
  wire  _T_47 = _T_25 & _T_46; // @[ForwardCtrl.scala 57:67]
  assign io_out_inst_0_src1_rdata = _T_27 ? io_in_forward_1_exe_wdata : _GEN_8; // @[ForwardCtrl.scala 53:9 54:35]
  assign io_out_inst_0_src2_rdata = _T_31 ? io_in_forward_1_exe_wdata : _GEN_9; // @[ForwardCtrl.scala 59:9 60:35]
  assign io_out_inst_1_src1_rdata = _T_43 ? io_in_forward_1_exe_wdata : _GEN_12; // @[ForwardCtrl.scala 53:9 54:35]
  assign io_out_inst_1_src2_rdata = _T_47 ? io_in_forward_1_exe_wdata : _GEN_13; // @[ForwardCtrl.scala 59:9 60:35]
endmodule
module DecoderUnit(
  output        io_instBuffer_inst_0_ready,
  input  [31:0] io_instBuffer_inst_0_bits_pc,
  input  [31:0] io_instBuffer_inst_0_bits_inst,
  input         io_instBuffer_inst_0_bits_tlb_invalid,
  output        io_instBuffer_inst_1_ready,
  input  [31:0] io_instBuffer_inst_1_bits_pc,
  input  [31:0] io_instBuffer_inst_1_bits_inst,
  input         io_instBuffer_inst_1_bits_tlb_invalid,
  input         io_instBuffer_info_inst0_is_in_delayslot,
  input         io_instBuffer_info_empty,
  input         io_instBuffer_info_almost_empty,
  output        io_instBuffer_inst0_is_jb,
  output [4:0]  io_regfile_0_src1_raddr,
  input  [31:0] io_regfile_0_src1_rdata,
  output [4:0]  io_regfile_0_src2_raddr,
  input  [31:0] io_regfile_0_src2_rdata,
  output [4:0]  io_regfile_1_src1_raddr,
  input  [31:0] io_regfile_1_src1_rdata,
  output [4:0]  io_regfile_1_src2_raddr,
  input  [31:0] io_regfile_1_src2_rdata,
  input         io_forward_0_exe_wen,
  input  [4:0]  io_forward_0_exe_waddr,
  input  [31:0] io_forward_0_exe_wdata,
  input         io_forward_0_exe_mem_ren,
  input         io_forward_0_mem_wen,
  input  [4:0]  io_forward_0_mem_waddr,
  input  [31:0] io_forward_0_mem_wdata,
  input         io_forward_1_exe_wen,
  input  [4:0]  io_forward_1_exe_waddr,
  input  [31:0] io_forward_1_exe_wdata,
  input         io_forward_1_exe_mem_ren,
  input         io_forward_1_mem_wen,
  input  [4:0]  io_forward_1_mem_waddr,
  input  [31:0] io_forward_1_mem_wdata,
  input         io_cp0_access_allowed,
  input         io_cp0_kernel_mode,
  input         io_cp0_intterupt_allowed,
  input  [7:0]  io_cp0_cause_ip,
  input  [7:0]  io_cp0_status_im,
  output        io_fetchUnit_branch,
  output [31:0] io_fetchUnit_target,
  output [31:0] io_bpu_pc,
  output [31:0] io_bpu_decoded_inst0_inst,
  input         io_bpu_inst_is_branch,
  input         io_bpu_pred_branch_flag,
  input  [31:0] io_bpu_branch_target,
  output [31:0] io_executeStage_inst0_pc,
  output [3:0]  io_executeStage_inst0_inst_info_fusel,
  output [6:0]  io_executeStage_inst0_inst_info_op,
  output        io_executeStage_inst0_inst_info_reg_wen,
  output [4:0]  io_executeStage_inst0_inst_info_reg_waddr,
  output [7:0]  io_executeStage_inst0_inst_info_cp0_addr,
  output [31:0] io_executeStage_inst0_inst_info_inst,
  output [31:0] io_executeStage_inst0_src_info_src1_data,
  output [31:0] io_executeStage_inst0_src_info_src2_data,
  output        io_executeStage_inst0_ex_flush_req,
  output        io_executeStage_inst0_ex_tlb_refill,
  output        io_executeStage_inst0_ex_eret,
  output [31:0] io_executeStage_inst0_ex_badvaddr,
  output        io_executeStage_inst0_ex_bd,
  output [4:0]  io_executeStage_inst0_ex_excode,
  output        io_executeStage_inst0_jb_info_jump_regiser_conflict,
  output        io_executeStage_inst0_jb_info_is_branch,
  output        io_executeStage_inst0_jb_info_pred_branch_flag,
  output [31:0] io_executeStage_inst0_jb_info_branch_target,
  output        io_executeStage_inst1_allow_to_go,
  output [31:0] io_executeStage_inst1_pc,
  output [3:0]  io_executeStage_inst1_inst_info_fusel,
  output [6:0]  io_executeStage_inst1_inst_info_op,
  output        io_executeStage_inst1_inst_info_reg_wen,
  output [4:0]  io_executeStage_inst1_inst_info_reg_waddr,
  output [31:0] io_executeStage_inst1_inst_info_inst,
  output [31:0] io_executeStage_inst1_src_info_src1_data,
  output [31:0] io_executeStage_inst1_src_info_src2_data,
  output        io_executeStage_inst1_ex_flush_req,
  output        io_executeStage_inst1_ex_tlb_refill,
  output        io_executeStage_inst1_ex_eret,
  output [31:0] io_executeStage_inst1_ex_badvaddr,
  output        io_executeStage_inst1_ex_bd,
  output [4:0]  io_executeStage_inst1_ex_excode,
  output        io_ctrl_inst0_src1_ren,
  output [4:0]  io_ctrl_inst0_src1_raddr,
  output        io_ctrl_inst0_src2_ren,
  output [4:0]  io_ctrl_inst0_src2_raddr,
  output        io_ctrl_branch_flag,
  input         io_ctrl_allow_to_go
);
  wire  Issue_io_allow_to_go; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_instBuffer_empty; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_instBuffer_almost_empty; // @[DecoderUnit.scala 70:27]
  wire [3:0] Issue_io_decodeInst_0_fusel; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_decodeInst_0_reg_wen; // @[DecoderUnit.scala 70:27]
  wire [4:0] Issue_io_decodeInst_0_reg_waddr; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_decodeInst_0_dual_issue; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_decodeInst_1_reg1_ren; // @[DecoderUnit.scala 70:27]
  wire [4:0] Issue_io_decodeInst_1_reg1_raddr; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_decodeInst_1_reg2_ren; // @[DecoderUnit.scala 70:27]
  wire [4:0] Issue_io_decodeInst_1_reg2_raddr; // @[DecoderUnit.scala 70:27]
  wire [3:0] Issue_io_decodeInst_1_fusel; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_decodeInst_1_dual_issue; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_execute_0_mem_ren; // @[DecoderUnit.scala 70:27]
  wire [4:0] Issue_io_execute_0_reg_waddr; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_execute_1_mem_ren; // @[DecoderUnit.scala 70:27]
  wire [4:0] Issue_io_execute_1_reg_waddr; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_inst1_is_in_delayslot; // @[DecoderUnit.scala 70:27]
  wire  Issue_io_inst1_allow_to_go; // @[DecoderUnit.scala 70:27]
  wire [31:0] decoder_0_io_in_inst; // @[DecoderUnit.scala 71:55]
  wire  decoder_0_io_out_inst_valid; // @[DecoderUnit.scala 71:55]
  wire  decoder_0_io_out_reg1_ren; // @[DecoderUnit.scala 71:55]
  wire [4:0] decoder_0_io_out_reg1_raddr; // @[DecoderUnit.scala 71:55]
  wire  decoder_0_io_out_reg2_ren; // @[DecoderUnit.scala 71:55]
  wire [4:0] decoder_0_io_out_reg2_raddr; // @[DecoderUnit.scala 71:55]
  wire [3:0] decoder_0_io_out_fusel; // @[DecoderUnit.scala 71:55]
  wire [6:0] decoder_0_io_out_op; // @[DecoderUnit.scala 71:55]
  wire  decoder_0_io_out_reg_wen; // @[DecoderUnit.scala 71:55]
  wire [4:0] decoder_0_io_out_reg_waddr; // @[DecoderUnit.scala 71:55]
  wire [31:0] decoder_0_io_out_imm32; // @[DecoderUnit.scala 71:55]
  wire [7:0] decoder_0_io_out_cp0_addr; // @[DecoderUnit.scala 71:55]
  wire  decoder_0_io_out_dual_issue; // @[DecoderUnit.scala 71:55]
  wire [31:0] decoder_0_io_out_inst; // @[DecoderUnit.scala 71:55]
  wire [31:0] decoder_1_io_in_inst; // @[DecoderUnit.scala 71:55]
  wire  decoder_1_io_out_inst_valid; // @[DecoderUnit.scala 71:55]
  wire  decoder_1_io_out_reg1_ren; // @[DecoderUnit.scala 71:55]
  wire [4:0] decoder_1_io_out_reg1_raddr; // @[DecoderUnit.scala 71:55]
  wire  decoder_1_io_out_reg2_ren; // @[DecoderUnit.scala 71:55]
  wire [4:0] decoder_1_io_out_reg2_raddr; // @[DecoderUnit.scala 71:55]
  wire [3:0] decoder_1_io_out_fusel; // @[DecoderUnit.scala 71:55]
  wire [6:0] decoder_1_io_out_op; // @[DecoderUnit.scala 71:55]
  wire  decoder_1_io_out_reg_wen; // @[DecoderUnit.scala 71:55]
  wire [4:0] decoder_1_io_out_reg_waddr; // @[DecoderUnit.scala 71:55]
  wire [31:0] decoder_1_io_out_imm32; // @[DecoderUnit.scala 71:55]
  wire [7:0] decoder_1_io_out_cp0_addr; // @[DecoderUnit.scala 71:55]
  wire  decoder_1_io_out_dual_issue; // @[DecoderUnit.scala 71:55]
  wire [31:0] decoder_1_io_out_inst; // @[DecoderUnit.scala 71:55]
  wire  JumpCtrl_io_in_allow_to_go; // @[DecoderUnit.scala 72:27]
  wire [31:0] JumpCtrl_io_in_pc; // @[DecoderUnit.scala 72:27]
  wire [4:0] JumpCtrl_io_in_decoded_inst0_reg1_raddr; // @[DecoderUnit.scala 72:27]
  wire [6:0] JumpCtrl_io_in_decoded_inst0_op; // @[DecoderUnit.scala 72:27]
  wire [31:0] JumpCtrl_io_in_decoded_inst0_inst; // @[DecoderUnit.scala 72:27]
  wire [31:0] JumpCtrl_io_in_reg1_data; // @[DecoderUnit.scala 72:27]
  wire  JumpCtrl_io_in_forward_0_exe_wen; // @[DecoderUnit.scala 72:27]
  wire [4:0] JumpCtrl_io_in_forward_0_exe_waddr; // @[DecoderUnit.scala 72:27]
  wire  JumpCtrl_io_in_forward_0_mem_wen; // @[DecoderUnit.scala 72:27]
  wire [4:0] JumpCtrl_io_in_forward_0_mem_waddr; // @[DecoderUnit.scala 72:27]
  wire  JumpCtrl_io_in_forward_1_exe_wen; // @[DecoderUnit.scala 72:27]
  wire [4:0] JumpCtrl_io_in_forward_1_exe_waddr; // @[DecoderUnit.scala 72:27]
  wire  JumpCtrl_io_in_forward_1_mem_wen; // @[DecoderUnit.scala 72:27]
  wire [4:0] JumpCtrl_io_in_forward_1_mem_waddr; // @[DecoderUnit.scala 72:27]
  wire  JumpCtrl_io_out_inst_is_jump; // @[DecoderUnit.scala 72:27]
  wire  JumpCtrl_io_out_jump_register; // @[DecoderUnit.scala 72:27]
  wire  JumpCtrl_io_out_jump_flag; // @[DecoderUnit.scala 72:27]
  wire [31:0] JumpCtrl_io_out_jump_target; // @[DecoderUnit.scala 72:27]
  wire  ForwardCtrl_io_in_forward_0_exe_wen; // @[DecoderUnit.scala 73:27]
  wire [4:0] ForwardCtrl_io_in_forward_0_exe_waddr; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_in_forward_0_exe_wdata; // @[DecoderUnit.scala 73:27]
  wire  ForwardCtrl_io_in_forward_0_exe_mem_ren; // @[DecoderUnit.scala 73:27]
  wire  ForwardCtrl_io_in_forward_0_mem_wen; // @[DecoderUnit.scala 73:27]
  wire [4:0] ForwardCtrl_io_in_forward_0_mem_waddr; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_in_forward_0_mem_wdata; // @[DecoderUnit.scala 73:27]
  wire  ForwardCtrl_io_in_forward_1_exe_wen; // @[DecoderUnit.scala 73:27]
  wire [4:0] ForwardCtrl_io_in_forward_1_exe_waddr; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_in_forward_1_exe_wdata; // @[DecoderUnit.scala 73:27]
  wire  ForwardCtrl_io_in_forward_1_exe_mem_ren; // @[DecoderUnit.scala 73:27]
  wire  ForwardCtrl_io_in_forward_1_mem_wen; // @[DecoderUnit.scala 73:27]
  wire [4:0] ForwardCtrl_io_in_forward_1_mem_waddr; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_in_forward_1_mem_wdata; // @[DecoderUnit.scala 73:27]
  wire [4:0] ForwardCtrl_io_in_regfile_0_src1_raddr; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_in_regfile_0_src1_rdata; // @[DecoderUnit.scala 73:27]
  wire [4:0] ForwardCtrl_io_in_regfile_0_src2_raddr; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_in_regfile_0_src2_rdata; // @[DecoderUnit.scala 73:27]
  wire [4:0] ForwardCtrl_io_in_regfile_1_src1_raddr; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_in_regfile_1_src1_rdata; // @[DecoderUnit.scala 73:27]
  wire [4:0] ForwardCtrl_io_in_regfile_1_src2_raddr; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_in_regfile_1_src2_rdata; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_out_inst_0_src1_rdata; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_out_inst_0_src2_rdata; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_out_inst_1_src1_rdata; // @[DecoderUnit.scala 73:27]
  wire [31:0] ForwardCtrl_io_out_inst_1_src2_rdata; // @[DecoderUnit.scala 73:27]
  wire [7:0] _interrupt_T = io_cp0_cause_ip & io_cp0_status_im; // @[DecoderUnit.scala 117:66]
  wire  interrupt = io_cp0_intterupt_allowed & |_interrupt_T & ~io_instBuffer_info_empty; // @[DecoderUnit.scala 117:92]
  wire  _io_executeStage_inst0_ex_flush_req_T_1 = io_executeStage_inst0_ex_excode != 5'h0 |
    io_executeStage_inst0_ex_tlb_refill; // @[DecoderUnit.scala 139:47]
  wire  _io_executeStage_inst0_ex_excode_T_4 = ~io_cp0_kernel_mode; // @[DecoderUnit.scala 151:43]
  wire  _io_executeStage_inst0_ex_excode_T_6 = |io_instBuffer_inst_0_bits_pc[1:0] | io_instBuffer_inst_0_bits_pc[31] & ~
    io_cp0_kernel_mode; // @[DecoderUnit.scala 151:26]
  wire  _io_executeStage_inst0_ex_excode_T_7 = decoder_0_io_out_inst_valid; // @[DecoderUnit.scala 152:32]
  wire  _io_executeStage_inst0_ex_excode_T_8 = decoder_0_io_out_op == 7'h44; // @[DecoderUnit.scala 153:24]
  wire  _io_executeStage_inst0_ex_excode_T_9 = decoder_0_io_out_op == 7'h45; // @[DecoderUnit.scala 154:24]
  wire  _io_executeStage_inst0_ex_excode_T_10 = ~io_cp0_access_allowed; // @[DecoderUnit.scala 155:8]
  wire [4:0] _io_executeStage_inst0_ex_excode_T_11 = _io_executeStage_inst0_ex_excode_T_10 ? 5'ha : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_executeStage_inst0_ex_excode_T_12 = _io_executeStage_inst0_ex_excode_T_9 ? 5'h8 :
    _io_executeStage_inst0_ex_excode_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_executeStage_inst0_ex_excode_T_13 = _io_executeStage_inst0_ex_excode_T_8 ? 5'h7 :
    _io_executeStage_inst0_ex_excode_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_executeStage_inst0_ex_excode_T_14 = _io_executeStage_inst0_ex_excode_T_7 ? 5'h9 :
    _io_executeStage_inst0_ex_excode_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_executeStage_inst0_ex_excode_T_15 = _io_executeStage_inst0_ex_excode_T_6 ? 5'h5 :
    _io_executeStage_inst0_ex_excode_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_executeStage_inst0_ex_excode_T_16 = io_instBuffer_inst_0_bits_tlb_invalid ? 5'h3 :
    _io_executeStage_inst0_ex_excode_T_15; // @[Mux.scala 101:16]
  wire  _io_executeStage_inst1_ex_excode_T_6 = |io_instBuffer_inst_1_bits_pc[1:0] | io_instBuffer_inst_1_bits_pc[31] &
    _io_executeStage_inst0_ex_excode_T_4; // @[DecoderUnit.scala 185:26]
  wire  _io_executeStage_inst1_ex_excode_T_7 = decoder_1_io_out_inst_valid; // @[DecoderUnit.scala 186:32]
  wire  _io_executeStage_inst1_ex_excode_T_8 = decoder_1_io_out_op == 7'h44; // @[DecoderUnit.scala 187:24]
  wire  _io_executeStage_inst1_ex_excode_T_9 = decoder_1_io_out_op == 7'h45; // @[DecoderUnit.scala 188:24]
  wire [4:0] _io_executeStage_inst1_ex_excode_T_12 = _io_executeStage_inst1_ex_excode_T_9 ? 5'h8 :
    _io_executeStage_inst0_ex_excode_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_executeStage_inst1_ex_excode_T_13 = _io_executeStage_inst1_ex_excode_T_8 ? 5'h7 :
    _io_executeStage_inst1_ex_excode_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_executeStage_inst1_ex_excode_T_14 = _io_executeStage_inst1_ex_excode_T_7 ? 5'h9 :
    _io_executeStage_inst1_ex_excode_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_executeStage_inst1_ex_excode_T_15 = _io_executeStage_inst1_ex_excode_T_6 ? 5'h5 :
    _io_executeStage_inst1_ex_excode_T_14; // @[Mux.scala 101:16]
  Issue Issue ( // @[DecoderUnit.scala 70:27]
    .io_allow_to_go(Issue_io_allow_to_go),
    .io_instBuffer_empty(Issue_io_instBuffer_empty),
    .io_instBuffer_almost_empty(Issue_io_instBuffer_almost_empty),
    .io_decodeInst_0_fusel(Issue_io_decodeInst_0_fusel),
    .io_decodeInst_0_reg_wen(Issue_io_decodeInst_0_reg_wen),
    .io_decodeInst_0_reg_waddr(Issue_io_decodeInst_0_reg_waddr),
    .io_decodeInst_0_dual_issue(Issue_io_decodeInst_0_dual_issue),
    .io_decodeInst_1_reg1_ren(Issue_io_decodeInst_1_reg1_ren),
    .io_decodeInst_1_reg1_raddr(Issue_io_decodeInst_1_reg1_raddr),
    .io_decodeInst_1_reg2_ren(Issue_io_decodeInst_1_reg2_ren),
    .io_decodeInst_1_reg2_raddr(Issue_io_decodeInst_1_reg2_raddr),
    .io_decodeInst_1_fusel(Issue_io_decodeInst_1_fusel),
    .io_decodeInst_1_dual_issue(Issue_io_decodeInst_1_dual_issue),
    .io_execute_0_mem_ren(Issue_io_execute_0_mem_ren),
    .io_execute_0_reg_waddr(Issue_io_execute_0_reg_waddr),
    .io_execute_1_mem_ren(Issue_io_execute_1_mem_ren),
    .io_execute_1_reg_waddr(Issue_io_execute_1_reg_waddr),
    .io_inst1_is_in_delayslot(Issue_io_inst1_is_in_delayslot),
    .io_inst1_allow_to_go(Issue_io_inst1_allow_to_go)
  );
  Decoder decoder_0 ( // @[DecoderUnit.scala 71:55]
    .io_in_inst(decoder_0_io_in_inst),
    .io_out_inst_valid(decoder_0_io_out_inst_valid),
    .io_out_reg1_ren(decoder_0_io_out_reg1_ren),
    .io_out_reg1_raddr(decoder_0_io_out_reg1_raddr),
    .io_out_reg2_ren(decoder_0_io_out_reg2_ren),
    .io_out_reg2_raddr(decoder_0_io_out_reg2_raddr),
    .io_out_fusel(decoder_0_io_out_fusel),
    .io_out_op(decoder_0_io_out_op),
    .io_out_reg_wen(decoder_0_io_out_reg_wen),
    .io_out_reg_waddr(decoder_0_io_out_reg_waddr),
    .io_out_imm32(decoder_0_io_out_imm32),
    .io_out_cp0_addr(decoder_0_io_out_cp0_addr),
    .io_out_dual_issue(decoder_0_io_out_dual_issue),
    .io_out_inst(decoder_0_io_out_inst)
  );
  Decoder decoder_1 ( // @[DecoderUnit.scala 71:55]
    .io_in_inst(decoder_1_io_in_inst),
    .io_out_inst_valid(decoder_1_io_out_inst_valid),
    .io_out_reg1_ren(decoder_1_io_out_reg1_ren),
    .io_out_reg1_raddr(decoder_1_io_out_reg1_raddr),
    .io_out_reg2_ren(decoder_1_io_out_reg2_ren),
    .io_out_reg2_raddr(decoder_1_io_out_reg2_raddr),
    .io_out_fusel(decoder_1_io_out_fusel),
    .io_out_op(decoder_1_io_out_op),
    .io_out_reg_wen(decoder_1_io_out_reg_wen),
    .io_out_reg_waddr(decoder_1_io_out_reg_waddr),
    .io_out_imm32(decoder_1_io_out_imm32),
    .io_out_cp0_addr(decoder_1_io_out_cp0_addr),
    .io_out_dual_issue(decoder_1_io_out_dual_issue),
    .io_out_inst(decoder_1_io_out_inst)
  );
  JumpCtrl JumpCtrl ( // @[DecoderUnit.scala 72:27]
    .io_in_allow_to_go(JumpCtrl_io_in_allow_to_go),
    .io_in_pc(JumpCtrl_io_in_pc),
    .io_in_decoded_inst0_reg1_raddr(JumpCtrl_io_in_decoded_inst0_reg1_raddr),
    .io_in_decoded_inst0_op(JumpCtrl_io_in_decoded_inst0_op),
    .io_in_decoded_inst0_inst(JumpCtrl_io_in_decoded_inst0_inst),
    .io_in_reg1_data(JumpCtrl_io_in_reg1_data),
    .io_in_forward_0_exe_wen(JumpCtrl_io_in_forward_0_exe_wen),
    .io_in_forward_0_exe_waddr(JumpCtrl_io_in_forward_0_exe_waddr),
    .io_in_forward_0_mem_wen(JumpCtrl_io_in_forward_0_mem_wen),
    .io_in_forward_0_mem_waddr(JumpCtrl_io_in_forward_0_mem_waddr),
    .io_in_forward_1_exe_wen(JumpCtrl_io_in_forward_1_exe_wen),
    .io_in_forward_1_exe_waddr(JumpCtrl_io_in_forward_1_exe_waddr),
    .io_in_forward_1_mem_wen(JumpCtrl_io_in_forward_1_mem_wen),
    .io_in_forward_1_mem_waddr(JumpCtrl_io_in_forward_1_mem_waddr),
    .io_out_inst_is_jump(JumpCtrl_io_out_inst_is_jump),
    .io_out_jump_register(JumpCtrl_io_out_jump_register),
    .io_out_jump_flag(JumpCtrl_io_out_jump_flag),
    .io_out_jump_target(JumpCtrl_io_out_jump_target)
  );
  ForwardCtrl ForwardCtrl ( // @[DecoderUnit.scala 73:27]
    .io_in_forward_0_exe_wen(ForwardCtrl_io_in_forward_0_exe_wen),
    .io_in_forward_0_exe_waddr(ForwardCtrl_io_in_forward_0_exe_waddr),
    .io_in_forward_0_exe_wdata(ForwardCtrl_io_in_forward_0_exe_wdata),
    .io_in_forward_0_exe_mem_ren(ForwardCtrl_io_in_forward_0_exe_mem_ren),
    .io_in_forward_0_mem_wen(ForwardCtrl_io_in_forward_0_mem_wen),
    .io_in_forward_0_mem_waddr(ForwardCtrl_io_in_forward_0_mem_waddr),
    .io_in_forward_0_mem_wdata(ForwardCtrl_io_in_forward_0_mem_wdata),
    .io_in_forward_1_exe_wen(ForwardCtrl_io_in_forward_1_exe_wen),
    .io_in_forward_1_exe_waddr(ForwardCtrl_io_in_forward_1_exe_waddr),
    .io_in_forward_1_exe_wdata(ForwardCtrl_io_in_forward_1_exe_wdata),
    .io_in_forward_1_exe_mem_ren(ForwardCtrl_io_in_forward_1_exe_mem_ren),
    .io_in_forward_1_mem_wen(ForwardCtrl_io_in_forward_1_mem_wen),
    .io_in_forward_1_mem_waddr(ForwardCtrl_io_in_forward_1_mem_waddr),
    .io_in_forward_1_mem_wdata(ForwardCtrl_io_in_forward_1_mem_wdata),
    .io_in_regfile_0_src1_raddr(ForwardCtrl_io_in_regfile_0_src1_raddr),
    .io_in_regfile_0_src1_rdata(ForwardCtrl_io_in_regfile_0_src1_rdata),
    .io_in_regfile_0_src2_raddr(ForwardCtrl_io_in_regfile_0_src2_raddr),
    .io_in_regfile_0_src2_rdata(ForwardCtrl_io_in_regfile_0_src2_rdata),
    .io_in_regfile_1_src1_raddr(ForwardCtrl_io_in_regfile_1_src1_raddr),
    .io_in_regfile_1_src1_rdata(ForwardCtrl_io_in_regfile_1_src1_rdata),
    .io_in_regfile_1_src2_raddr(ForwardCtrl_io_in_regfile_1_src2_raddr),
    .io_in_regfile_1_src2_rdata(ForwardCtrl_io_in_regfile_1_src2_rdata),
    .io_out_inst_0_src1_rdata(ForwardCtrl_io_out_inst_0_src1_rdata),
    .io_out_inst_0_src2_rdata(ForwardCtrl_io_out_inst_0_src2_rdata),
    .io_out_inst_1_src1_rdata(ForwardCtrl_io_out_inst_1_src1_rdata),
    .io_out_inst_1_src2_rdata(ForwardCtrl_io_out_inst_1_src2_rdata)
  );
  assign io_instBuffer_inst_0_ready = io_ctrl_allow_to_go; // @[DecoderUnit.scala 98:31]
  assign io_instBuffer_inst_1_ready = Issue_io_inst1_allow_to_go; // @[DecoderUnit.scala 99:31]
  assign io_instBuffer_inst0_is_jb = JumpCtrl_io_out_inst_is_jump | io_bpu_inst_is_branch; // @[DecoderUnit.scala 92:49]
  assign io_regfile_0_src1_raddr = decoder_0_io_out_reg1_raddr; // @[DecoderUnit.scala 75:28]
  assign io_regfile_0_src2_raddr = decoder_0_io_out_reg2_raddr; // @[DecoderUnit.scala 76:28]
  assign io_regfile_1_src1_raddr = decoder_1_io_out_reg1_raddr; // @[DecoderUnit.scala 77:28]
  assign io_regfile_1_src2_raddr = decoder_1_io_out_reg2_raddr; // @[DecoderUnit.scala 78:28]
  assign io_fetchUnit_branch = JumpCtrl_io_out_jump_flag | io_bpu_pred_branch_flag; // @[DecoderUnit.scala 93:46]
  assign io_fetchUnit_target = io_bpu_pred_branch_flag ? io_bpu_branch_target : JumpCtrl_io_out_jump_target; // @[DecoderUnit.scala 96:29]
  assign io_bpu_pc = io_instBuffer_inst_0_bits_pc; // @[DecoderUnit.scala 103:25]
  assign io_bpu_decoded_inst0_inst = decoder_0_io_out_inst; // @[DecoderUnit.scala 104:25]
  assign io_executeStage_inst0_pc = io_instBuffer_inst_0_bits_pc; // @[DecoderUnit.scala 126:35]
  assign io_executeStage_inst0_inst_info_fusel = decoder_0_io_out_fusel; // @[DecoderUnit.scala 127:35]
  assign io_executeStage_inst0_inst_info_op = decoder_0_io_out_op; // @[DecoderUnit.scala 127:35]
  assign io_executeStage_inst0_inst_info_reg_wen = decoder_0_io_out_reg_wen; // @[DecoderUnit.scala 127:35]
  assign io_executeStage_inst0_inst_info_reg_waddr = decoder_0_io_out_reg_waddr; // @[DecoderUnit.scala 127:35]
  assign io_executeStage_inst0_inst_info_cp0_addr = decoder_0_io_out_cp0_addr; // @[DecoderUnit.scala 127:35]
  assign io_executeStage_inst0_inst_info_inst = decoder_0_io_out_inst; // @[DecoderUnit.scala 127:35]
  assign io_executeStage_inst0_src_info_src1_data = decoder_0_io_out_reg1_ren ? ForwardCtrl_io_out_inst_0_src1_rdata :
    decoder_0_io_out_imm32; // @[DecoderUnit.scala 128:50]
  assign io_executeStage_inst0_src_info_src2_data = decoder_0_io_out_reg2_ren ? ForwardCtrl_io_out_inst_0_src2_rdata :
    decoder_0_io_out_imm32; // @[DecoderUnit.scala 133:50]
  assign io_executeStage_inst0_ex_flush_req = _io_executeStage_inst0_ex_flush_req_T_1 | io_executeStage_inst0_ex_eret; // @[DecoderUnit.scala 140:43]
  assign io_executeStage_inst0_ex_tlb_refill = 1'h0; // @[DecoderUnit.scala 142:39]
  assign io_executeStage_inst0_ex_eret = decoder_0_io_out_op == 7'h46; // @[DecoderUnit.scala 143:58]
  assign io_executeStage_inst0_ex_badvaddr = io_instBuffer_inst_0_bits_pc; // @[DecoderUnit.scala 144:39]
  assign io_executeStage_inst0_ex_bd = io_instBuffer_info_inst0_is_in_delayslot; // @[DecoderUnit.scala 145:39]
  assign io_executeStage_inst0_ex_excode = interrupt ? 5'h1 : _io_executeStage_inst0_ex_excode_T_16; // @[Mux.scala 101:16]
  assign io_executeStage_inst0_jb_info_jump_regiser_conflict = JumpCtrl_io_out_jump_register; // @[DecoderUnit.scala 158:55]
  assign io_executeStage_inst0_jb_info_is_branch = io_bpu_inst_is_branch; // @[DecoderUnit.scala 159:55]
  assign io_executeStage_inst0_jb_info_pred_branch_flag = io_bpu_pred_branch_flag; // @[DecoderUnit.scala 160:55]
  assign io_executeStage_inst0_jb_info_branch_target = io_bpu_branch_target; // @[DecoderUnit.scala 161:55]
  assign io_executeStage_inst1_allow_to_go = Issue_io_inst1_allow_to_go; // @[DecoderUnit.scala 163:37]
  assign io_executeStage_inst1_pc = io_instBuffer_inst_1_bits_pc; // @[DecoderUnit.scala 164:37]
  assign io_executeStage_inst1_inst_info_fusel = decoder_1_io_out_fusel; // @[DecoderUnit.scala 165:37]
  assign io_executeStage_inst1_inst_info_op = decoder_1_io_out_op; // @[DecoderUnit.scala 165:37]
  assign io_executeStage_inst1_inst_info_reg_wen = decoder_1_io_out_reg_wen; // @[DecoderUnit.scala 165:37]
  assign io_executeStage_inst1_inst_info_reg_waddr = decoder_1_io_out_reg_waddr; // @[DecoderUnit.scala 165:37]
  assign io_executeStage_inst1_inst_info_inst = decoder_1_io_out_inst; // @[DecoderUnit.scala 165:37]
  assign io_executeStage_inst1_src_info_src1_data = decoder_1_io_out_reg1_ren ? ForwardCtrl_io_out_inst_1_src1_rdata :
    decoder_1_io_out_imm32; // @[DecoderUnit.scala 166:50]
  assign io_executeStage_inst1_src_info_src2_data = decoder_1_io_out_reg2_ren ? ForwardCtrl_io_out_inst_1_src2_rdata :
    decoder_1_io_out_imm32; // @[DecoderUnit.scala 171:50]
  assign io_executeStage_inst1_ex_flush_req = io_executeStage_inst1_ex_excode != 5'h0 |
    io_executeStage_inst1_ex_tlb_refill; // @[DecoderUnit.scala 176:83]
  assign io_executeStage_inst1_ex_tlb_refill = 1'h0; // @[DecoderUnit.scala 177:39]
  assign io_executeStage_inst1_ex_eret = decoder_1_io_out_op == 7'h46; // @[DecoderUnit.scala 178:58]
  assign io_executeStage_inst1_ex_badvaddr = io_instBuffer_inst_1_bits_pc; // @[DecoderUnit.scala 179:39]
  assign io_executeStage_inst1_ex_bd = Issue_io_inst1_is_in_delayslot; // @[DecoderUnit.scala 180:39]
  assign io_executeStage_inst1_ex_excode = io_instBuffer_inst_1_bits_tlb_invalid ? 5'h3 :
    _io_executeStage_inst1_ex_excode_T_15; // @[Mux.scala 101:16]
  assign io_ctrl_inst0_src1_ren = decoder_0_io_out_reg1_ren; // @[DecoderUnit.scala 106:28]
  assign io_ctrl_inst0_src1_raddr = decoder_0_io_out_reg1_raddr; // @[DecoderUnit.scala 107:28]
  assign io_ctrl_inst0_src2_ren = decoder_0_io_out_reg2_ren; // @[DecoderUnit.scala 108:28]
  assign io_ctrl_inst0_src2_raddr = decoder_0_io_out_reg2_raddr; // @[DecoderUnit.scala 109:28]
  assign io_ctrl_branch_flag = JumpCtrl_io_out_jump_flag | io_bpu_pred_branch_flag; // @[DecoderUnit.scala 93:46]
  assign Issue_io_allow_to_go = io_ctrl_allow_to_go; // @[DecoderUnit.scala 83:21]
  assign Issue_io_instBuffer_empty = io_instBuffer_info_empty; // @[DecoderUnit.scala 84:21]
  assign Issue_io_instBuffer_almost_empty = io_instBuffer_info_almost_empty; // @[DecoderUnit.scala 84:21]
  assign Issue_io_decodeInst_0_fusel = decoder_0_io_out_fusel; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_0_reg_wen = decoder_0_io_out_reg_wen; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_0_reg_waddr = decoder_0_io_out_reg_waddr; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_0_dual_issue = decoder_0_io_out_dual_issue; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_1_reg1_ren = decoder_1_io_out_reg1_ren; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_1_reg1_raddr = decoder_1_io_out_reg1_raddr; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_1_reg2_ren = decoder_1_io_out_reg2_ren; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_1_reg2_raddr = decoder_1_io_out_reg2_raddr; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_1_fusel = decoder_1_io_out_fusel; // @[DecoderUnit.scala 121:32]
  assign Issue_io_decodeInst_1_dual_issue = decoder_1_io_out_dual_issue; // @[DecoderUnit.scala 121:32]
  assign Issue_io_execute_0_mem_ren = io_forward_0_exe_mem_ren; // @[DecoderUnit.scala 122:32]
  assign Issue_io_execute_0_reg_waddr = io_forward_0_exe_waddr; // @[DecoderUnit.scala 123:32]
  assign Issue_io_execute_1_mem_ren = io_forward_1_exe_mem_ren; // @[DecoderUnit.scala 122:32]
  assign Issue_io_execute_1_reg_waddr = io_forward_1_exe_waddr; // @[DecoderUnit.scala 123:32]
  assign decoder_0_io_in_inst = io_instBuffer_inst_0_bits_inst; // @[DecoderUnit.scala 120:32]
  assign decoder_1_io_in_inst = io_instBuffer_inst_1_bits_inst; // @[DecoderUnit.scala 120:32]
  assign JumpCtrl_io_in_allow_to_go = io_ctrl_allow_to_go; // @[DecoderUnit.scala 86:29]
  assign JumpCtrl_io_in_pc = io_instBuffer_inst_0_bits_pc; // @[DecoderUnit.scala 89:29]
  assign JumpCtrl_io_in_decoded_inst0_reg1_raddr = decoder_0_io_out_reg1_raddr; // @[DecoderUnit.scala 87:29]
  assign JumpCtrl_io_in_decoded_inst0_op = decoder_0_io_out_op; // @[DecoderUnit.scala 87:29]
  assign JumpCtrl_io_in_decoded_inst0_inst = decoder_0_io_out_inst; // @[DecoderUnit.scala 87:29]
  assign JumpCtrl_io_in_reg1_data = io_regfile_0_src1_rdata; // @[DecoderUnit.scala 90:29]
  assign JumpCtrl_io_in_forward_0_exe_wen = io_forward_0_exe_wen; // @[DecoderUnit.scala 88:29]
  assign JumpCtrl_io_in_forward_0_exe_waddr = io_forward_0_exe_waddr; // @[DecoderUnit.scala 88:29]
  assign JumpCtrl_io_in_forward_0_mem_wen = io_forward_0_mem_wen; // @[DecoderUnit.scala 88:29]
  assign JumpCtrl_io_in_forward_0_mem_waddr = io_forward_0_mem_waddr; // @[DecoderUnit.scala 88:29]
  assign JumpCtrl_io_in_forward_1_exe_wen = io_forward_1_exe_wen; // @[DecoderUnit.scala 88:29]
  assign JumpCtrl_io_in_forward_1_exe_waddr = io_forward_1_exe_waddr; // @[DecoderUnit.scala 88:29]
  assign JumpCtrl_io_in_forward_1_mem_wen = io_forward_1_mem_wen; // @[DecoderUnit.scala 88:29]
  assign JumpCtrl_io_in_forward_1_mem_waddr = io_forward_1_mem_waddr; // @[DecoderUnit.scala 88:29]
  assign ForwardCtrl_io_in_forward_0_exe_wen = io_forward_0_exe_wen; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_0_exe_waddr = io_forward_0_exe_waddr; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_0_exe_wdata = io_forward_0_exe_wdata; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_0_exe_mem_ren = io_forward_0_exe_mem_ren; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_0_mem_wen = io_forward_0_mem_wen; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_0_mem_waddr = io_forward_0_mem_waddr; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_0_mem_wdata = io_forward_0_mem_wdata; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_1_exe_wen = io_forward_1_exe_wen; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_1_exe_waddr = io_forward_1_exe_waddr; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_1_exe_wdata = io_forward_1_exe_wdata; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_1_exe_mem_ren = io_forward_1_exe_mem_ren; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_1_mem_wen = io_forward_1_mem_wen; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_1_mem_waddr = io_forward_1_mem_waddr; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_forward_1_mem_wdata = io_forward_1_mem_wdata; // @[DecoderUnit.scala 80:26]
  assign ForwardCtrl_io_in_regfile_0_src1_raddr = io_regfile_0_src1_raddr; // @[DecoderUnit.scala 81:26]
  assign ForwardCtrl_io_in_regfile_0_src1_rdata = io_regfile_0_src1_rdata; // @[DecoderUnit.scala 81:26]
  assign ForwardCtrl_io_in_regfile_0_src2_raddr = io_regfile_0_src2_raddr; // @[DecoderUnit.scala 81:26]
  assign ForwardCtrl_io_in_regfile_0_src2_rdata = io_regfile_0_src2_rdata; // @[DecoderUnit.scala 81:26]
  assign ForwardCtrl_io_in_regfile_1_src1_raddr = io_regfile_1_src1_raddr; // @[DecoderUnit.scala 81:26]
  assign ForwardCtrl_io_in_regfile_1_src1_rdata = io_regfile_1_src1_rdata; // @[DecoderUnit.scala 81:26]
  assign ForwardCtrl_io_in_regfile_1_src2_raddr = io_regfile_1_src2_raddr; // @[DecoderUnit.scala 81:26]
  assign ForwardCtrl_io_in_regfile_1_src2_rdata = io_regfile_1_src2_rdata; // @[DecoderUnit.scala 81:26]
endmodule
module ARegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_read_0_src1_raddr,
  output [31:0] io_read_0_src1_rdata,
  input  [4:0]  io_read_0_src2_raddr,
  output [31:0] io_read_0_src2_rdata,
  input  [4:0]  io_read_1_src1_raddr,
  output [31:0] io_read_1_src1_rdata,
  input  [4:0]  io_read_1_src2_raddr,
  output [31:0] io_read_1_src2_rdata,
  input         io_write_0_wen,
  input  [4:0]  io_write_0_waddr,
  input  [31:0] io_write_0_wdata,
  input         io_write_1_wen,
  input  [4:0]  io_write_1_waddr,
  input  [31:0] io_write_1_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[ARegfile.scala 32:21]
  reg [31:0] regs_1; // @[ARegfile.scala 32:21]
  reg [31:0] regs_2; // @[ARegfile.scala 32:21]
  reg [31:0] regs_3; // @[ARegfile.scala 32:21]
  reg [31:0] regs_4; // @[ARegfile.scala 32:21]
  reg [31:0] regs_5; // @[ARegfile.scala 32:21]
  reg [31:0] regs_6; // @[ARegfile.scala 32:21]
  reg [31:0] regs_7; // @[ARegfile.scala 32:21]
  reg [31:0] regs_8; // @[ARegfile.scala 32:21]
  reg [31:0] regs_9; // @[ARegfile.scala 32:21]
  reg [31:0] regs_10; // @[ARegfile.scala 32:21]
  reg [31:0] regs_11; // @[ARegfile.scala 32:21]
  reg [31:0] regs_12; // @[ARegfile.scala 32:21]
  reg [31:0] regs_13; // @[ARegfile.scala 32:21]
  reg [31:0] regs_14; // @[ARegfile.scala 32:21]
  reg [31:0] regs_15; // @[ARegfile.scala 32:21]
  reg [31:0] regs_16; // @[ARegfile.scala 32:21]
  reg [31:0] regs_17; // @[ARegfile.scala 32:21]
  reg [31:0] regs_18; // @[ARegfile.scala 32:21]
  reg [31:0] regs_19; // @[ARegfile.scala 32:21]
  reg [31:0] regs_20; // @[ARegfile.scala 32:21]
  reg [31:0] regs_21; // @[ARegfile.scala 32:21]
  reg [31:0] regs_22; // @[ARegfile.scala 32:21]
  reg [31:0] regs_23; // @[ARegfile.scala 32:21]
  reg [31:0] regs_24; // @[ARegfile.scala 32:21]
  reg [31:0] regs_25; // @[ARegfile.scala 32:21]
  reg [31:0] regs_26; // @[ARegfile.scala 32:21]
  reg [31:0] regs_27; // @[ARegfile.scala 32:21]
  reg [31:0] regs_28; // @[ARegfile.scala 32:21]
  reg [31:0] regs_29; // @[ARegfile.scala 32:21]
  reg [31:0] regs_30; // @[ARegfile.scala 32:21]
  reg [31:0] regs_31; // @[ARegfile.scala 32:21]
  wire [31:0] _GEN_0 = 5'h0 == io_write_0_waddr ? io_write_0_wdata : regs_0; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_1 = 5'h1 == io_write_0_waddr ? io_write_0_wdata : regs_1; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_2 = 5'h2 == io_write_0_waddr ? io_write_0_wdata : regs_2; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_3 = 5'h3 == io_write_0_waddr ? io_write_0_wdata : regs_3; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_4 = 5'h4 == io_write_0_waddr ? io_write_0_wdata : regs_4; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_5 = 5'h5 == io_write_0_waddr ? io_write_0_wdata : regs_5; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_6 = 5'h6 == io_write_0_waddr ? io_write_0_wdata : regs_6; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_7 = 5'h7 == io_write_0_waddr ? io_write_0_wdata : regs_7; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_8 = 5'h8 == io_write_0_waddr ? io_write_0_wdata : regs_8; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_9 = 5'h9 == io_write_0_waddr ? io_write_0_wdata : regs_9; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_10 = 5'ha == io_write_0_waddr ? io_write_0_wdata : regs_10; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_11 = 5'hb == io_write_0_waddr ? io_write_0_wdata : regs_11; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_12 = 5'hc == io_write_0_waddr ? io_write_0_wdata : regs_12; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_13 = 5'hd == io_write_0_waddr ? io_write_0_wdata : regs_13; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_14 = 5'he == io_write_0_waddr ? io_write_0_wdata : regs_14; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_15 = 5'hf == io_write_0_waddr ? io_write_0_wdata : regs_15; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_16 = 5'h10 == io_write_0_waddr ? io_write_0_wdata : regs_16; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_17 = 5'h11 == io_write_0_waddr ? io_write_0_wdata : regs_17; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_18 = 5'h12 == io_write_0_waddr ? io_write_0_wdata : regs_18; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_19 = 5'h13 == io_write_0_waddr ? io_write_0_wdata : regs_19; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_20 = 5'h14 == io_write_0_waddr ? io_write_0_wdata : regs_20; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_21 = 5'h15 == io_write_0_waddr ? io_write_0_wdata : regs_21; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_22 = 5'h16 == io_write_0_waddr ? io_write_0_wdata : regs_22; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_23 = 5'h17 == io_write_0_waddr ? io_write_0_wdata : regs_23; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_24 = 5'h18 == io_write_0_waddr ? io_write_0_wdata : regs_24; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_25 = 5'h19 == io_write_0_waddr ? io_write_0_wdata : regs_25; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_26 = 5'h1a == io_write_0_waddr ? io_write_0_wdata : regs_26; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_27 = 5'h1b == io_write_0_waddr ? io_write_0_wdata : regs_27; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_28 = 5'h1c == io_write_0_waddr ? io_write_0_wdata : regs_28; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_29 = 5'h1d == io_write_0_waddr ? io_write_0_wdata : regs_29; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_30 = 5'h1e == io_write_0_waddr ? io_write_0_wdata : regs_30; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_31 = 5'h1f == io_write_0_waddr ? io_write_0_wdata : regs_31; // @[ARegfile.scala 32:21 37:{31,31}]
  wire [31:0] _GEN_32 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_0 : regs_0; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_33 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_1 : regs_1; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_34 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_2 : regs_2; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_35 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_3 : regs_3; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_36 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_4 : regs_4; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_37 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_5 : regs_5; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_38 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_6 : regs_6; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_39 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_7 : regs_7; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_40 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_8 : regs_8; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_41 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_9 : regs_9; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_42 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_10 : regs_10; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_43 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_11 : regs_11; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_44 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_12 : regs_12; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_45 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_13 : regs_13; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_46 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_14 : regs_14; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_47 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_15 : regs_15; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_48 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_16 : regs_16; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_49 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_17 : regs_17; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_50 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_18 : regs_18; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_51 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_19 : regs_19; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_52 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_20 : regs_20; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_53 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_21 : regs_21; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_54 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_22 : regs_22; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_55 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_23 : regs_23; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_56 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_24 : regs_24; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_57 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_25 : regs_25; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_58 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_26 : regs_26; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_59 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_27 : regs_27; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_60 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_28 : regs_28; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_61 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_29 : regs_29; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_62 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_30 : regs_30; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_63 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_31 : regs_31; // @[ARegfile.scala 32:21 36:56]
  wire [31:0] _GEN_129 = 5'h1 == io_read_0_src1_raddr ? regs_1 : regs_0; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_130 = 5'h2 == io_read_0_src1_raddr ? regs_2 : _GEN_129; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_131 = 5'h3 == io_read_0_src1_raddr ? regs_3 : _GEN_130; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_132 = 5'h4 == io_read_0_src1_raddr ? regs_4 : _GEN_131; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_133 = 5'h5 == io_read_0_src1_raddr ? regs_5 : _GEN_132; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_134 = 5'h6 == io_read_0_src1_raddr ? regs_6 : _GEN_133; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_135 = 5'h7 == io_read_0_src1_raddr ? regs_7 : _GEN_134; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_136 = 5'h8 == io_read_0_src1_raddr ? regs_8 : _GEN_135; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_137 = 5'h9 == io_read_0_src1_raddr ? regs_9 : _GEN_136; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_138 = 5'ha == io_read_0_src1_raddr ? regs_10 : _GEN_137; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_139 = 5'hb == io_read_0_src1_raddr ? regs_11 : _GEN_138; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_140 = 5'hc == io_read_0_src1_raddr ? regs_12 : _GEN_139; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_141 = 5'hd == io_read_0_src1_raddr ? regs_13 : _GEN_140; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_142 = 5'he == io_read_0_src1_raddr ? regs_14 : _GEN_141; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_143 = 5'hf == io_read_0_src1_raddr ? regs_15 : _GEN_142; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_144 = 5'h10 == io_read_0_src1_raddr ? regs_16 : _GEN_143; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_145 = 5'h11 == io_read_0_src1_raddr ? regs_17 : _GEN_144; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_146 = 5'h12 == io_read_0_src1_raddr ? regs_18 : _GEN_145; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_147 = 5'h13 == io_read_0_src1_raddr ? regs_19 : _GEN_146; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_148 = 5'h14 == io_read_0_src1_raddr ? regs_20 : _GEN_147; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_149 = 5'h15 == io_read_0_src1_raddr ? regs_21 : _GEN_148; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_150 = 5'h16 == io_read_0_src1_raddr ? regs_22 : _GEN_149; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_151 = 5'h17 == io_read_0_src1_raddr ? regs_23 : _GEN_150; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_152 = 5'h18 == io_read_0_src1_raddr ? regs_24 : _GEN_151; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_153 = 5'h19 == io_read_0_src1_raddr ? regs_25 : _GEN_152; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_154 = 5'h1a == io_read_0_src1_raddr ? regs_26 : _GEN_153; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_155 = 5'h1b == io_read_0_src1_raddr ? regs_27 : _GEN_154; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_156 = 5'h1c == io_read_0_src1_raddr ? regs_28 : _GEN_155; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_157 = 5'h1d == io_read_0_src1_raddr ? regs_29 : _GEN_156; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_158 = 5'h1e == io_read_0_src1_raddr ? regs_30 : _GEN_157; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_159 = 5'h1f == io_read_0_src1_raddr ? regs_31 : _GEN_158; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_160 = io_write_0_wen & io_read_0_src1_raddr == io_write_0_waddr ? io_write_0_wdata : _GEN_159; // @[ARegfile.scala 47:29 49:78 50:33]
  wire [31:0] _GEN_161 = io_write_1_wen & io_read_0_src1_raddr == io_write_1_waddr ? io_write_1_wdata : _GEN_160; // @[ARegfile.scala 49:78 50:33]
  wire [31:0] _GEN_164 = 5'h1 == io_read_0_src2_raddr ? regs_1 : regs_0; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_165 = 5'h2 == io_read_0_src2_raddr ? regs_2 : _GEN_164; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_166 = 5'h3 == io_read_0_src2_raddr ? regs_3 : _GEN_165; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_167 = 5'h4 == io_read_0_src2_raddr ? regs_4 : _GEN_166; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_168 = 5'h5 == io_read_0_src2_raddr ? regs_5 : _GEN_167; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_169 = 5'h6 == io_read_0_src2_raddr ? regs_6 : _GEN_168; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_170 = 5'h7 == io_read_0_src2_raddr ? regs_7 : _GEN_169; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_171 = 5'h8 == io_read_0_src2_raddr ? regs_8 : _GEN_170; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_172 = 5'h9 == io_read_0_src2_raddr ? regs_9 : _GEN_171; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_173 = 5'ha == io_read_0_src2_raddr ? regs_10 : _GEN_172; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_174 = 5'hb == io_read_0_src2_raddr ? regs_11 : _GEN_173; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_175 = 5'hc == io_read_0_src2_raddr ? regs_12 : _GEN_174; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_176 = 5'hd == io_read_0_src2_raddr ? regs_13 : _GEN_175; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_177 = 5'he == io_read_0_src2_raddr ? regs_14 : _GEN_176; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_178 = 5'hf == io_read_0_src2_raddr ? regs_15 : _GEN_177; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_179 = 5'h10 == io_read_0_src2_raddr ? regs_16 : _GEN_178; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_180 = 5'h11 == io_read_0_src2_raddr ? regs_17 : _GEN_179; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_181 = 5'h12 == io_read_0_src2_raddr ? regs_18 : _GEN_180; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_182 = 5'h13 == io_read_0_src2_raddr ? regs_19 : _GEN_181; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_183 = 5'h14 == io_read_0_src2_raddr ? regs_20 : _GEN_182; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_184 = 5'h15 == io_read_0_src2_raddr ? regs_21 : _GEN_183; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_185 = 5'h16 == io_read_0_src2_raddr ? regs_22 : _GEN_184; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_186 = 5'h17 == io_read_0_src2_raddr ? regs_23 : _GEN_185; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_187 = 5'h18 == io_read_0_src2_raddr ? regs_24 : _GEN_186; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_188 = 5'h19 == io_read_0_src2_raddr ? regs_25 : _GEN_187; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_189 = 5'h1a == io_read_0_src2_raddr ? regs_26 : _GEN_188; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_190 = 5'h1b == io_read_0_src2_raddr ? regs_27 : _GEN_189; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_191 = 5'h1c == io_read_0_src2_raddr ? regs_28 : _GEN_190; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_192 = 5'h1d == io_read_0_src2_raddr ? regs_29 : _GEN_191; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_193 = 5'h1e == io_read_0_src2_raddr ? regs_30 : _GEN_192; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_194 = 5'h1f == io_read_0_src2_raddr ? regs_31 : _GEN_193; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_195 = io_write_0_wen & io_read_0_src2_raddr == io_write_0_waddr ? io_write_0_wdata : _GEN_194; // @[ARegfile.scala 58:29 60:78 61:33]
  wire [31:0] _GEN_196 = io_write_1_wen & io_read_0_src2_raddr == io_write_1_waddr ? io_write_1_wdata : _GEN_195; // @[ARegfile.scala 60:78 61:33]
  wire [31:0] _GEN_199 = 5'h1 == io_read_1_src1_raddr ? regs_1 : regs_0; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_200 = 5'h2 == io_read_1_src1_raddr ? regs_2 : _GEN_199; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_201 = 5'h3 == io_read_1_src1_raddr ? regs_3 : _GEN_200; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_202 = 5'h4 == io_read_1_src1_raddr ? regs_4 : _GEN_201; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_203 = 5'h5 == io_read_1_src1_raddr ? regs_5 : _GEN_202; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_204 = 5'h6 == io_read_1_src1_raddr ? regs_6 : _GEN_203; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_205 = 5'h7 == io_read_1_src1_raddr ? regs_7 : _GEN_204; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_206 = 5'h8 == io_read_1_src1_raddr ? regs_8 : _GEN_205; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_207 = 5'h9 == io_read_1_src1_raddr ? regs_9 : _GEN_206; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_208 = 5'ha == io_read_1_src1_raddr ? regs_10 : _GEN_207; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_209 = 5'hb == io_read_1_src1_raddr ? regs_11 : _GEN_208; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_210 = 5'hc == io_read_1_src1_raddr ? regs_12 : _GEN_209; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_211 = 5'hd == io_read_1_src1_raddr ? regs_13 : _GEN_210; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_212 = 5'he == io_read_1_src1_raddr ? regs_14 : _GEN_211; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_213 = 5'hf == io_read_1_src1_raddr ? regs_15 : _GEN_212; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_214 = 5'h10 == io_read_1_src1_raddr ? regs_16 : _GEN_213; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_215 = 5'h11 == io_read_1_src1_raddr ? regs_17 : _GEN_214; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_216 = 5'h12 == io_read_1_src1_raddr ? regs_18 : _GEN_215; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_217 = 5'h13 == io_read_1_src1_raddr ? regs_19 : _GEN_216; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_218 = 5'h14 == io_read_1_src1_raddr ? regs_20 : _GEN_217; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_219 = 5'h15 == io_read_1_src1_raddr ? regs_21 : _GEN_218; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_220 = 5'h16 == io_read_1_src1_raddr ? regs_22 : _GEN_219; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_221 = 5'h17 == io_read_1_src1_raddr ? regs_23 : _GEN_220; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_222 = 5'h18 == io_read_1_src1_raddr ? regs_24 : _GEN_221; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_223 = 5'h19 == io_read_1_src1_raddr ? regs_25 : _GEN_222; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_224 = 5'h1a == io_read_1_src1_raddr ? regs_26 : _GEN_223; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_225 = 5'h1b == io_read_1_src1_raddr ? regs_27 : _GEN_224; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_226 = 5'h1c == io_read_1_src1_raddr ? regs_28 : _GEN_225; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_227 = 5'h1d == io_read_1_src1_raddr ? regs_29 : _GEN_226; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_228 = 5'h1e == io_read_1_src1_raddr ? regs_30 : _GEN_227; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_229 = 5'h1f == io_read_1_src1_raddr ? regs_31 : _GEN_228; // @[ARegfile.scala 47:{29,29}]
  wire [31:0] _GEN_230 = io_write_0_wen & io_read_1_src1_raddr == io_write_0_waddr ? io_write_0_wdata : _GEN_229; // @[ARegfile.scala 47:29 49:78 50:33]
  wire [31:0] _GEN_231 = io_write_1_wen & io_read_1_src1_raddr == io_write_1_waddr ? io_write_1_wdata : _GEN_230; // @[ARegfile.scala 49:78 50:33]
  wire [31:0] _GEN_234 = 5'h1 == io_read_1_src2_raddr ? regs_1 : regs_0; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_235 = 5'h2 == io_read_1_src2_raddr ? regs_2 : _GEN_234; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_236 = 5'h3 == io_read_1_src2_raddr ? regs_3 : _GEN_235; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_237 = 5'h4 == io_read_1_src2_raddr ? regs_4 : _GEN_236; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_238 = 5'h5 == io_read_1_src2_raddr ? regs_5 : _GEN_237; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_239 = 5'h6 == io_read_1_src2_raddr ? regs_6 : _GEN_238; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_240 = 5'h7 == io_read_1_src2_raddr ? regs_7 : _GEN_239; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_241 = 5'h8 == io_read_1_src2_raddr ? regs_8 : _GEN_240; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_242 = 5'h9 == io_read_1_src2_raddr ? regs_9 : _GEN_241; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_243 = 5'ha == io_read_1_src2_raddr ? regs_10 : _GEN_242; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_244 = 5'hb == io_read_1_src2_raddr ? regs_11 : _GEN_243; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_245 = 5'hc == io_read_1_src2_raddr ? regs_12 : _GEN_244; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_246 = 5'hd == io_read_1_src2_raddr ? regs_13 : _GEN_245; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_247 = 5'he == io_read_1_src2_raddr ? regs_14 : _GEN_246; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_248 = 5'hf == io_read_1_src2_raddr ? regs_15 : _GEN_247; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_249 = 5'h10 == io_read_1_src2_raddr ? regs_16 : _GEN_248; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_250 = 5'h11 == io_read_1_src2_raddr ? regs_17 : _GEN_249; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_251 = 5'h12 == io_read_1_src2_raddr ? regs_18 : _GEN_250; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_252 = 5'h13 == io_read_1_src2_raddr ? regs_19 : _GEN_251; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_253 = 5'h14 == io_read_1_src2_raddr ? regs_20 : _GEN_252; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_254 = 5'h15 == io_read_1_src2_raddr ? regs_21 : _GEN_253; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_255 = 5'h16 == io_read_1_src2_raddr ? regs_22 : _GEN_254; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_256 = 5'h17 == io_read_1_src2_raddr ? regs_23 : _GEN_255; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_257 = 5'h18 == io_read_1_src2_raddr ? regs_24 : _GEN_256; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_258 = 5'h19 == io_read_1_src2_raddr ? regs_25 : _GEN_257; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_259 = 5'h1a == io_read_1_src2_raddr ? regs_26 : _GEN_258; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_260 = 5'h1b == io_read_1_src2_raddr ? regs_27 : _GEN_259; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_261 = 5'h1c == io_read_1_src2_raddr ? regs_28 : _GEN_260; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_262 = 5'h1d == io_read_1_src2_raddr ? regs_29 : _GEN_261; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_263 = 5'h1e == io_read_1_src2_raddr ? regs_30 : _GEN_262; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_264 = 5'h1f == io_read_1_src2_raddr ? regs_31 : _GEN_263; // @[ARegfile.scala 58:{29,29}]
  wire [31:0] _GEN_265 = io_write_0_wen & io_read_1_src2_raddr == io_write_0_waddr ? io_write_0_wdata : _GEN_264; // @[ARegfile.scala 58:29 60:78 61:33]
  wire [31:0] _GEN_266 = io_write_1_wen & io_read_1_src2_raddr == io_write_1_waddr ? io_write_1_wdata : _GEN_265; // @[ARegfile.scala 60:78 61:33]
  assign io_read_0_src1_rdata = io_read_0_src1_raddr == 5'h0 ? 32'h0 : _GEN_161; // @[ARegfile.scala 44:41 45:29]
  assign io_read_0_src2_rdata = io_read_0_src2_raddr == 5'h0 ? 32'h0 : _GEN_196; // @[ARegfile.scala 55:41 56:29]
  assign io_read_1_src1_rdata = io_read_1_src1_raddr == 5'h0 ? 32'h0 : _GEN_231; // @[ARegfile.scala 44:41 45:29]
  assign io_read_1_src2_rdata = io_read_1_src2_raddr == 5'h0 ? 32'h0 : _GEN_266; // @[ARegfile.scala 55:41 56:29]
  always @(posedge clock) begin
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_0 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h0 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_0 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_0 <= _GEN_32;
      end
    end else begin
      regs_0 <= _GEN_32;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_1 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h1 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_1 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_1 <= _GEN_33;
      end
    end else begin
      regs_1 <= _GEN_33;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_2 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h2 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_2 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_2 <= _GEN_34;
      end
    end else begin
      regs_2 <= _GEN_34;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_3 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h3 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_3 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_3 <= _GEN_35;
      end
    end else begin
      regs_3 <= _GEN_35;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_4 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h4 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_4 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_4 <= _GEN_36;
      end
    end else begin
      regs_4 <= _GEN_36;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_5 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h5 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_5 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_5 <= _GEN_37;
      end
    end else begin
      regs_5 <= _GEN_37;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_6 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h6 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_6 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_6 <= _GEN_38;
      end
    end else begin
      regs_6 <= _GEN_38;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_7 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h7 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_7 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_7 <= _GEN_39;
      end
    end else begin
      regs_7 <= _GEN_39;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_8 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h8 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_8 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_8 <= _GEN_40;
      end
    end else begin
      regs_8 <= _GEN_40;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_9 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h9 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_9 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_9 <= _GEN_41;
      end
    end else begin
      regs_9 <= _GEN_41;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_10 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'ha == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_10 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_10 <= _GEN_42;
      end
    end else begin
      regs_10 <= _GEN_42;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_11 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'hb == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_11 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_11 <= _GEN_43;
      end
    end else begin
      regs_11 <= _GEN_43;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_12 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'hc == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_12 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_12 <= _GEN_44;
      end
    end else begin
      regs_12 <= _GEN_44;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_13 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'hd == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_13 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_13 <= _GEN_45;
      end
    end else begin
      regs_13 <= _GEN_45;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_14 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'he == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_14 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_14 <= _GEN_46;
      end
    end else begin
      regs_14 <= _GEN_46;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_15 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'hf == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_15 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_15 <= _GEN_47;
      end
    end else begin
      regs_15 <= _GEN_47;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_16 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h10 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_16 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_16 <= _GEN_48;
      end
    end else begin
      regs_16 <= _GEN_48;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_17 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h11 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_17 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_17 <= _GEN_49;
      end
    end else begin
      regs_17 <= _GEN_49;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_18 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h12 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_18 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_18 <= _GEN_50;
      end
    end else begin
      regs_18 <= _GEN_50;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_19 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h13 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_19 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_19 <= _GEN_51;
      end
    end else begin
      regs_19 <= _GEN_51;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_20 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h14 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_20 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_20 <= _GEN_52;
      end
    end else begin
      regs_20 <= _GEN_52;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_21 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h15 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_21 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_21 <= _GEN_53;
      end
    end else begin
      regs_21 <= _GEN_53;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_22 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h16 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_22 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_22 <= _GEN_54;
      end
    end else begin
      regs_22 <= _GEN_54;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_23 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h17 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_23 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_23 <= _GEN_55;
      end
    end else begin
      regs_23 <= _GEN_55;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_24 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h18 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_24 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_24 <= _GEN_56;
      end
    end else begin
      regs_24 <= _GEN_56;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_25 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h19 == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_25 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_25 <= _GEN_57;
      end
    end else begin
      regs_25 <= _GEN_57;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_26 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h1a == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_26 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_26 <= _GEN_58;
      end
    end else begin
      regs_26 <= _GEN_58;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_27 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h1b == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_27 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_27 <= _GEN_59;
      end
    end else begin
      regs_27 <= _GEN_59;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_28 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h1c == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_28 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_28 <= _GEN_60;
      end
    end else begin
      regs_28 <= _GEN_60;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_29 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h1d == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_29 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_29 <= _GEN_61;
      end
    end else begin
      regs_29 <= _GEN_61;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_30 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h1e == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_30 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_30 <= _GEN_62;
      end
    end else begin
      regs_30 <= _GEN_62;
    end
    if (reset) begin // @[ARegfile.scala 32:21]
      regs_31 <= 32'h0; // @[ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[ARegfile.scala 36:56]
      if (5'h1f == io_write_1_waddr) begin // @[ARegfile.scala 37:31]
        regs_31 <= io_write_1_wdata; // @[ARegfile.scala 37:31]
      end else begin
        regs_31 <= _GEN_63;
      end
    end else begin
      regs_31 <= _GEN_63;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ExecuteStage(
  input         clock,
  input         reset,
  input         io_ctrl_inst0_allow_to_go,
  input         io_ctrl_clear_0,
  input         io_ctrl_clear_1,
  input  [31:0] io_decoderUnit_inst0_pc,
  input  [3:0]  io_decoderUnit_inst0_inst_info_fusel,
  input  [6:0]  io_decoderUnit_inst0_inst_info_op,
  input         io_decoderUnit_inst0_inst_info_reg_wen,
  input  [4:0]  io_decoderUnit_inst0_inst_info_reg_waddr,
  input  [7:0]  io_decoderUnit_inst0_inst_info_cp0_addr,
  input  [31:0] io_decoderUnit_inst0_inst_info_inst,
  input  [31:0] io_decoderUnit_inst0_src_info_src1_data,
  input  [31:0] io_decoderUnit_inst0_src_info_src2_data,
  input         io_decoderUnit_inst0_ex_flush_req,
  input         io_decoderUnit_inst0_ex_eret,
  input  [31:0] io_decoderUnit_inst0_ex_badvaddr,
  input         io_decoderUnit_inst0_ex_bd,
  input  [4:0]  io_decoderUnit_inst0_ex_excode,
  input         io_decoderUnit_inst0_jb_info_jump_regiser_conflict,
  input         io_decoderUnit_inst0_jb_info_is_branch,
  input         io_decoderUnit_inst0_jb_info_pred_branch_flag,
  input  [31:0] io_decoderUnit_inst0_jb_info_branch_target,
  input         io_decoderUnit_inst1_allow_to_go,
  input  [31:0] io_decoderUnit_inst1_pc,
  input  [3:0]  io_decoderUnit_inst1_inst_info_fusel,
  input  [6:0]  io_decoderUnit_inst1_inst_info_op,
  input         io_decoderUnit_inst1_inst_info_reg_wen,
  input  [4:0]  io_decoderUnit_inst1_inst_info_reg_waddr,
  input  [31:0] io_decoderUnit_inst1_inst_info_inst,
  input  [31:0] io_decoderUnit_inst1_src_info_src1_data,
  input  [31:0] io_decoderUnit_inst1_src_info_src2_data,
  input         io_decoderUnit_inst1_ex_flush_req,
  input         io_decoderUnit_inst1_ex_eret,
  input  [31:0] io_decoderUnit_inst1_ex_badvaddr,
  input         io_decoderUnit_inst1_ex_bd,
  input  [4:0]  io_decoderUnit_inst1_ex_excode,
  output [31:0] io_executeUnit_inst0_pc,
  output [3:0]  io_executeUnit_inst0_inst_info_fusel,
  output [6:0]  io_executeUnit_inst0_inst_info_op,
  output        io_executeUnit_inst0_inst_info_reg_wen,
  output [4:0]  io_executeUnit_inst0_inst_info_reg_waddr,
  output [7:0]  io_executeUnit_inst0_inst_info_cp0_addr,
  output [31:0] io_executeUnit_inst0_inst_info_inst,
  output [31:0] io_executeUnit_inst0_src_info_src1_data,
  output [31:0] io_executeUnit_inst0_src_info_src2_data,
  output        io_executeUnit_inst0_ex_flush_req,
  output        io_executeUnit_inst0_ex_eret,
  output [31:0] io_executeUnit_inst0_ex_badvaddr,
  output        io_executeUnit_inst0_ex_bd,
  output [4:0]  io_executeUnit_inst0_ex_excode,
  output        io_executeUnit_inst0_jb_info_jump_regiser_conflict,
  output        io_executeUnit_inst0_jb_info_is_branch,
  output        io_executeUnit_inst0_jb_info_pred_branch_flag,
  output [31:0] io_executeUnit_inst0_jb_info_branch_target,
  output [31:0] io_executeUnit_inst1_pc,
  output [3:0]  io_executeUnit_inst1_inst_info_fusel,
  output [6:0]  io_executeUnit_inst1_inst_info_op,
  output        io_executeUnit_inst1_inst_info_reg_wen,
  output [4:0]  io_executeUnit_inst1_inst_info_reg_waddr,
  output [31:0] io_executeUnit_inst1_inst_info_inst,
  output [31:0] io_executeUnit_inst1_src_info_src1_data,
  output [31:0] io_executeUnit_inst1_src_info_src2_data,
  output        io_executeUnit_inst1_ex_flush_req,
  output        io_executeUnit_inst1_ex_eret,
  output [31:0] io_executeUnit_inst1_ex_badvaddr,
  output        io_executeUnit_inst1_ex_bd,
  output [4:0]  io_executeUnit_inst1_ex_excode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] inst0_pc; // @[ExecuteStage.scala 47:22]
  reg [3:0] inst0_inst_info_fusel; // @[ExecuteStage.scala 47:22]
  reg [6:0] inst0_inst_info_op; // @[ExecuteStage.scala 47:22]
  reg  inst0_inst_info_reg_wen; // @[ExecuteStage.scala 47:22]
  reg [4:0] inst0_inst_info_reg_waddr; // @[ExecuteStage.scala 47:22]
  reg [7:0] inst0_inst_info_cp0_addr; // @[ExecuteStage.scala 47:22]
  reg [31:0] inst0_inst_info_inst; // @[ExecuteStage.scala 47:22]
  reg [31:0] inst0_src_info_src1_data; // @[ExecuteStage.scala 47:22]
  reg [31:0] inst0_src_info_src2_data; // @[ExecuteStage.scala 47:22]
  reg  inst0_ex_flush_req; // @[ExecuteStage.scala 47:22]
  reg  inst0_ex_eret; // @[ExecuteStage.scala 47:22]
  reg [31:0] inst0_ex_badvaddr; // @[ExecuteStage.scala 47:22]
  reg  inst0_ex_bd; // @[ExecuteStage.scala 47:22]
  reg [4:0] inst0_ex_excode; // @[ExecuteStage.scala 47:22]
  reg  inst0_jb_info_jump_regiser_conflict; // @[ExecuteStage.scala 47:22]
  reg  inst0_jb_info_is_branch; // @[ExecuteStage.scala 47:22]
  reg  inst0_jb_info_pred_branch_flag; // @[ExecuteStage.scala 47:22]
  reg [31:0] inst0_jb_info_branch_target; // @[ExecuteStage.scala 47:22]
  reg [31:0] inst1_pc; // @[ExecuteStage.scala 48:22]
  reg [3:0] inst1_inst_info_fusel; // @[ExecuteStage.scala 48:22]
  reg [6:0] inst1_inst_info_op; // @[ExecuteStage.scala 48:22]
  reg  inst1_inst_info_reg_wen; // @[ExecuteStage.scala 48:22]
  reg [4:0] inst1_inst_info_reg_waddr; // @[ExecuteStage.scala 48:22]
  reg [31:0] inst1_inst_info_inst; // @[ExecuteStage.scala 48:22]
  reg [31:0] inst1_src_info_src1_data; // @[ExecuteStage.scala 48:22]
  reg [31:0] inst1_src_info_src2_data; // @[ExecuteStage.scala 48:22]
  reg  inst1_ex_flush_req; // @[ExecuteStage.scala 48:22]
  reg  inst1_ex_eret; // @[ExecuteStage.scala 48:22]
  reg [31:0] inst1_ex_badvaddr; // @[ExecuteStage.scala 48:22]
  reg  inst1_ex_bd; // @[ExecuteStage.scala 48:22]
  reg [4:0] inst1_ex_excode; // @[ExecuteStage.scala 48:22]
  assign io_executeUnit_inst0_pc = inst0_pc; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_inst_info_fusel = inst0_inst_info_fusel; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_inst_info_op = inst0_inst_info_op; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_inst_info_reg_wen = inst0_inst_info_reg_wen; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_inst_info_reg_waddr = inst0_inst_info_reg_waddr; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_inst_info_cp0_addr = inst0_inst_info_cp0_addr; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_inst_info_inst = inst0_inst_info_inst; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_src_info_src1_data = inst0_src_info_src1_data; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_src_info_src2_data = inst0_src_info_src2_data; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_ex_flush_req = inst0_ex_flush_req; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_ex_eret = inst0_ex_eret; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_ex_badvaddr = inst0_ex_badvaddr; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_ex_bd = inst0_ex_bd; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_ex_excode = inst0_ex_excode; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_jb_info_jump_regiser_conflict = inst0_jb_info_jump_regiser_conflict; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_jb_info_is_branch = inst0_jb_info_is_branch; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_jb_info_pred_branch_flag = inst0_jb_info_pred_branch_flag; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst0_jb_info_branch_target = inst0_jb_info_branch_target; // @[ExecuteStage.scala 62:24]
  assign io_executeUnit_inst1_pc = inst1_pc; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_inst_info_fusel = inst1_inst_info_fusel; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_inst_info_op = inst1_inst_info_op; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_inst_info_reg_wen = inst1_inst_info_reg_wen; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_inst_info_reg_waddr = inst1_inst_info_reg_waddr; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_inst_info_inst = inst1_inst_info_inst; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_src_info_src1_data = inst1_src_info_src1_data; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_src_info_src2_data = inst1_src_info_src2_data; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_ex_flush_req = inst1_ex_flush_req; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_ex_eret = inst1_ex_eret; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_ex_badvaddr = inst1_ex_badvaddr; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_ex_bd = inst1_ex_bd; // @[ExecuteStage.scala 63:24]
  assign io_executeUnit_inst1_ex_excode = inst1_ex_excode; // @[ExecuteStage.scala 63:24]
  always @(posedge clock) begin
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_pc <= 32'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_pc <= 32'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_pc <= io_decoderUnit_inst0_pc; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_inst_info_fusel <= 4'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_inst_info_fusel <= 4'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_inst_info_fusel <= io_decoderUnit_inst0_inst_info_fusel; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_inst_info_op <= 7'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_inst_info_op <= 7'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_inst_info_op <= io_decoderUnit_inst0_inst_info_op; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_inst_info_reg_wen <= 1'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_inst_info_reg_wen <= 1'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_inst_info_reg_wen <= io_decoderUnit_inst0_inst_info_reg_wen; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_inst_info_reg_waddr <= 5'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_inst_info_reg_waddr <= 5'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_inst_info_reg_waddr <= io_decoderUnit_inst0_inst_info_reg_waddr; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_inst_info_cp0_addr <= 8'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_inst_info_cp0_addr <= 8'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_inst_info_cp0_addr <= io_decoderUnit_inst0_inst_info_cp0_addr; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_inst_info_inst <= 32'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_inst_info_inst <= 32'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_inst_info_inst <= io_decoderUnit_inst0_inst_info_inst; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_src_info_src1_data <= 32'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_src_info_src1_data <= 32'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_src_info_src1_data <= io_decoderUnit_inst0_src_info_src1_data; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_src_info_src2_data <= 32'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_src_info_src2_data <= 32'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_src_info_src2_data <= io_decoderUnit_inst0_src_info_src2_data; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_ex_flush_req <= 1'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_ex_flush_req <= 1'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_ex_flush_req <= io_decoderUnit_inst0_ex_flush_req; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_ex_eret <= 1'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_ex_eret <= 1'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_ex_eret <= io_decoderUnit_inst0_ex_eret; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_ex_badvaddr <= 32'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_ex_badvaddr <= 32'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_ex_badvaddr <= io_decoderUnit_inst0_ex_badvaddr; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_ex_bd <= 1'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_ex_bd <= 1'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_ex_bd <= io_decoderUnit_inst0_ex_bd; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_ex_excode <= 5'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_ex_excode <= 5'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_ex_excode <= io_decoderUnit_inst0_ex_excode; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_jb_info_jump_regiser_conflict <= 1'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_jb_info_jump_regiser_conflict <= 1'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_jb_info_jump_regiser_conflict <= io_decoderUnit_inst0_jb_info_jump_regiser_conflict; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_jb_info_is_branch <= 1'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_jb_info_is_branch <= 1'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_jb_info_is_branch <= io_decoderUnit_inst0_jb_info_is_branch; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_jb_info_pred_branch_flag <= 1'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_jb_info_pred_branch_flag <= 1'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_jb_info_pred_branch_flag <= io_decoderUnit_inst0_jb_info_pred_branch_flag; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 47:22]
      inst0_jb_info_branch_target <= 32'h0; // @[ExecuteStage.scala 47:22]
    end else if (io_ctrl_clear_0) begin // @[ExecuteStage.scala 50:26]
      inst0_jb_info_branch_target <= 32'h0; // @[ExecuteStage.scala 51:11]
    end else if (io_ctrl_inst0_allow_to_go) begin // @[ExecuteStage.scala 52:41]
      inst0_jb_info_branch_target <= io_decoderUnit_inst0_jb_info_branch_target; // @[ExecuteStage.scala 53:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_pc <= 32'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_pc <= 32'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_pc <= io_decoderUnit_inst1_pc; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_inst_info_fusel <= 4'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_inst_info_fusel <= 4'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_inst_info_fusel <= io_decoderUnit_inst1_inst_info_fusel; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_inst_info_op <= 7'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_inst_info_op <= 7'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_inst_info_op <= io_decoderUnit_inst1_inst_info_op; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_inst_info_reg_wen <= 1'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_inst_info_reg_wen <= 1'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_inst_info_reg_wen <= io_decoderUnit_inst1_inst_info_reg_wen; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_inst_info_reg_waddr <= 5'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_inst_info_reg_waddr <= 5'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_inst_info_reg_waddr <= io_decoderUnit_inst1_inst_info_reg_waddr; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_inst_info_inst <= 32'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_inst_info_inst <= 32'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_inst_info_inst <= io_decoderUnit_inst1_inst_info_inst; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_src_info_src1_data <= 32'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_src_info_src1_data <= 32'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_src_info_src1_data <= io_decoderUnit_inst1_src_info_src1_data; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_src_info_src2_data <= 32'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_src_info_src2_data <= 32'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_src_info_src2_data <= io_decoderUnit_inst1_src_info_src2_data; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_ex_flush_req <= 1'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_ex_flush_req <= 1'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_ex_flush_req <= io_decoderUnit_inst1_ex_flush_req; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_ex_eret <= 1'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_ex_eret <= 1'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_ex_eret <= io_decoderUnit_inst1_ex_eret; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_ex_badvaddr <= 32'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_ex_badvaddr <= 32'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_ex_badvaddr <= io_decoderUnit_inst1_ex_badvaddr; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_ex_bd <= 1'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_ex_bd <= 1'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_ex_bd <= io_decoderUnit_inst1_ex_bd; // @[ExecuteStage.scala 59:11]
    end
    if (reset) begin // @[ExecuteStage.scala 48:22]
      inst1_ex_excode <= 5'h0; // @[ExecuteStage.scala 48:22]
    end else if (io_ctrl_clear_1) begin // @[ExecuteStage.scala 56:26]
      inst1_ex_excode <= 5'h0; // @[ExecuteStage.scala 57:11]
    end else if (io_decoderUnit_inst1_allow_to_go) begin // @[ExecuteStage.scala 58:48]
      inst1_ex_excode <= io_decoderUnit_inst1_ex_excode; // @[ExecuteStage.scala 59:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst0_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  inst0_inst_info_fusel = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  inst0_inst_info_op = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  inst0_inst_info_reg_wen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  inst0_inst_info_reg_waddr = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  inst0_inst_info_cp0_addr = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  inst0_inst_info_inst = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  inst0_src_info_src1_data = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  inst0_src_info_src2_data = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  inst0_ex_flush_req = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  inst0_ex_eret = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inst0_ex_badvaddr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  inst0_ex_bd = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inst0_ex_excode = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  inst0_jb_info_jump_regiser_conflict = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  inst0_jb_info_is_branch = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  inst0_jb_info_pred_branch_flag = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  inst0_jb_info_branch_target = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  inst1_pc = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inst1_inst_info_fusel = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  inst1_inst_info_op = _RAND_20[6:0];
  _RAND_21 = {1{`RANDOM}};
  inst1_inst_info_reg_wen = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  inst1_inst_info_reg_waddr = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  inst1_inst_info_inst = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  inst1_src_info_src1_data = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  inst1_src_info_src2_data = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  inst1_ex_flush_req = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  inst1_ex_eret = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  inst1_ex_badvaddr = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inst1_ex_bd = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  inst1_ex_excode = _RAND_30[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Alu(
  input  [6:0]  io_inst_info_op,
  input  [31:0] io_src_info_src1_data,
  input  [31:0] io_src_info_src2_data,
  input  [31:0] io_cp0_rdata,
  input  [63:0] io_hilo_rdata,
  output [63:0] io_hilo_wdata,
  input         io_mul_ready,
  input  [63:0] io_mul_result,
  output        io_mul_start,
  output        io_mul_signed,
  input         io_div_ready,
  input  [63:0] io_div_result,
  output        io_div_start,
  output        io_div_signed,
  output [31:0] io_result,
  output        io_overflow
);
  wire [31:0] sum = io_src_info_src1_data + io_src_info_src2_data; // @[ALU.scala 34:19]
  wire [31:0] diff = io_src_info_src1_data - io_src_info_src2_data; // @[ALU.scala 35:19]
  wire  slt = $signed(io_src_info_src1_data) < $signed(io_src_info_src2_data); // @[ALU.scala 36:28]
  wire  sltu = io_src_info_src1_data < io_src_info_src2_data; // @[ALU.scala 37:19]
  wire [5:0] _GEN_0 = ~io_src_info_src1_data[0] ? 6'h1f : 6'h20; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_1 = ~io_src_info_src1_data[0] ? 6'h20 : 6'h1f; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_2 = ~io_src_info_src1_data[1] ? 6'h1e : _GEN_0; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_3 = ~io_src_info_src1_data[1] ? _GEN_1 : 6'h1e; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_4 = ~io_src_info_src1_data[2] ? 6'h1d : _GEN_2; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_5 = ~io_src_info_src1_data[2] ? _GEN_3 : 6'h1d; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_6 = ~io_src_info_src1_data[3] ? 6'h1c : _GEN_4; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_7 = ~io_src_info_src1_data[3] ? _GEN_5 : 6'h1c; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_8 = ~io_src_info_src1_data[4] ? 6'h1b : _GEN_6; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_9 = ~io_src_info_src1_data[4] ? _GEN_7 : 6'h1b; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_10 = ~io_src_info_src1_data[5] ? 6'h1a : _GEN_8; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_11 = ~io_src_info_src1_data[5] ? _GEN_9 : 6'h1a; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_12 = ~io_src_info_src1_data[6] ? 6'h19 : _GEN_10; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_13 = ~io_src_info_src1_data[6] ? _GEN_11 : 6'h19; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_14 = ~io_src_info_src1_data[7] ? 6'h18 : _GEN_12; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_15 = ~io_src_info_src1_data[7] ? _GEN_13 : 6'h18; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_16 = ~io_src_info_src1_data[8] ? 6'h17 : _GEN_14; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_17 = ~io_src_info_src1_data[8] ? _GEN_15 : 6'h17; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_18 = ~io_src_info_src1_data[9] ? 6'h16 : _GEN_16; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_19 = ~io_src_info_src1_data[9] ? _GEN_17 : 6'h16; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_20 = ~io_src_info_src1_data[10] ? 6'h15 : _GEN_18; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_21 = ~io_src_info_src1_data[10] ? _GEN_19 : 6'h15; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_22 = ~io_src_info_src1_data[11] ? 6'h14 : _GEN_20; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_23 = ~io_src_info_src1_data[11] ? _GEN_21 : 6'h14; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_24 = ~io_src_info_src1_data[12] ? 6'h13 : _GEN_22; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_25 = ~io_src_info_src1_data[12] ? _GEN_23 : 6'h13; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_26 = ~io_src_info_src1_data[13] ? 6'h12 : _GEN_24; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_27 = ~io_src_info_src1_data[13] ? _GEN_25 : 6'h12; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_28 = ~io_src_info_src1_data[14] ? 6'h11 : _GEN_26; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_29 = ~io_src_info_src1_data[14] ? _GEN_27 : 6'h11; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_30 = ~io_src_info_src1_data[15] ? 6'h10 : _GEN_28; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_31 = ~io_src_info_src1_data[15] ? _GEN_29 : 6'h10; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_32 = ~io_src_info_src1_data[16] ? 6'hf : _GEN_30; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_33 = ~io_src_info_src1_data[16] ? _GEN_31 : 6'hf; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_34 = ~io_src_info_src1_data[17] ? 6'he : _GEN_32; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_35 = ~io_src_info_src1_data[17] ? _GEN_33 : 6'he; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_36 = ~io_src_info_src1_data[18] ? 6'hd : _GEN_34; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_37 = ~io_src_info_src1_data[18] ? _GEN_35 : 6'hd; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_38 = ~io_src_info_src1_data[19] ? 6'hc : _GEN_36; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_39 = ~io_src_info_src1_data[19] ? _GEN_37 : 6'hc; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_40 = ~io_src_info_src1_data[20] ? 6'hb : _GEN_38; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_41 = ~io_src_info_src1_data[20] ? _GEN_39 : 6'hb; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_42 = ~io_src_info_src1_data[21] ? 6'ha : _GEN_40; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_43 = ~io_src_info_src1_data[21] ? _GEN_41 : 6'ha; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_44 = ~io_src_info_src1_data[22] ? 6'h9 : _GEN_42; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_45 = ~io_src_info_src1_data[22] ? _GEN_43 : 6'h9; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_46 = ~io_src_info_src1_data[23] ? 6'h8 : _GEN_44; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_47 = ~io_src_info_src1_data[23] ? _GEN_45 : 6'h8; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_48 = ~io_src_info_src1_data[24] ? 6'h7 : _GEN_46; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_49 = ~io_src_info_src1_data[24] ? _GEN_47 : 6'h7; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_50 = ~io_src_info_src1_data[25] ? 6'h6 : _GEN_48; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_51 = ~io_src_info_src1_data[25] ? _GEN_49 : 6'h6; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_52 = ~io_src_info_src1_data[26] ? 6'h5 : _GEN_50; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_53 = ~io_src_info_src1_data[26] ? _GEN_51 : 6'h5; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_54 = ~io_src_info_src1_data[27] ? 6'h4 : _GEN_52; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_55 = ~io_src_info_src1_data[27] ? _GEN_53 : 6'h4; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_56 = ~io_src_info_src1_data[28] ? 6'h3 : _GEN_54; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_57 = ~io_src_info_src1_data[28] ? _GEN_55 : 6'h3; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_58 = ~io_src_info_src1_data[29] ? 6'h2 : _GEN_56; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_59 = ~io_src_info_src1_data[29] ? _GEN_57 : 6'h2; // @[ALU.scala 41:20 44:11]
  wire [5:0] _GEN_60 = ~io_src_info_src1_data[30] ? 6'h1 : _GEN_58; // @[ALU.scala 41:20 42:11]
  wire [5:0] _GEN_61 = ~io_src_info_src1_data[30] ? _GEN_59 : 6'h1; // @[ALU.scala 41:20 44:11]
  wire [5:0] clo = ~io_src_info_src1_data[31] ? 6'h0 : _GEN_60; // @[ALU.scala 41:20 42:11]
  wire [5:0] clz = ~io_src_info_src1_data[31] ? _GEN_61 : 6'h0; // @[ALU.scala 41:20 44:11]
  wire [63:0] _io_hilo_wdata_T_1 = {io_src_info_src1_data,io_hilo_rdata[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _io_hilo_wdata_T_3 = {io_hilo_rdata[63:32],io_src_info_src1_data}; // @[Cat.scala 33:92]
  wire [63:0] _io_hilo_wdata_T_4 = io_mul_ready ? io_mul_result : 64'h0; // @[ALU.scala 56:23]
  wire [63:0] _io_hilo_wdata_T_7 = io_hilo_rdata + io_mul_result; // @[ALU.scala 58:43]
  wire [63:0] _io_hilo_wdata_T_8 = io_mul_ready ? _io_hilo_wdata_T_7 : 64'h0; // @[ALU.scala 58:23]
  wire [63:0] _io_hilo_wdata_T_13 = io_hilo_rdata - io_mul_result; // @[ALU.scala 60:43]
  wire [63:0] _io_hilo_wdata_T_14 = io_mul_ready ? _io_hilo_wdata_T_13 : 64'h0; // @[ALU.scala 60:23]
  wire [63:0] _io_hilo_wdata_T_18 = io_div_ready ? io_div_result : 64'h0; // @[ALU.scala 62:23]
  wire [63:0] _io_hilo_wdata_T_21 = 7'he == io_inst_info_op ? _io_hilo_wdata_T_1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_hilo_wdata_T_23 = 7'h10 == io_inst_info_op ? _io_hilo_wdata_T_3 : _io_hilo_wdata_T_21; // @[Mux.scala 81:58]
  wire  _io_hilo_wdata_T_24 = 7'h1b == io_inst_info_op; // @[Mux.scala 81:61]
  wire [63:0] _io_hilo_wdata_T_25 = 7'h1b == io_inst_info_op ? _io_hilo_wdata_T_4 : _io_hilo_wdata_T_23; // @[Mux.scala 81:58]
  wire  _io_hilo_wdata_T_26 = 7'h1c == io_inst_info_op; // @[Mux.scala 81:61]
  wire [63:0] _io_hilo_wdata_T_27 = 7'h1c == io_inst_info_op ? _io_hilo_wdata_T_4 : _io_hilo_wdata_T_25; // @[Mux.scala 81:58]
  wire  _io_hilo_wdata_T_28 = 7'h1e == io_inst_info_op; // @[Mux.scala 81:61]
  wire [63:0] _io_hilo_wdata_T_29 = 7'h1e == io_inst_info_op ? _io_hilo_wdata_T_8 : _io_hilo_wdata_T_27; // @[Mux.scala 81:58]
  wire  _io_hilo_wdata_T_30 = 7'h1f == io_inst_info_op; // @[Mux.scala 81:61]
  wire [63:0] _io_hilo_wdata_T_31 = 7'h1f == io_inst_info_op ? _io_hilo_wdata_T_8 : _io_hilo_wdata_T_29; // @[Mux.scala 81:58]
  wire  _io_hilo_wdata_T_32 = 7'h20 == io_inst_info_op; // @[Mux.scala 81:61]
  wire [63:0] _io_hilo_wdata_T_33 = 7'h20 == io_inst_info_op ? _io_hilo_wdata_T_14 : _io_hilo_wdata_T_31; // @[Mux.scala 81:58]
  wire  _io_hilo_wdata_T_34 = 7'h21 == io_inst_info_op; // @[Mux.scala 81:61]
  wire [63:0] _io_hilo_wdata_T_35 = 7'h21 == io_inst_info_op ? _io_hilo_wdata_T_14 : _io_hilo_wdata_T_33; // @[Mux.scala 81:58]
  wire  _io_hilo_wdata_T_36 = 7'h22 == io_inst_info_op; // @[Mux.scala 81:61]
  wire [63:0] _io_hilo_wdata_T_37 = 7'h22 == io_inst_info_op ? _io_hilo_wdata_T_18 : _io_hilo_wdata_T_35; // @[Mux.scala 81:58]
  wire  _io_hilo_wdata_T_38 = 7'h23 == io_inst_info_op; // @[Mux.scala 81:61]
  wire  _io_mul_start_T_11 = _io_hilo_wdata_T_24 | _io_hilo_wdata_T_26 | _io_hilo_wdata_T_28 | _io_hilo_wdata_T_32 |
    _io_hilo_wdata_T_30 | _io_hilo_wdata_T_34; // @[ALU.scala 69:84]
  wire  _io_mul_start_T_12 = ~io_mul_ready; // @[ALU.scala 70:5]
  wire [31:0] _io_result_T = io_src_info_src1_data & io_src_info_src2_data; // @[ALU.scala 88:24]
  wire [31:0] _io_result_T_1 = io_src_info_src1_data | io_src_info_src2_data; // @[ALU.scala 89:24]
  wire [31:0] _io_result_T_3 = ~_io_result_T_1; // @[ALU.scala 90:19]
  wire [31:0] _io_result_T_4 = io_src_info_src1_data ^ io_src_info_src2_data; // @[ALU.scala 91:24]
  wire [62:0] _GEN_64 = {{31'd0}, io_src_info_src2_data}; // @[ALU.scala 93:24]
  wire [62:0] _io_result_T_6 = _GEN_64 << io_src_info_src1_data[4:0]; // @[ALU.scala 93:24]
  wire [31:0] _io_result_T_8 = io_src_info_src2_data >> io_src_info_src1_data[4:0]; // @[ALU.scala 94:24]
  wire [31:0] _io_result_T_12 = $signed(io_src_info_src2_data) >>> io_src_info_src1_data[4:0]; // @[ALU.scala 95:47]
  wire [31:0] _io_result_T_16 = io_mul_ready ? io_mul_result[31:0] : 32'h0; // @[ALU.scala 108:23]
  wire [31:0] _io_result_T_20 = 7'h15 == io_inst_info_op ? sum : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_22 = 7'h16 == io_inst_info_op ? sum : _io_result_T_20; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_24 = 7'h17 == io_inst_info_op ? diff : _io_result_T_22; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_26 = 7'h18 == io_inst_info_op ? diff : _io_result_T_24; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_28 = 7'h13 == io_inst_info_op ? {{31'd0}, slt} : _io_result_T_26; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_30 = 7'h14 == io_inst_info_op ? {{31'd0}, sltu} : _io_result_T_28; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_32 = 7'h1 == io_inst_info_op ? _io_result_T : _io_result_T_30; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_34 = 7'h2 == io_inst_info_op ? _io_result_T_1 : _io_result_T_32; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_36 = 7'h4 == io_inst_info_op ? _io_result_T_3 : _io_result_T_34; // @[Mux.scala 81:58]
  wire [31:0] _io_result_T_38 = 7'h3 == io_inst_info_op ? _io_result_T_4 : _io_result_T_36; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_40 = 7'h5 == io_inst_info_op ? _io_result_T_6 : {{31'd0}, _io_result_T_38}; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_42 = 7'h7 == io_inst_info_op ? {{31'd0}, _io_result_T_8} : _io_result_T_40; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_44 = 7'h9 == io_inst_info_op ? {{31'd0}, _io_result_T_12} : _io_result_T_42; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_46 = 7'hd == io_inst_info_op ? {{31'd0}, io_hilo_rdata[63:32]} : _io_result_T_44; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_48 = 7'hf == io_inst_info_op ? {{31'd0}, io_hilo_rdata[31:0]} : _io_result_T_46; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_50 = 7'h11 == io_inst_info_op ? {{31'd0}, io_cp0_rdata} : _io_result_T_48; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_52 = 7'hc == io_inst_info_op ? {{31'd0}, io_src_info_src1_data} : _io_result_T_50; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_54 = 7'hc == io_inst_info_op ? {{31'd0}, io_src_info_src1_data} : _io_result_T_52; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_56 = 7'h19 == io_inst_info_op ? {{57'd0}, clz} : _io_result_T_54; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_58 = 7'h1a == io_inst_info_op ? {{57'd0}, clo} : _io_result_T_56; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_60 = 7'h39 == io_inst_info_op ? 63'h1 : _io_result_T_58; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_62 = 7'h1b == io_inst_info_op ? {{31'd0}, _io_result_T_16} : _io_result_T_60; // @[Mux.scala 81:58]
  wire [62:0] _io_result_T_64 = 7'h1c == io_inst_info_op ? {{31'd0}, _io_result_T_16} : _io_result_T_62; // @[Mux.scala 81:58]
  wire  _io_overflow_T_6 = io_src_info_src1_data[31] == io_src_info_src2_data[31] & io_src_info_src1_data[31] != sum[31]
    ; // @[ALU.scala 117:43]
  wire  _io_overflow_T_13 = io_src_info_src1_data[31] != io_src_info_src2_data[31] & io_src_info_src1_data[31] != diff[
    31]; // @[ALU.scala 118:43]
  assign io_hilo_wdata = 7'h23 == io_inst_info_op ? _io_hilo_wdata_T_18 : _io_hilo_wdata_T_37; // @[Mux.scala 81:58]
  assign io_mul_start = _io_mul_start_T_11 & _io_mul_start_T_12; // @[ALU.scala 68:22]
  assign io_mul_signed = _io_hilo_wdata_T_24 | _io_hilo_wdata_T_28 | _io_hilo_wdata_T_32; // @[ALU.scala 67:70]
  assign io_div_start = (_io_hilo_wdata_T_36 | _io_hilo_wdata_T_38) & ~io_div_ready; // @[ALU.scala 74:23]
  assign io_div_signed = 7'h22 == io_inst_info_op; // @[ALU.scala 73:49]
  assign io_result = _io_result_T_64[31:0]; // @[ALU.scala 76:13]
  assign io_overflow = 7'h17 == io_inst_info_op ? _io_overflow_T_13 : 7'h15 == io_inst_info_op & _io_overflow_T_6; // @[Mux.scala 81:58]
endmodule
module Mul(
  input         clock,
  input         reset,
  input  [31:0] io_src1,
  input  [31:0] io_src2,
  input         io_signed,
  input         io_start,
  output [63:0] io_result,
  output        io_ready
);
  wire  MulBlackBox_clk; // @[Mul.scala 33:19]
  wire  MulBlackBox_rst; // @[Mul.scala 33:19]
  wire [31:0] MulBlackBox_a; // @[Mul.scala 33:19]
  wire [31:0] MulBlackBox_b; // @[Mul.scala 33:19]
  wire  MulBlackBox_sign; // @[Mul.scala 33:19]
  wire  MulBlackBox_start; // @[Mul.scala 33:19]
  wire [63:0] MulBlackBox_result; // @[Mul.scala 33:19]
  wire  MulBlackBox_ready; // @[Mul.scala 33:19]
  MulBlackBox MulBlackBox ( // @[Mul.scala 33:19]
    .clk(MulBlackBox_clk),
    .rst(MulBlackBox_rst),
    .a(MulBlackBox_a),
    .b(MulBlackBox_b),
    .sign(MulBlackBox_sign),
    .start(MulBlackBox_start),
    .result(MulBlackBox_result),
    .ready(MulBlackBox_ready)
  );
  assign io_result = MulBlackBox_result; // @[Mul.scala 40:13]
  assign io_ready = MulBlackBox_ready; // @[Mul.scala 41:13]
  assign MulBlackBox_clk = clock; // @[Mul.scala 34:13]
  assign MulBlackBox_rst = reset; // @[Mul.scala 35:13]
  assign MulBlackBox_a = io_src1; // @[Mul.scala 36:13]
  assign MulBlackBox_b = io_src2; // @[Mul.scala 37:13]
  assign MulBlackBox_sign = io_signed; // @[Mul.scala 38:13]
  assign MulBlackBox_start = io_start; // @[Mul.scala 39:13]
endmodule
module Div(
  input         clock,
  input         reset,
  input  [31:0] io_src1,
  input  [31:0] io_src2,
  input         io_signed,
  input         io_start,
  output        io_ready,
  output [63:0] io_result
);
  wire  DivBlackBox_clk; // @[Div.scala 37:19]
  wire  DivBlackBox_rst; // @[Div.scala 37:19]
  wire  DivBlackBox_signed_div_i; // @[Div.scala 37:19]
  wire  DivBlackBox_start_i; // @[Div.scala 37:19]
  wire  DivBlackBox_annul_i; // @[Div.scala 37:19]
  wire [31:0] DivBlackBox_opdata1_i; // @[Div.scala 37:19]
  wire [31:0] DivBlackBox_opdata2_i; // @[Div.scala 37:19]
  wire [63:0] DivBlackBox_result_o; // @[Div.scala 37:19]
  wire  DivBlackBox_ready_o; // @[Div.scala 37:19]
  DivBlackBox DivBlackBox ( // @[Div.scala 37:19]
    .clk(DivBlackBox_clk),
    .rst(DivBlackBox_rst),
    .signed_div_i(DivBlackBox_signed_div_i),
    .start_i(DivBlackBox_start_i),
    .annul_i(DivBlackBox_annul_i),
    .opdata1_i(DivBlackBox_opdata1_i),
    .opdata2_i(DivBlackBox_opdata2_i),
    .result_o(DivBlackBox_result_o),
    .ready_o(DivBlackBox_ready_o)
  );
  assign io_ready = DivBlackBox_ready_o; // @[Div.scala 45:20]
  assign io_result = DivBlackBox_result_o; // @[Div.scala 46:20]
  assign DivBlackBox_clk = clock; // @[Div.scala 38:20]
  assign DivBlackBox_rst = reset; // @[Div.scala 39:20]
  assign DivBlackBox_signed_div_i = io_signed; // @[Div.scala 40:20]
  assign DivBlackBox_start_i = io_start; // @[Div.scala 41:20]
  assign DivBlackBox_annul_i = 1'h0; // @[Div.scala 42:20]
  assign DivBlackBox_opdata1_i = io_src1; // @[Div.scala 43:20]
  assign DivBlackBox_opdata2_i = io_src2; // @[Div.scala 44:20]
endmodule
module HiLo(
  input         clock,
  input         reset,
  input         io_wen,
  input  [63:0] io_wdata,
  output [63:0] io_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] hilo; // @[HiLo.scala 15:21]
  assign io_rdata = hilo; // @[HiLo.scala 21:12]
  always @(posedge clock) begin
    if (reset) begin // @[HiLo.scala 15:21]
      hilo <= 64'h0; // @[HiLo.scala 15:21]
    end else if (io_wen) begin // @[HiLo.scala 17:16]
      hilo <= io_wdata; // @[HiLo.scala 18:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  hilo = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BranchCtrl(
  input  [6:0]  io_in_inst_info_op,
  input  [31:0] io_in_src_info_src1_data,
  input  [31:0] io_in_src_info_src2_data,
  input         io_in_pred_branch_flag,
  output        io_out_branch_flag,
  output        io_out_pred_fail
);
  wire  _io_out_branch_flag_T = io_in_src_info_src1_data == io_in_src_info_src2_data; // @[BranchCtrl.scala 27:27]
  wire  _io_out_branch_flag_T_1 = io_in_src_info_src1_data != io_in_src_info_src2_data; // @[BranchCtrl.scala 28:27]
  wire  _io_out_branch_flag_T_3 = ~io_in_src_info_src1_data[31]; // @[BranchCtrl.scala 29:22]
  wire  _io_out_branch_flag_T_5 = ~io_in_src_info_src1_data[31] & io_in_src_info_src1_data != 32'h0; // @[BranchCtrl.scala 29:32]
  wire  _io_out_branch_flag_T_8 = io_in_src_info_src1_data[31] | io_in_src_info_src1_data == 32'h0; // @[BranchCtrl.scala 30:31]
  wire  _io_out_branch_flag_T_18 = 7'h2f == io_in_inst_info_op ? _io_out_branch_flag_T_1 : 7'h28 == io_in_inst_info_op
     & _io_out_branch_flag_T; // @[Mux.scala 81:58]
  wire  _io_out_branch_flag_T_20 = 7'h2b == io_in_inst_info_op ? _io_out_branch_flag_T_5 : _io_out_branch_flag_T_18; // @[Mux.scala 81:58]
  wire  _io_out_branch_flag_T_22 = 7'h2c == io_in_inst_info_op ? _io_out_branch_flag_T_8 : _io_out_branch_flag_T_20; // @[Mux.scala 81:58]
  wire  _io_out_branch_flag_T_24 = 7'h29 == io_in_inst_info_op ? _io_out_branch_flag_T_3 : _io_out_branch_flag_T_22; // @[Mux.scala 81:58]
  wire  _io_out_branch_flag_T_26 = 7'h2a == io_in_inst_info_op ? _io_out_branch_flag_T_3 : _io_out_branch_flag_T_24; // @[Mux.scala 81:58]
  wire  _io_out_branch_flag_T_28 = 7'h2d == io_in_inst_info_op ? io_in_src_info_src1_data[31] : _io_out_branch_flag_T_26
    ; // @[Mux.scala 81:58]
  assign io_out_branch_flag = 7'h2e == io_in_inst_info_op ? io_in_src_info_src1_data[31] : _io_out_branch_flag_T_28; // @[Mux.scala 81:58]
  assign io_out_pred_fail = io_in_pred_branch_flag != io_out_branch_flag; // @[BranchCtrl.scala 22:46]
endmodule
module Fu(
  input         clock,
  input         reset,
  input         io_ctrl_allow_to_go,
  input         io_ctrl_do_flush,
  input  [31:0] io_inst_0_pc,
  input         io_inst_0_hilo_wen,
  input         io_inst_0_mul_en,
  input         io_inst_0_div_en,
  input  [6:0]  io_inst_0_inst_info_op,
  input  [31:0] io_inst_0_src_info_src1_data,
  input  [31:0] io_inst_0_src_info_src2_data,
  input         io_inst_0_ex_in_flush_req,
  input         io_inst_0_ex_in_eret,
  input  [31:0] io_inst_0_ex_in_badvaddr,
  input         io_inst_0_ex_in_bd,
  input  [4:0]  io_inst_0_ex_in_excode,
  output        io_inst_0_ex_out_flush_req,
  output        io_inst_0_ex_out_eret,
  output [31:0] io_inst_0_ex_out_badvaddr,
  output        io_inst_0_ex_out_bd,
  output [4:0]  io_inst_0_ex_out_excode,
  output [31:0] io_inst_0_result,
  input         io_inst_1_hilo_wen,
  input         io_inst_1_mul_en,
  input         io_inst_1_div_en,
  input  [6:0]  io_inst_1_inst_info_op,
  input  [31:0] io_inst_1_src_info_src1_data,
  input  [31:0] io_inst_1_src_info_src2_data,
  input         io_inst_1_ex_in_flush_req,
  input         io_inst_1_ex_in_eret,
  input  [31:0] io_inst_1_ex_in_badvaddr,
  input         io_inst_1_ex_in_bd,
  input  [4:0]  io_inst_1_ex_in_excode,
  output        io_inst_1_ex_out_flush_req,
  output        io_inst_1_ex_out_eret,
  output [31:0] io_inst_1_ex_out_badvaddr,
  output        io_inst_1_ex_out_bd,
  output [4:0]  io_inst_1_ex_out_excode,
  output [31:0] io_inst_1_result,
  input  [31:0] io_cp0_rdata,
  output        io_stall_req,
  input         io_branch_pred_branch_flag,
  output        io_branch_branch_flag,
  output        io_branch_pred_fail
);
  wire [6:0] alu_0_io_inst_info_op; // @[Fu.scala 40:54]
  wire [31:0] alu_0_io_src_info_src1_data; // @[Fu.scala 40:54]
  wire [31:0] alu_0_io_src_info_src2_data; // @[Fu.scala 40:54]
  wire [31:0] alu_0_io_cp0_rdata; // @[Fu.scala 40:54]
  wire [63:0] alu_0_io_hilo_rdata; // @[Fu.scala 40:54]
  wire [63:0] alu_0_io_hilo_wdata; // @[Fu.scala 40:54]
  wire  alu_0_io_mul_ready; // @[Fu.scala 40:54]
  wire [63:0] alu_0_io_mul_result; // @[Fu.scala 40:54]
  wire  alu_0_io_mul_start; // @[Fu.scala 40:54]
  wire  alu_0_io_mul_signed; // @[Fu.scala 40:54]
  wire  alu_0_io_div_ready; // @[Fu.scala 40:54]
  wire [63:0] alu_0_io_div_result; // @[Fu.scala 40:54]
  wire  alu_0_io_div_start; // @[Fu.scala 40:54]
  wire  alu_0_io_div_signed; // @[Fu.scala 40:54]
  wire [31:0] alu_0_io_result; // @[Fu.scala 40:54]
  wire  alu_0_io_overflow; // @[Fu.scala 40:54]
  wire [6:0] alu_1_io_inst_info_op; // @[Fu.scala 40:54]
  wire [31:0] alu_1_io_src_info_src1_data; // @[Fu.scala 40:54]
  wire [31:0] alu_1_io_src_info_src2_data; // @[Fu.scala 40:54]
  wire [31:0] alu_1_io_cp0_rdata; // @[Fu.scala 40:54]
  wire [63:0] alu_1_io_hilo_rdata; // @[Fu.scala 40:54]
  wire [63:0] alu_1_io_hilo_wdata; // @[Fu.scala 40:54]
  wire  alu_1_io_mul_ready; // @[Fu.scala 40:54]
  wire [63:0] alu_1_io_mul_result; // @[Fu.scala 40:54]
  wire  alu_1_io_mul_start; // @[Fu.scala 40:54]
  wire  alu_1_io_mul_signed; // @[Fu.scala 40:54]
  wire  alu_1_io_div_ready; // @[Fu.scala 40:54]
  wire [63:0] alu_1_io_div_result; // @[Fu.scala 40:54]
  wire  alu_1_io_div_start; // @[Fu.scala 40:54]
  wire  alu_1_io_div_signed; // @[Fu.scala 40:54]
  wire [31:0] alu_1_io_result; // @[Fu.scala 40:54]
  wire  alu_1_io_overflow; // @[Fu.scala 40:54]
  wire  Mul_clock; // @[Fu.scala 41:26]
  wire  Mul_reset; // @[Fu.scala 41:26]
  wire [31:0] Mul_io_src1; // @[Fu.scala 41:26]
  wire [31:0] Mul_io_src2; // @[Fu.scala 41:26]
  wire  Mul_io_signed; // @[Fu.scala 41:26]
  wire  Mul_io_start; // @[Fu.scala 41:26]
  wire [63:0] Mul_io_result; // @[Fu.scala 41:26]
  wire  Mul_io_ready; // @[Fu.scala 41:26]
  wire  Div_clock; // @[Fu.scala 42:26]
  wire  Div_reset; // @[Fu.scala 42:26]
  wire [31:0] Div_io_src1; // @[Fu.scala 42:26]
  wire [31:0] Div_io_src2; // @[Fu.scala 42:26]
  wire  Div_io_signed; // @[Fu.scala 42:26]
  wire  Div_io_start; // @[Fu.scala 42:26]
  wire  Div_io_ready; // @[Fu.scala 42:26]
  wire [63:0] Div_io_result; // @[Fu.scala 42:26]
  wire  HiLo_clock; // @[Fu.scala 43:26]
  wire  HiLo_reset; // @[Fu.scala 43:26]
  wire  HiLo_io_wen; // @[Fu.scala 43:26]
  wire [63:0] HiLo_io_wdata; // @[Fu.scala 43:26]
  wire [63:0] HiLo_io_rdata; // @[Fu.scala 43:26]
  wire [6:0] BranchCtrl_io_in_inst_info_op; // @[Fu.scala 44:26]
  wire [31:0] BranchCtrl_io_in_src_info_src1_data; // @[Fu.scala 44:26]
  wire [31:0] BranchCtrl_io_in_src_info_src2_data; // @[Fu.scala 44:26]
  wire  BranchCtrl_io_in_pred_branch_flag; // @[Fu.scala 44:26]
  wire  BranchCtrl_io_out_branch_flag; // @[Fu.scala 44:26]
  wire  BranchCtrl_io_out_pred_fail; // @[Fu.scala 44:26]
  wire  _io_inst_0_ex_out_excode_T = io_inst_0_ex_in_excode != 5'h0; // @[Fu.scala 65:34]
  wire [4:0] _io_inst_0_ex_out_excode_T_1 = alu_0_io_overflow ? 5'hb : io_inst_0_ex_in_excode; // @[Mux.scala 101:16]
  wire  _io_inst_1_ex_out_excode_T = io_inst_1_ex_in_excode != 5'h0; // @[Fu.scala 65:34]
  wire [4:0] _io_inst_1_ex_out_excode_T_1 = alu_1_io_overflow ? 5'hb : io_inst_1_ex_in_excode; // @[Mux.scala 101:16]
  wire  _io_stall_req_T_5 = (io_inst_0_div_en | io_inst_1_div_en) & ~Div_io_ready; // @[Fu.scala 85:43]
  wire  _io_inst_0_result_T_7 = 7'h25 == io_inst_0_inst_info_op | 7'h26 == io_inst_0_inst_info_op | 7'h2a ==
    io_inst_0_inst_info_op | 7'h2e == io_inst_0_inst_info_op; // @[Fu.scala 88:64]
  wire [31:0] _io_inst_0_result_T_9 = io_inst_0_pc + 32'h8; // @[Fu.scala 89:19]
  wire  _T_12 = io_inst_1_hilo_wen & ~io_inst_1_ex_out_flush_req; // @[Fu.scala 95:26]
  wire  _T_13 = io_inst_0_hilo_wen & ~(io_inst_0_ex_out_flush_req | io_inst_1_ex_out_flush_req) | _T_12; // @[Fu.scala 94:89]
  Alu alu_0 ( // @[Fu.scala 40:54]
    .io_inst_info_op(alu_0_io_inst_info_op),
    .io_src_info_src1_data(alu_0_io_src_info_src1_data),
    .io_src_info_src2_data(alu_0_io_src_info_src2_data),
    .io_cp0_rdata(alu_0_io_cp0_rdata),
    .io_hilo_rdata(alu_0_io_hilo_rdata),
    .io_hilo_wdata(alu_0_io_hilo_wdata),
    .io_mul_ready(alu_0_io_mul_ready),
    .io_mul_result(alu_0_io_mul_result),
    .io_mul_start(alu_0_io_mul_start),
    .io_mul_signed(alu_0_io_mul_signed),
    .io_div_ready(alu_0_io_div_ready),
    .io_div_result(alu_0_io_div_result),
    .io_div_start(alu_0_io_div_start),
    .io_div_signed(alu_0_io_div_signed),
    .io_result(alu_0_io_result),
    .io_overflow(alu_0_io_overflow)
  );
  Alu alu_1 ( // @[Fu.scala 40:54]
    .io_inst_info_op(alu_1_io_inst_info_op),
    .io_src_info_src1_data(alu_1_io_src_info_src1_data),
    .io_src_info_src2_data(alu_1_io_src_info_src2_data),
    .io_cp0_rdata(alu_1_io_cp0_rdata),
    .io_hilo_rdata(alu_1_io_hilo_rdata),
    .io_hilo_wdata(alu_1_io_hilo_wdata),
    .io_mul_ready(alu_1_io_mul_ready),
    .io_mul_result(alu_1_io_mul_result),
    .io_mul_start(alu_1_io_mul_start),
    .io_mul_signed(alu_1_io_mul_signed),
    .io_div_ready(alu_1_io_div_ready),
    .io_div_result(alu_1_io_div_result),
    .io_div_start(alu_1_io_div_start),
    .io_div_signed(alu_1_io_div_signed),
    .io_result(alu_1_io_result),
    .io_overflow(alu_1_io_overflow)
  );
  Mul Mul ( // @[Fu.scala 41:26]
    .clock(Mul_clock),
    .reset(Mul_reset),
    .io_src1(Mul_io_src1),
    .io_src2(Mul_io_src2),
    .io_signed(Mul_io_signed),
    .io_start(Mul_io_start),
    .io_result(Mul_io_result),
    .io_ready(Mul_io_ready)
  );
  Div Div ( // @[Fu.scala 42:26]
    .clock(Div_clock),
    .reset(Div_reset),
    .io_src1(Div_io_src1),
    .io_src2(Div_io_src2),
    .io_signed(Div_io_signed),
    .io_start(Div_io_start),
    .io_ready(Div_io_ready),
    .io_result(Div_io_result)
  );
  HiLo HiLo ( // @[Fu.scala 43:26]
    .clock(HiLo_clock),
    .reset(HiLo_reset),
    .io_wen(HiLo_io_wen),
    .io_wdata(HiLo_io_wdata),
    .io_rdata(HiLo_io_rdata)
  );
  BranchCtrl BranchCtrl ( // @[Fu.scala 44:26]
    .io_in_inst_info_op(BranchCtrl_io_in_inst_info_op),
    .io_in_src_info_src1_data(BranchCtrl_io_in_src_info_src1_data),
    .io_in_src_info_src2_data(BranchCtrl_io_in_src_info_src2_data),
    .io_in_pred_branch_flag(BranchCtrl_io_in_pred_branch_flag),
    .io_out_branch_flag(BranchCtrl_io_out_branch_flag),
    .io_out_pred_fail(BranchCtrl_io_out_pred_fail)
  );
  assign io_inst_0_ex_out_flush_req = io_inst_0_ex_in_flush_req | alu_0_io_overflow; // @[Fu.scala 61:63]
  assign io_inst_0_ex_out_eret = io_inst_0_ex_in_eret; // @[Fu.scala 60:33]
  assign io_inst_0_ex_out_badvaddr = io_inst_0_ex_in_badvaddr; // @[Fu.scala 60:33]
  assign io_inst_0_ex_out_bd = io_inst_0_ex_in_bd; // @[Fu.scala 60:33]
  assign io_inst_0_ex_out_excode = _io_inst_0_ex_out_excode_T ? io_inst_0_ex_in_excode : _io_inst_0_ex_out_excode_T_1; // @[Mux.scala 101:16]
  assign io_inst_0_result = _io_inst_0_result_T_7 ? _io_inst_0_result_T_9 : alu_0_io_result; // @[Fu.scala 87:27]
  assign io_inst_1_ex_out_flush_req = io_inst_1_ex_in_flush_req | alu_1_io_overflow; // @[Fu.scala 61:63]
  assign io_inst_1_ex_out_eret = io_inst_1_ex_in_eret; // @[Fu.scala 60:33]
  assign io_inst_1_ex_out_badvaddr = io_inst_1_ex_in_badvaddr; // @[Fu.scala 60:33]
  assign io_inst_1_ex_out_bd = io_inst_1_ex_in_bd; // @[Fu.scala 60:33]
  assign io_inst_1_ex_out_excode = _io_inst_1_ex_out_excode_T ? io_inst_1_ex_in_excode : _io_inst_1_ex_out_excode_T_1; // @[Mux.scala 101:16]
  assign io_inst_1_result = alu_1_io_result; // @[Fu.scala 92:21]
  assign io_stall_req = (io_inst_0_mul_en | io_inst_1_mul_en) & ~Mul_io_ready | _io_stall_req_T_5; // @[Fu.scala 84:72]
  assign io_branch_branch_flag = BranchCtrl_io_out_branch_flag; // @[Fu.scala 49:34]
  assign io_branch_pred_fail = BranchCtrl_io_out_pred_fail; // @[Fu.scala 50:34]
  assign alu_0_io_inst_info_op = io_inst_0_inst_info_op; // @[Fu.scala 53:33]
  assign alu_0_io_src_info_src1_data = io_inst_0_src_info_src1_data; // @[Fu.scala 54:33]
  assign alu_0_io_src_info_src2_data = io_inst_0_src_info_src2_data; // @[Fu.scala 54:33]
  assign alu_0_io_cp0_rdata = io_cp0_rdata; // @[Fu.scala 70:23]
  assign alu_0_io_hilo_rdata = HiLo_io_rdata; // @[Fu.scala 55:33]
  assign alu_0_io_mul_ready = Mul_io_ready; // @[Fu.scala 56:33]
  assign alu_0_io_mul_result = Mul_io_result; // @[Fu.scala 57:33]
  assign alu_0_io_div_ready = Div_io_ready; // @[Fu.scala 58:33]
  assign alu_0_io_div_result = Div_io_result; // @[Fu.scala 59:33]
  assign alu_1_io_inst_info_op = io_inst_1_inst_info_op; // @[Fu.scala 53:33]
  assign alu_1_io_src_info_src1_data = io_inst_1_src_info_src1_data; // @[Fu.scala 54:33]
  assign alu_1_io_src_info_src2_data = io_inst_1_src_info_src2_data; // @[Fu.scala 54:33]
  assign alu_1_io_cp0_rdata = 32'h0; // @[Fu.scala 71:23]
  assign alu_1_io_hilo_rdata = HiLo_io_rdata; // @[Fu.scala 55:33]
  assign alu_1_io_mul_ready = Mul_io_ready; // @[Fu.scala 56:33]
  assign alu_1_io_mul_result = Mul_io_result; // @[Fu.scala 57:33]
  assign alu_1_io_div_ready = Div_io_ready; // @[Fu.scala 58:33]
  assign alu_1_io_div_result = Div_io_result; // @[Fu.scala 59:33]
  assign Mul_clock = clock;
  assign Mul_reset = reset;
  assign Mul_io_src1 = io_inst_0_mul_en ? io_inst_0_src_info_src1_data : io_inst_1_src_info_src1_data; // @[Fu.scala 73:20]
  assign Mul_io_src2 = io_inst_0_mul_en ? io_inst_0_src_info_src2_data : io_inst_1_src_info_src2_data; // @[Fu.scala 74:20]
  assign Mul_io_signed = io_inst_0_mul_en ? alu_0_io_mul_signed : alu_1_io_mul_signed; // @[Fu.scala 75:20]
  assign Mul_io_start = io_inst_0_mul_en ? alu_0_io_mul_start : alu_1_io_mul_start; // @[Fu.scala 76:20]
  assign Div_clock = clock;
  assign Div_reset = reset;
  assign Div_io_src1 = io_inst_0_div_en ? io_inst_0_src_info_src1_data : io_inst_1_src_info_src1_data; // @[Fu.scala 78:20]
  assign Div_io_src2 = io_inst_0_div_en ? io_inst_0_src_info_src2_data : io_inst_1_src_info_src2_data; // @[Fu.scala 79:20]
  assign Div_io_signed = io_inst_0_div_en ? alu_0_io_div_signed : alu_1_io_div_signed; // @[Fu.scala 80:20]
  assign Div_io_start = io_inst_0_div_en ? alu_0_io_div_start : alu_1_io_div_start; // @[Fu.scala 81:20]
  assign HiLo_clock = clock;
  assign HiLo_reset = reset;
  assign HiLo_io_wen = _T_13 & io_ctrl_allow_to_go & ~io_ctrl_do_flush; // @[Fu.scala 95:83]
  assign HiLo_io_wdata = io_inst_1_hilo_wen ? alu_1_io_hilo_wdata : alu_0_io_hilo_wdata; // @[Fu.scala 96:20]
  assign BranchCtrl_io_in_inst_info_op = io_inst_0_inst_info_op; // @[Fu.scala 46:34]
  assign BranchCtrl_io_in_src_info_src1_data = io_inst_0_src_info_src1_data; // @[Fu.scala 47:34]
  assign BranchCtrl_io_in_src_info_src2_data = io_inst_0_src_info_src2_data; // @[Fu.scala 47:34]
  assign BranchCtrl_io_in_pred_branch_flag = io_branch_pred_branch_flag; // @[Fu.scala 48:34]
endmodule
module ExeAccessMemCtrl(
  output        io_mem_out_en,
  output [6:0]  io_mem_out_inst_info_op,
  output [31:0] io_mem_out_addr,
  output [31:0] io_mem_out_wdata,
  input  [3:0]  io_inst_0_inst_info_fusel,
  input  [6:0]  io_inst_0_inst_info_op,
  input  [31:0] io_inst_0_inst_info_inst,
  input  [31:0] io_inst_0_src_info_src1_data,
  input  [31:0] io_inst_0_src_info_src2_data,
  input         io_inst_0_ex_in_flush_req,
  input         io_inst_0_ex_in_eret,
  input  [31:0] io_inst_0_ex_in_badvaddr,
  input         io_inst_0_ex_in_bd,
  input  [4:0]  io_inst_0_ex_in_excode,
  output        io_inst_0_ex_out_flush_req,
  output        io_inst_0_ex_out_eret,
  output [31:0] io_inst_0_ex_out_badvaddr,
  output        io_inst_0_ex_out_bd,
  output [4:0]  io_inst_0_ex_out_excode,
  output        io_inst_0_mem_sel,
  input  [3:0]  io_inst_1_inst_info_fusel,
  input  [6:0]  io_inst_1_inst_info_op,
  input  [31:0] io_inst_1_inst_info_inst,
  input  [31:0] io_inst_1_src_info_src1_data,
  input  [31:0] io_inst_1_src_info_src2_data,
  input         io_inst_1_ex_in_flush_req,
  input         io_inst_1_ex_in_eret,
  input  [31:0] io_inst_1_ex_in_badvaddr,
  input         io_inst_1_ex_in_bd,
  input  [4:0]  io_inst_1_ex_in_excode,
  output        io_inst_1_ex_out_flush_req,
  output        io_inst_1_ex_out_eret,
  output [31:0] io_inst_1_ex_out_badvaddr,
  output        io_inst_1_ex_out_bd,
  output [4:0]  io_inst_1_ex_out_excode,
  output        io_inst_1_mem_sel
);
  wire  _io_mem_out_inst_info_T = io_inst_0_inst_info_fusel == 4'h4; // @[ExeAccessMemCtrl.scala 43:35]
  wire  _io_mem_out_inst_info_T_1 = io_inst_1_inst_info_fusel == 4'h4; // @[ExeAccessMemCtrl.scala 44:35]
  wire [6:0] _io_mem_out_inst_info_T_2_op = _io_mem_out_inst_info_T_1 ? io_inst_1_inst_info_op : 7'h0; // @[Mux.scala 101:16]
  wire [15:0] _mem_addr_0_T_3 = io_inst_0_inst_info_inst[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _mem_addr_0_T_4 = {_mem_addr_0_T_3,io_inst_0_inst_info_inst[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] mem_addr_0 = io_inst_0_src_info_src1_data + _mem_addr_0_T_4; // @[ExeAccessMemCtrl.scala 48:48]
  wire [15:0] _mem_addr_1_T_3 = io_inst_1_inst_info_inst[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _mem_addr_1_T_4 = {_mem_addr_1_T_3,io_inst_1_inst_info_inst[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] mem_addr_1 = io_inst_1_src_info_src1_data + _mem_addr_1_T_4; // @[ExeAccessMemCtrl.scala 49:48]
  wire [31:0] _io_mem_out_addr_T_2 = _io_mem_out_inst_info_T_1 ? mem_addr_1 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _io_mem_out_wdata_T_2 = _io_mem_out_inst_info_T_1 ? io_inst_1_src_info_src2_data : 32'h0; // @[Mux.scala 101:16]
  wire  _mem_adel_0_T_5 = mem_addr_0[1:0] != 2'h0; // @[ExeAccessMemCtrl.scala 68:99]
  wire  _mem_adel_0_T_13 = (7'h32 == io_inst_0_inst_info_op | 7'h33 == io_inst_0_inst_info_op) & mem_addr_0[0]; // @[ExeAccessMemCtrl.scala 69:66]
  wire  mem_adel_0 = (7'h35 == io_inst_0_inst_info_op | 7'h34 == io_inst_0_inst_info_op) & mem_addr_0[1:0] != 2'h0 |
    _mem_adel_0_T_13; // @[ExeAccessMemCtrl.scala 68:107]
  wire  _mem_adel_1_T_5 = mem_addr_1[1:0] != 2'h0; // @[ExeAccessMemCtrl.scala 68:99]
  wire  _mem_adel_1_T_13 = (7'h32 == io_inst_1_inst_info_op | 7'h33 == io_inst_1_inst_info_op) & mem_addr_1[0]; // @[ExeAccessMemCtrl.scala 69:66]
  wire  mem_adel_1 = (7'h35 == io_inst_1_inst_info_op | 7'h34 == io_inst_1_inst_info_op) & mem_addr_1[1:0] != 2'h0 |
    _mem_adel_1_T_13; // @[ExeAccessMemCtrl.scala 68:107]
  wire  _mem_ades_0_T_10 = io_inst_0_inst_info_op == 7'h3a & mem_addr_0[0]; // @[ExeAccessMemCtrl.scala 74:42]
  wire  mem_ades_0 = (7'h3b == io_inst_0_inst_info_op | 7'h39 == io_inst_0_inst_info_op) & _mem_adel_0_T_5 |
    _mem_ades_0_T_10; // @[ExeAccessMemCtrl.scala 73:107]
  wire  _mem_ades_1_T_10 = io_inst_1_inst_info_op == 7'h3a & mem_addr_1[0]; // @[ExeAccessMemCtrl.scala 74:42]
  wire  mem_ades_1 = (7'h3b == io_inst_1_inst_info_op | 7'h39 == io_inst_1_inst_info_op) & _mem_adel_1_T_5 |
    _mem_ades_1_T_10; // @[ExeAccessMemCtrl.scala 73:107]
  wire  _io_inst_0_ex_out_excode_T = io_inst_0_ex_in_excode != 5'h0; // @[ExeAccessMemCtrl.scala 82:34]
  wire [4:0] _io_inst_0_ex_out_excode_T_1 = mem_ades_0 ? 5'h6 : io_inst_0_ex_in_excode; // @[Mux.scala 101:16]
  wire [4:0] _io_inst_0_ex_out_excode_T_2 = mem_adel_0 ? 5'h5 : _io_inst_0_ex_out_excode_T_1; // @[Mux.scala 101:16]
  wire  _io_inst_0_ex_out_badvaddr_T_3 = 5'h5 == io_inst_0_ex_in_excode | 5'h6 == io_inst_0_ex_in_excode; // @[ExeAccessMemCtrl.scala 88:41]
  wire  _io_inst_1_ex_out_excode_T = io_inst_1_ex_in_excode != 5'h0; // @[ExeAccessMemCtrl.scala 82:34]
  wire [4:0] _io_inst_1_ex_out_excode_T_1 = mem_ades_1 ? 5'h6 : io_inst_1_ex_in_excode; // @[Mux.scala 101:16]
  wire [4:0] _io_inst_1_ex_out_excode_T_2 = mem_adel_1 ? 5'h5 : _io_inst_1_ex_out_excode_T_1; // @[Mux.scala 101:16]
  wire  _io_inst_1_ex_out_badvaddr_T_3 = 5'h5 == io_inst_1_ex_in_excode | 5'h6 == io_inst_1_ex_in_excode; // @[ExeAccessMemCtrl.scala 88:41]
  wire  _io_inst_0_mem_sel_T_1 = ~io_inst_0_ex_out_flush_req; // @[ExeAccessMemCtrl.scala 95:5]
  wire  _io_inst_1_mem_sel_T_2 = _io_mem_out_inst_info_T_1 & _io_inst_0_mem_sel_T_1; // @[ExeAccessMemCtrl.scala 96:63]
  assign io_mem_out_en = io_inst_0_mem_sel | io_inst_1_mem_sel; // @[ExeAccessMemCtrl.scala 35:52]
  assign io_mem_out_inst_info_op = _io_mem_out_inst_info_T ? io_inst_0_inst_info_op : _io_mem_out_inst_info_T_2_op; // @[Mux.scala 101:16]
  assign io_mem_out_addr = _io_mem_out_inst_info_T ? mem_addr_0 : _io_mem_out_addr_T_2; // @[Mux.scala 101:16]
  assign io_mem_out_wdata = _io_mem_out_inst_info_T ? io_inst_0_src_info_src2_data : _io_mem_out_wdata_T_2; // @[Mux.scala 101:16]
  assign io_inst_0_ex_out_flush_req = io_inst_0_ex_in_flush_req | io_inst_0_ex_out_excode != 5'h0; // @[ExeAccessMemCtrl.scala 92:63]
  assign io_inst_0_ex_out_eret = io_inst_0_ex_in_eret; // @[ExeAccessMemCtrl.scala 78:23]
  assign io_inst_0_ex_out_badvaddr = _io_inst_0_ex_out_badvaddr_T_3 ? io_inst_0_ex_in_badvaddr : mem_addr_0; // @[ExeAccessMemCtrl.scala 87:38]
  assign io_inst_0_ex_out_bd = io_inst_0_ex_in_bd; // @[ExeAccessMemCtrl.scala 78:23]
  assign io_inst_0_ex_out_excode = _io_inst_0_ex_out_excode_T ? io_inst_0_ex_in_excode : _io_inst_0_ex_out_excode_T_2; // @[Mux.scala 101:16]
  assign io_inst_0_mem_sel = _io_mem_out_inst_info_T & _io_inst_0_mem_sel_T_1; // @[ExeAccessMemCtrl.scala 94:63]
  assign io_inst_1_ex_out_flush_req = io_inst_1_ex_in_flush_req | io_inst_1_ex_out_excode != 5'h0; // @[ExeAccessMemCtrl.scala 92:63]
  assign io_inst_1_ex_out_eret = io_inst_1_ex_in_eret; // @[ExeAccessMemCtrl.scala 78:23]
  assign io_inst_1_ex_out_badvaddr = _io_inst_1_ex_out_badvaddr_T_3 ? io_inst_1_ex_in_badvaddr : mem_addr_1; // @[ExeAccessMemCtrl.scala 87:38]
  assign io_inst_1_ex_out_bd = io_inst_1_ex_in_bd; // @[ExeAccessMemCtrl.scala 78:23]
  assign io_inst_1_ex_out_excode = _io_inst_1_ex_out_excode_T ? io_inst_1_ex_in_excode : _io_inst_1_ex_out_excode_T_2; // @[Mux.scala 101:16]
  assign io_inst_1_mem_sel = _io_inst_1_mem_sel_T_2 & ~io_inst_1_ex_out_flush_req; // @[ExeAccessMemCtrl.scala 97:34]
endmodule
module ExecuteUnit(
  input         clock,
  input         reset,
  output        io_ctrl_inst_0_mem_ren,
  output [4:0]  io_ctrl_inst_0_reg_waddr,
  output        io_ctrl_inst_1_mem_ren,
  output [4:0]  io_ctrl_inst_1_reg_waddr,
  output        io_ctrl_fu_stall,
  output        io_ctrl_branch_flag,
  input         io_ctrl_allow_to_go,
  input         io_ctrl_fu_allow_to_go,
  input         io_ctrl_fu_do_flush,
  input  [31:0] io_executeStage_inst0_pc,
  input  [3:0]  io_executeStage_inst0_inst_info_fusel,
  input  [6:0]  io_executeStage_inst0_inst_info_op,
  input         io_executeStage_inst0_inst_info_reg_wen,
  input  [4:0]  io_executeStage_inst0_inst_info_reg_waddr,
  input  [7:0]  io_executeStage_inst0_inst_info_cp0_addr,
  input  [31:0] io_executeStage_inst0_inst_info_inst,
  input  [31:0] io_executeStage_inst0_src_info_src1_data,
  input  [31:0] io_executeStage_inst0_src_info_src2_data,
  input         io_executeStage_inst0_ex_flush_req,
  input         io_executeStage_inst0_ex_eret,
  input  [31:0] io_executeStage_inst0_ex_badvaddr,
  input         io_executeStage_inst0_ex_bd,
  input  [4:0]  io_executeStage_inst0_ex_excode,
  input         io_executeStage_inst0_jb_info_jump_regiser_conflict,
  input         io_executeStage_inst0_jb_info_is_branch,
  input         io_executeStage_inst0_jb_info_pred_branch_flag,
  input  [31:0] io_executeStage_inst0_jb_info_branch_target,
  input  [31:0] io_executeStage_inst1_pc,
  input  [3:0]  io_executeStage_inst1_inst_info_fusel,
  input  [6:0]  io_executeStage_inst1_inst_info_op,
  input         io_executeStage_inst1_inst_info_reg_wen,
  input  [4:0]  io_executeStage_inst1_inst_info_reg_waddr,
  input  [31:0] io_executeStage_inst1_inst_info_inst,
  input  [31:0] io_executeStage_inst1_src_info_src1_data,
  input  [31:0] io_executeStage_inst1_src_info_src2_data,
  input         io_executeStage_inst1_ex_flush_req,
  input         io_executeStage_inst1_ex_eret,
  input  [31:0] io_executeStage_inst1_ex_badvaddr,
  input         io_executeStage_inst1_ex_bd,
  input  [4:0]  io_executeStage_inst1_ex_excode,
  output [6:0]  io_cp0_in_inst_info_op,
  output [7:0]  io_cp0_in_inst_info_cp0_addr,
  output [31:0] io_cp0_in_mtc0_wdata,
  input  [31:0] io_cp0_out_cp0_rdata,
  input  [31:0] io_cp0_out_debug_cp0_count,
  input  [31:0] io_cp0_out_debug_cp0_random,
  input  [31:0] io_cp0_out_debug_cp0_cause,
  output [31:0] io_bpu_pc,
  output        io_bpu_branch_flag,
  output        io_bpu_inst0_is_branch,
  output        io_fetchStage_branch,
  output [31:0] io_fetchStage_target,
  output        io_decoderUnit_forward_0_exe_wen,
  output [4:0]  io_decoderUnit_forward_0_exe_waddr,
  output [31:0] io_decoderUnit_forward_0_exe_wdata,
  output        io_decoderUnit_forward_0_exe_mem_ren,
  output        io_decoderUnit_forward_1_exe_wen,
  output [4:0]  io_decoderUnit_forward_1_exe_waddr,
  output [31:0] io_decoderUnit_forward_1_exe_wdata,
  output        io_decoderUnit_forward_1_exe_mem_ren,
  input         io_decoderUnit_inst0_bd,
  output [31:0] io_memoryStage_inst0_pc,
  output [3:0]  io_memoryStage_inst0_inst_info_fusel,
  output [6:0]  io_memoryStage_inst0_inst_info_op,
  output        io_memoryStage_inst0_inst_info_reg_wen,
  output [4:0]  io_memoryStage_inst0_inst_info_reg_waddr,
  output [31:0] io_memoryStage_inst0_inst_info_inst,
  output [31:0] io_memoryStage_inst0_rd_info_wdata,
  output        io_memoryStage_inst0_ex_flush_req,
  output        io_memoryStage_inst0_ex_eret,
  output [31:0] io_memoryStage_inst0_ex_badvaddr,
  output        io_memoryStage_inst0_ex_bd,
  output [4:0]  io_memoryStage_inst0_ex_excode,
  output [31:0] io_memoryStage_inst0_cp0_cp0_count,
  output [31:0] io_memoryStage_inst0_cp0_cp0_random,
  output [31:0] io_memoryStage_inst0_cp0_cp0_cause,
  output        io_memoryStage_inst0_mem_en,
  output [6:0]  io_memoryStage_inst0_mem_inst_info_op,
  output [31:0] io_memoryStage_inst0_mem_addr,
  output [31:0] io_memoryStage_inst0_mem_wdata,
  output        io_memoryStage_inst0_mem_sel_0,
  output        io_memoryStage_inst0_mem_sel_1,
  output [31:0] io_memoryStage_inst1_pc,
  output [3:0]  io_memoryStage_inst1_inst_info_fusel,
  output        io_memoryStage_inst1_inst_info_reg_wen,
  output [4:0]  io_memoryStage_inst1_inst_info_reg_waddr,
  output [31:0] io_memoryStage_inst1_rd_info_wdata,
  output        io_memoryStage_inst1_ex_flush_req,
  output        io_memoryStage_inst1_ex_eret,
  output [31:0] io_memoryStage_inst1_ex_badvaddr,
  output        io_memoryStage_inst1_ex_bd,
  output [4:0]  io_memoryStage_inst1_ex_excode
);
  wire  Fu_clock; // @[ExecuteUnit.scala 40:29]
  wire  Fu_reset; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_ctrl_allow_to_go; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_ctrl_do_flush; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_0_pc; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_hilo_wen; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_mul_en; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_div_en; // @[ExecuteUnit.scala 40:29]
  wire [6:0] Fu_io_inst_0_inst_info_op; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_0_src_info_src1_data; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_0_src_info_src2_data; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_ex_in_flush_req; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_ex_in_eret; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_0_ex_in_badvaddr; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_ex_in_bd; // @[ExecuteUnit.scala 40:29]
  wire [4:0] Fu_io_inst_0_ex_in_excode; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_ex_out_flush_req; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_ex_out_eret; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_0_ex_out_badvaddr; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_0_ex_out_bd; // @[ExecuteUnit.scala 40:29]
  wire [4:0] Fu_io_inst_0_ex_out_excode; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_0_result; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_hilo_wen; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_mul_en; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_div_en; // @[ExecuteUnit.scala 40:29]
  wire [6:0] Fu_io_inst_1_inst_info_op; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_1_src_info_src1_data; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_1_src_info_src2_data; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_ex_in_flush_req; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_ex_in_eret; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_1_ex_in_badvaddr; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_ex_in_bd; // @[ExecuteUnit.scala 40:29]
  wire [4:0] Fu_io_inst_1_ex_in_excode; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_ex_out_flush_req; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_ex_out_eret; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_1_ex_out_badvaddr; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_inst_1_ex_out_bd; // @[ExecuteUnit.scala 40:29]
  wire [4:0] Fu_io_inst_1_ex_out_excode; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_inst_1_result; // @[ExecuteUnit.scala 40:29]
  wire [31:0] Fu_io_cp0_rdata; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_stall_req; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_branch_pred_branch_flag; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_branch_branch_flag; // @[ExecuteUnit.scala 40:29]
  wire  Fu_io_branch_pred_fail; // @[ExecuteUnit.scala 40:29]
  wire  ExeAccessMemCtrl_io_mem_out_en; // @[ExecuteUnit.scala 41:29]
  wire [6:0] ExeAccessMemCtrl_io_mem_out_inst_info_op; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_mem_out_addr; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_mem_out_wdata; // @[ExecuteUnit.scala 41:29]
  wire [3:0] ExeAccessMemCtrl_io_inst_0_inst_info_fusel; // @[ExecuteUnit.scala 41:29]
  wire [6:0] ExeAccessMemCtrl_io_inst_0_inst_info_op; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_0_inst_info_inst; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_0_src_info_src1_data; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_0_src_info_src2_data; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_0_ex_in_flush_req; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_0_ex_in_eret; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_0_ex_in_badvaddr; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_0_ex_in_bd; // @[ExecuteUnit.scala 41:29]
  wire [4:0] ExeAccessMemCtrl_io_inst_0_ex_in_excode; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_0_ex_out_flush_req; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_0_ex_out_eret; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_0_ex_out_badvaddr; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_0_ex_out_bd; // @[ExecuteUnit.scala 41:29]
  wire [4:0] ExeAccessMemCtrl_io_inst_0_ex_out_excode; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_0_mem_sel; // @[ExecuteUnit.scala 41:29]
  wire [3:0] ExeAccessMemCtrl_io_inst_1_inst_info_fusel; // @[ExecuteUnit.scala 41:29]
  wire [6:0] ExeAccessMemCtrl_io_inst_1_inst_info_op; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_1_inst_info_inst; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_1_src_info_src1_data; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_1_src_info_src2_data; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_1_ex_in_flush_req; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_1_ex_in_eret; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_1_ex_in_badvaddr; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_1_ex_in_bd; // @[ExecuteUnit.scala 41:29]
  wire [4:0] ExeAccessMemCtrl_io_inst_1_ex_in_excode; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_1_ex_out_flush_req; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_1_ex_out_eret; // @[ExecuteUnit.scala 41:29]
  wire [31:0] ExeAccessMemCtrl_io_inst_1_ex_out_badvaddr; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_1_ex_out_bd; // @[ExecuteUnit.scala 41:29]
  wire [4:0] ExeAccessMemCtrl_io_inst_1_ex_out_excode; // @[ExecuteUnit.scala 41:29]
  wire  ExeAccessMemCtrl_io_inst_1_mem_sel; // @[ExecuteUnit.scala 41:29]
  wire  _io_ctrl_inst_0_mem_ren_T = io_executeStage_inst0_inst_info_fusel == 4'h4; // @[ExecuteUnit.scala 43:68]
  wire  _io_ctrl_inst_1_mem_ren_T = io_executeStage_inst1_inst_info_fusel == 4'h4; // @[ExecuteUnit.scala 46:68]
  wire  _io_ctrl_branch_flag_T = io_executeStage_inst0_jb_info_jump_regiser_conflict | Fu_io_branch_pred_fail; // @[ExecuteUnit.scala 50:58]
  wire  _io_cp0_in_inst_info_T = ~io_executeStage_inst0_ex_flush_req; // @[ExecuteUnit.scala 54:5]
  wire [31:0] _io_fetchStage_target_T_1 = io_executeStage_inst0_pc + 32'h4; // @[ExecuteUnit.scala 94:30]
  wire  _io_fetchStage_target_T_2 = Fu_io_branch_pred_fail & Fu_io_branch_branch_flag; // @[ExecuteUnit.scala 96:28]
  wire  _io_fetchStage_target_T_4 = Fu_io_branch_pred_fail & ~Fu_io_branch_branch_flag; // @[ExecuteUnit.scala 97:28]
  wire  _io_fetchStage_target_T_5 = io_decoderUnit_inst0_bd | io_executeStage_inst1_ex_bd; // @[ExecuteUnit.scala 98:33]
  wire [31:0] _io_fetchStage_target_T_7 = io_executeStage_inst0_pc + 32'h8; // @[ExecuteUnit.scala 99:34]
  wire [31:0] _io_fetchStage_target_T_10 = _io_fetchStage_target_T_5 ? _io_fetchStage_target_T_7 :
    _io_fetchStage_target_T_1; // @[ExecuteUnit.scala 97:61]
  wire [31:0] _io_fetchStage_target_T_11 = io_executeStage_inst0_jb_info_jump_regiser_conflict ?
    io_executeStage_inst0_src_info_src1_data : _io_fetchStage_target_T_1; // @[Mux.scala 101:16]
  wire [31:0] _io_fetchStage_target_T_12 = _io_fetchStage_target_T_4 ? _io_fetchStage_target_T_10 :
    _io_fetchStage_target_T_11; // @[Mux.scala 101:16]
  wire  _io_memoryStage_inst0_inst_info_reg_wen_T = io_executeStage_inst0_src_info_src2_data != 32'h0; // @[ExecuteUnit.scala 122:61]
  wire  _io_memoryStage_inst0_inst_info_reg_wen_T_1 = io_executeStage_inst0_src_info_src2_data == 32'h0; // @[ExecuteUnit.scala 123:61]
  wire  _io_memoryStage_inst0_inst_info_reg_wen_T_3 = 7'hc == io_executeStage_inst0_inst_info_op ?
    _io_memoryStage_inst0_inst_info_reg_wen_T : io_executeStage_inst0_inst_info_reg_wen; // @[Mux.scala 81:58]
  wire  _io_memoryStage_inst1_inst_info_reg_wen_T = io_executeStage_inst1_src_info_src2_data != 32'h0; // @[ExecuteUnit.scala 140:61]
  wire  _io_memoryStage_inst1_inst_info_reg_wen_T_1 = io_executeStage_inst1_src_info_src2_data == 32'h0; // @[ExecuteUnit.scala 141:61]
  wire  _io_memoryStage_inst1_inst_info_reg_wen_T_3 = 7'hc == io_executeStage_inst1_inst_info_op ?
    _io_memoryStage_inst1_inst_info_reg_wen_T : io_executeStage_inst1_inst_info_reg_wen; // @[Mux.scala 81:58]
  Fu Fu ( // @[ExecuteUnit.scala 40:29]
    .clock(Fu_clock),
    .reset(Fu_reset),
    .io_ctrl_allow_to_go(Fu_io_ctrl_allow_to_go),
    .io_ctrl_do_flush(Fu_io_ctrl_do_flush),
    .io_inst_0_pc(Fu_io_inst_0_pc),
    .io_inst_0_hilo_wen(Fu_io_inst_0_hilo_wen),
    .io_inst_0_mul_en(Fu_io_inst_0_mul_en),
    .io_inst_0_div_en(Fu_io_inst_0_div_en),
    .io_inst_0_inst_info_op(Fu_io_inst_0_inst_info_op),
    .io_inst_0_src_info_src1_data(Fu_io_inst_0_src_info_src1_data),
    .io_inst_0_src_info_src2_data(Fu_io_inst_0_src_info_src2_data),
    .io_inst_0_ex_in_flush_req(Fu_io_inst_0_ex_in_flush_req),
    .io_inst_0_ex_in_eret(Fu_io_inst_0_ex_in_eret),
    .io_inst_0_ex_in_badvaddr(Fu_io_inst_0_ex_in_badvaddr),
    .io_inst_0_ex_in_bd(Fu_io_inst_0_ex_in_bd),
    .io_inst_0_ex_in_excode(Fu_io_inst_0_ex_in_excode),
    .io_inst_0_ex_out_flush_req(Fu_io_inst_0_ex_out_flush_req),
    .io_inst_0_ex_out_eret(Fu_io_inst_0_ex_out_eret),
    .io_inst_0_ex_out_badvaddr(Fu_io_inst_0_ex_out_badvaddr),
    .io_inst_0_ex_out_bd(Fu_io_inst_0_ex_out_bd),
    .io_inst_0_ex_out_excode(Fu_io_inst_0_ex_out_excode),
    .io_inst_0_result(Fu_io_inst_0_result),
    .io_inst_1_hilo_wen(Fu_io_inst_1_hilo_wen),
    .io_inst_1_mul_en(Fu_io_inst_1_mul_en),
    .io_inst_1_div_en(Fu_io_inst_1_div_en),
    .io_inst_1_inst_info_op(Fu_io_inst_1_inst_info_op),
    .io_inst_1_src_info_src1_data(Fu_io_inst_1_src_info_src1_data),
    .io_inst_1_src_info_src2_data(Fu_io_inst_1_src_info_src2_data),
    .io_inst_1_ex_in_flush_req(Fu_io_inst_1_ex_in_flush_req),
    .io_inst_1_ex_in_eret(Fu_io_inst_1_ex_in_eret),
    .io_inst_1_ex_in_badvaddr(Fu_io_inst_1_ex_in_badvaddr),
    .io_inst_1_ex_in_bd(Fu_io_inst_1_ex_in_bd),
    .io_inst_1_ex_in_excode(Fu_io_inst_1_ex_in_excode),
    .io_inst_1_ex_out_flush_req(Fu_io_inst_1_ex_out_flush_req),
    .io_inst_1_ex_out_eret(Fu_io_inst_1_ex_out_eret),
    .io_inst_1_ex_out_badvaddr(Fu_io_inst_1_ex_out_badvaddr),
    .io_inst_1_ex_out_bd(Fu_io_inst_1_ex_out_bd),
    .io_inst_1_ex_out_excode(Fu_io_inst_1_ex_out_excode),
    .io_inst_1_result(Fu_io_inst_1_result),
    .io_cp0_rdata(Fu_io_cp0_rdata),
    .io_stall_req(Fu_io_stall_req),
    .io_branch_pred_branch_flag(Fu_io_branch_pred_branch_flag),
    .io_branch_branch_flag(Fu_io_branch_branch_flag),
    .io_branch_pred_fail(Fu_io_branch_pred_fail)
  );
  ExeAccessMemCtrl ExeAccessMemCtrl ( // @[ExecuteUnit.scala 41:29]
    .io_mem_out_en(ExeAccessMemCtrl_io_mem_out_en),
    .io_mem_out_inst_info_op(ExeAccessMemCtrl_io_mem_out_inst_info_op),
    .io_mem_out_addr(ExeAccessMemCtrl_io_mem_out_addr),
    .io_mem_out_wdata(ExeAccessMemCtrl_io_mem_out_wdata),
    .io_inst_0_inst_info_fusel(ExeAccessMemCtrl_io_inst_0_inst_info_fusel),
    .io_inst_0_inst_info_op(ExeAccessMemCtrl_io_inst_0_inst_info_op),
    .io_inst_0_inst_info_inst(ExeAccessMemCtrl_io_inst_0_inst_info_inst),
    .io_inst_0_src_info_src1_data(ExeAccessMemCtrl_io_inst_0_src_info_src1_data),
    .io_inst_0_src_info_src2_data(ExeAccessMemCtrl_io_inst_0_src_info_src2_data),
    .io_inst_0_ex_in_flush_req(ExeAccessMemCtrl_io_inst_0_ex_in_flush_req),
    .io_inst_0_ex_in_eret(ExeAccessMemCtrl_io_inst_0_ex_in_eret),
    .io_inst_0_ex_in_badvaddr(ExeAccessMemCtrl_io_inst_0_ex_in_badvaddr),
    .io_inst_0_ex_in_bd(ExeAccessMemCtrl_io_inst_0_ex_in_bd),
    .io_inst_0_ex_in_excode(ExeAccessMemCtrl_io_inst_0_ex_in_excode),
    .io_inst_0_ex_out_flush_req(ExeAccessMemCtrl_io_inst_0_ex_out_flush_req),
    .io_inst_0_ex_out_eret(ExeAccessMemCtrl_io_inst_0_ex_out_eret),
    .io_inst_0_ex_out_badvaddr(ExeAccessMemCtrl_io_inst_0_ex_out_badvaddr),
    .io_inst_0_ex_out_bd(ExeAccessMemCtrl_io_inst_0_ex_out_bd),
    .io_inst_0_ex_out_excode(ExeAccessMemCtrl_io_inst_0_ex_out_excode),
    .io_inst_0_mem_sel(ExeAccessMemCtrl_io_inst_0_mem_sel),
    .io_inst_1_inst_info_fusel(ExeAccessMemCtrl_io_inst_1_inst_info_fusel),
    .io_inst_1_inst_info_op(ExeAccessMemCtrl_io_inst_1_inst_info_op),
    .io_inst_1_inst_info_inst(ExeAccessMemCtrl_io_inst_1_inst_info_inst),
    .io_inst_1_src_info_src1_data(ExeAccessMemCtrl_io_inst_1_src_info_src1_data),
    .io_inst_1_src_info_src2_data(ExeAccessMemCtrl_io_inst_1_src_info_src2_data),
    .io_inst_1_ex_in_flush_req(ExeAccessMemCtrl_io_inst_1_ex_in_flush_req),
    .io_inst_1_ex_in_eret(ExeAccessMemCtrl_io_inst_1_ex_in_eret),
    .io_inst_1_ex_in_badvaddr(ExeAccessMemCtrl_io_inst_1_ex_in_badvaddr),
    .io_inst_1_ex_in_bd(ExeAccessMemCtrl_io_inst_1_ex_in_bd),
    .io_inst_1_ex_in_excode(ExeAccessMemCtrl_io_inst_1_ex_in_excode),
    .io_inst_1_ex_out_flush_req(ExeAccessMemCtrl_io_inst_1_ex_out_flush_req),
    .io_inst_1_ex_out_eret(ExeAccessMemCtrl_io_inst_1_ex_out_eret),
    .io_inst_1_ex_out_badvaddr(ExeAccessMemCtrl_io_inst_1_ex_out_badvaddr),
    .io_inst_1_ex_out_bd(ExeAccessMemCtrl_io_inst_1_ex_out_bd),
    .io_inst_1_ex_out_excode(ExeAccessMemCtrl_io_inst_1_ex_out_excode),
    .io_inst_1_mem_sel(ExeAccessMemCtrl_io_inst_1_mem_sel)
  );
  assign io_ctrl_inst_0_mem_ren = io_executeStage_inst0_inst_info_fusel == 4'h4 &
    io_executeStage_inst0_inst_info_reg_wen; // @[ExecuteUnit.scala 43:79]
  assign io_ctrl_inst_0_reg_waddr = io_executeStage_inst0_inst_info_reg_waddr; // @[ExecuteUnit.scala 45:29]
  assign io_ctrl_inst_1_mem_ren = io_executeStage_inst1_inst_info_fusel == 4'h4 &
    io_executeStage_inst1_inst_info_reg_wen; // @[ExecuteUnit.scala 46:79]
  assign io_ctrl_inst_1_reg_waddr = io_executeStage_inst1_inst_info_reg_waddr; // @[ExecuteUnit.scala 48:29]
  assign io_ctrl_fu_stall = Fu_io_stall_req; // @[ExecuteUnit.scala 106:20]
  assign io_ctrl_branch_flag = io_ctrl_allow_to_go & _io_ctrl_branch_flag_T; // @[ExecuteUnit.scala 49:46]
  assign io_cp0_in_inst_info_op = _io_cp0_in_inst_info_T ? io_executeStage_inst0_inst_info_op : 7'h0; // @[ExecuteUnit.scala 53:29]
  assign io_cp0_in_inst_info_cp0_addr = _io_cp0_in_inst_info_T ? io_executeStage_inst0_inst_info_cp0_addr : 8'h0; // @[ExecuteUnit.scala 53:29]
  assign io_cp0_in_mtc0_wdata = io_executeStage_inst0_src_info_src2_data; // @[ExecuteUnit.scala 52:24]
  assign io_bpu_pc = io_executeStage_inst0_pc; // @[ExecuteUnit.scala 87:26]
  assign io_bpu_branch_flag = Fu_io_branch_branch_flag; // @[ExecuteUnit.scala 88:26]
  assign io_bpu_inst0_is_branch = io_executeStage_inst0_jb_info_is_branch; // @[ExecuteUnit.scala 89:26]
  assign io_fetchStage_branch = io_ctrl_allow_to_go & _io_ctrl_branch_flag_T; // @[ExecuteUnit.scala 91:47]
  assign io_fetchStage_target = _io_fetchStage_target_T_2 ? io_executeStage_inst0_jb_info_branch_target :
    _io_fetchStage_target_T_12; // @[Mux.scala 101:16]
  assign io_decoderUnit_forward_0_exe_wen = io_memoryStage_inst0_inst_info_reg_wen; // @[ExecuteUnit.scala 151:39]
  assign io_decoderUnit_forward_0_exe_waddr = io_memoryStage_inst0_inst_info_reg_waddr; // @[ExecuteUnit.scala 152:39]
  assign io_decoderUnit_forward_0_exe_wdata = io_memoryStage_inst0_rd_info_wdata; // @[ExecuteUnit.scala 153:39]
  assign io_decoderUnit_forward_0_exe_mem_ren = io_memoryStage_inst0_inst_info_fusel == 4'h4 &
    io_memoryStage_inst0_inst_info_reg_wen; // @[ExecuteUnit.scala 154:92]
  assign io_decoderUnit_forward_1_exe_wen = io_memoryStage_inst1_inst_info_reg_wen; // @[ExecuteUnit.scala 157:39]
  assign io_decoderUnit_forward_1_exe_waddr = io_memoryStage_inst1_inst_info_reg_waddr; // @[ExecuteUnit.scala 158:39]
  assign io_decoderUnit_forward_1_exe_wdata = io_memoryStage_inst1_rd_info_wdata; // @[ExecuteUnit.scala 159:39]
  assign io_decoderUnit_forward_1_exe_mem_ren = io_memoryStage_inst1_inst_info_fusel == 4'h4 &
    io_memoryStage_inst1_inst_info_reg_wen; // @[ExecuteUnit.scala 160:92]
  assign io_memoryStage_inst0_pc = io_executeStage_inst0_pc; // @[ExecuteUnit.scala 116:34]
  assign io_memoryStage_inst0_inst_info_fusel = io_executeStage_inst0_inst_info_fusel; // @[ExecuteUnit.scala 117:34]
  assign io_memoryStage_inst0_inst_info_op = io_executeStage_inst0_inst_info_op; // @[ExecuteUnit.scala 117:34]
  assign io_memoryStage_inst0_inst_info_reg_wen = 7'hb == io_executeStage_inst0_inst_info_op ?
    _io_memoryStage_inst0_inst_info_reg_wen_T_1 : _io_memoryStage_inst0_inst_info_reg_wen_T_3; // @[Mux.scala 81:58]
  assign io_memoryStage_inst0_inst_info_reg_waddr = io_executeStage_inst0_inst_info_reg_waddr; // @[ExecuteUnit.scala 117:34]
  assign io_memoryStage_inst0_inst_info_inst = io_executeStage_inst0_inst_info_inst; // @[ExecuteUnit.scala 117:34]
  assign io_memoryStage_inst0_rd_info_wdata = Fu_io_inst_0_result; // @[ExecuteUnit.scala 126:38]
  assign io_memoryStage_inst0_ex_flush_req = _io_ctrl_inst_0_mem_ren_T ? ExeAccessMemCtrl_io_inst_0_ex_out_flush_req :
    Fu_io_inst_0_ex_out_flush_req; // @[ExecuteUnit.scala 127:33]
  assign io_memoryStage_inst0_ex_eret = _io_ctrl_inst_0_mem_ren_T ? ExeAccessMemCtrl_io_inst_0_ex_out_eret :
    Fu_io_inst_0_ex_out_eret; // @[ExecuteUnit.scala 127:33]
  assign io_memoryStage_inst0_ex_badvaddr = _io_ctrl_inst_0_mem_ren_T ? ExeAccessMemCtrl_io_inst_0_ex_out_badvaddr :
    Fu_io_inst_0_ex_out_badvaddr; // @[ExecuteUnit.scala 127:33]
  assign io_memoryStage_inst0_ex_bd = _io_ctrl_inst_0_mem_ren_T ? ExeAccessMemCtrl_io_inst_0_ex_out_bd :
    Fu_io_inst_0_ex_out_bd; // @[ExecuteUnit.scala 127:33]
  assign io_memoryStage_inst0_ex_excode = _io_ctrl_inst_0_mem_ren_T ? ExeAccessMemCtrl_io_inst_0_ex_out_excode :
    Fu_io_inst_0_ex_out_excode; // @[ExecuteUnit.scala 127:33]
  assign io_memoryStage_inst0_cp0_cp0_count = io_cp0_out_debug_cp0_count; // @[ExecuteUnit.scala 132:28]
  assign io_memoryStage_inst0_cp0_cp0_random = io_cp0_out_debug_cp0_random; // @[ExecuteUnit.scala 132:28]
  assign io_memoryStage_inst0_cp0_cp0_cause = io_cp0_out_debug_cp0_cause; // @[ExecuteUnit.scala 132:28]
  assign io_memoryStage_inst0_mem_en = ExeAccessMemCtrl_io_mem_out_en; // @[ExecuteUnit.scala 108:38]
  assign io_memoryStage_inst0_mem_inst_info_op = ExeAccessMemCtrl_io_mem_out_inst_info_op; // @[ExecuteUnit.scala 114:38]
  assign io_memoryStage_inst0_mem_addr = ExeAccessMemCtrl_io_mem_out_addr; // @[ExecuteUnit.scala 111:38]
  assign io_memoryStage_inst0_mem_wdata = ExeAccessMemCtrl_io_mem_out_wdata; // @[ExecuteUnit.scala 112:38]
  assign io_memoryStage_inst0_mem_sel_0 = ExeAccessMemCtrl_io_inst_0_mem_sel; // @[ExecuteUnit.scala 113:38]
  assign io_memoryStage_inst0_mem_sel_1 = ExeAccessMemCtrl_io_inst_1_mem_sel; // @[ExecuteUnit.scala 113:38]
  assign io_memoryStage_inst1_pc = io_executeStage_inst1_pc; // @[ExecuteUnit.scala 134:34]
  assign io_memoryStage_inst1_inst_info_fusel = io_executeStage_inst1_inst_info_fusel; // @[ExecuteUnit.scala 135:34]
  assign io_memoryStage_inst1_inst_info_reg_wen = 7'hb == io_executeStage_inst1_inst_info_op ?
    _io_memoryStage_inst1_inst_info_reg_wen_T_1 : _io_memoryStage_inst1_inst_info_reg_wen_T_3; // @[Mux.scala 81:58]
  assign io_memoryStage_inst1_inst_info_reg_waddr = io_executeStage_inst1_inst_info_reg_waddr; // @[ExecuteUnit.scala 135:34]
  assign io_memoryStage_inst1_rd_info_wdata = Fu_io_inst_1_result; // @[ExecuteUnit.scala 144:38]
  assign io_memoryStage_inst1_ex_flush_req = _io_ctrl_inst_1_mem_ren_T ? ExeAccessMemCtrl_io_inst_1_ex_out_flush_req :
    Fu_io_inst_1_ex_out_flush_req; // @[ExecuteUnit.scala 145:33]
  assign io_memoryStage_inst1_ex_eret = _io_ctrl_inst_1_mem_ren_T ? ExeAccessMemCtrl_io_inst_1_ex_out_eret :
    Fu_io_inst_1_ex_out_eret; // @[ExecuteUnit.scala 145:33]
  assign io_memoryStage_inst1_ex_badvaddr = _io_ctrl_inst_1_mem_ren_T ? ExeAccessMemCtrl_io_inst_1_ex_out_badvaddr :
    Fu_io_inst_1_ex_out_badvaddr; // @[ExecuteUnit.scala 145:33]
  assign io_memoryStage_inst1_ex_bd = _io_ctrl_inst_1_mem_ren_T ? ExeAccessMemCtrl_io_inst_1_ex_out_bd :
    Fu_io_inst_1_ex_out_bd; // @[ExecuteUnit.scala 145:33]
  assign io_memoryStage_inst1_ex_excode = _io_ctrl_inst_1_mem_ren_T ? ExeAccessMemCtrl_io_inst_1_ex_out_excode :
    Fu_io_inst_1_ex_out_excode; // @[ExecuteUnit.scala 145:33]
  assign Fu_clock = clock;
  assign Fu_reset = reset;
  assign Fu_io_ctrl_allow_to_go = io_ctrl_fu_allow_to_go; // @[ExecuteUnit.scala 68:30]
  assign Fu_io_ctrl_do_flush = io_ctrl_fu_do_flush; // @[ExecuteUnit.scala 69:30]
  assign Fu_io_inst_0_pc = io_executeStage_inst0_pc; // @[ExecuteUnit.scala 70:30]
  assign Fu_io_inst_0_hilo_wen = 4'hb == io_executeStage_inst0_inst_info_fusel | 4'hc ==
    io_executeStage_inst0_inst_info_fusel | 4'h9 == io_executeStage_inst0_inst_info_fusel; // @[ExecuteUnit.scala 71:76]
  assign Fu_io_inst_0_mul_en = io_executeStage_inst0_inst_info_fusel == 4'hb; // @[ExecuteUnit.scala 72:71]
  assign Fu_io_inst_0_div_en = io_executeStage_inst0_inst_info_fusel == 4'hc; // @[ExecuteUnit.scala 73:71]
  assign Fu_io_inst_0_inst_info_op = io_executeStage_inst0_inst_info_op; // @[ExecuteUnit.scala 74:30]
  assign Fu_io_inst_0_src_info_src1_data = io_executeStage_inst0_src_info_src1_data; // @[ExecuteUnit.scala 75:30]
  assign Fu_io_inst_0_src_info_src2_data = io_executeStage_inst0_src_info_src2_data; // @[ExecuteUnit.scala 75:30]
  assign Fu_io_inst_0_ex_in_flush_req = io_executeStage_inst0_ex_flush_req; // @[ExecuteUnit.scala 76:30]
  assign Fu_io_inst_0_ex_in_eret = io_executeStage_inst0_ex_eret; // @[ExecuteUnit.scala 76:30]
  assign Fu_io_inst_0_ex_in_badvaddr = io_executeStage_inst0_ex_badvaddr; // @[ExecuteUnit.scala 76:30]
  assign Fu_io_inst_0_ex_in_bd = io_executeStage_inst0_ex_bd; // @[ExecuteUnit.scala 76:30]
  assign Fu_io_inst_0_ex_in_excode = io_executeStage_inst0_ex_excode; // @[ExecuteUnit.scala 76:30]
  assign Fu_io_inst_1_hilo_wen = 4'hb == io_executeStage_inst1_inst_info_fusel | 4'hc ==
    io_executeStage_inst1_inst_info_fusel | 4'h9 == io_executeStage_inst1_inst_info_fusel; // @[ExecuteUnit.scala 78:76]
  assign Fu_io_inst_1_mul_en = io_executeStage_inst1_inst_info_fusel == 4'hb; // @[ExecuteUnit.scala 79:71]
  assign Fu_io_inst_1_div_en = io_executeStage_inst1_inst_info_fusel == 4'hc; // @[ExecuteUnit.scala 80:71]
  assign Fu_io_inst_1_inst_info_op = io_executeStage_inst1_inst_info_op; // @[ExecuteUnit.scala 81:30]
  assign Fu_io_inst_1_src_info_src1_data = io_executeStage_inst1_src_info_src1_data; // @[ExecuteUnit.scala 82:30]
  assign Fu_io_inst_1_src_info_src2_data = io_executeStage_inst1_src_info_src2_data; // @[ExecuteUnit.scala 82:30]
  assign Fu_io_inst_1_ex_in_flush_req = io_executeStage_inst1_ex_flush_req; // @[ExecuteUnit.scala 83:30]
  assign Fu_io_inst_1_ex_in_eret = io_executeStage_inst1_ex_eret; // @[ExecuteUnit.scala 83:30]
  assign Fu_io_inst_1_ex_in_badvaddr = io_executeStage_inst1_ex_badvaddr; // @[ExecuteUnit.scala 83:30]
  assign Fu_io_inst_1_ex_in_bd = io_executeStage_inst1_ex_bd; // @[ExecuteUnit.scala 83:30]
  assign Fu_io_inst_1_ex_in_excode = io_executeStage_inst1_ex_excode; // @[ExecuteUnit.scala 83:30]
  assign Fu_io_cp0_rdata = io_cp0_out_cp0_rdata; // @[ExecuteUnit.scala 84:30]
  assign Fu_io_branch_pred_branch_flag = io_executeStage_inst0_jb_info_pred_branch_flag; // @[ExecuteUnit.scala 85:30]
  assign ExeAccessMemCtrl_io_inst_0_inst_info_fusel = io_executeStage_inst0_inst_info_fusel; // @[ExecuteUnit.scala 60:35]
  assign ExeAccessMemCtrl_io_inst_0_inst_info_op = io_executeStage_inst0_inst_info_op; // @[ExecuteUnit.scala 60:35]
  assign ExeAccessMemCtrl_io_inst_0_inst_info_inst = io_executeStage_inst0_inst_info_inst; // @[ExecuteUnit.scala 60:35]
  assign ExeAccessMemCtrl_io_inst_0_src_info_src1_data = io_executeStage_inst0_src_info_src1_data; // @[ExecuteUnit.scala 61:35]
  assign ExeAccessMemCtrl_io_inst_0_src_info_src2_data = io_executeStage_inst0_src_info_src2_data; // @[ExecuteUnit.scala 61:35]
  assign ExeAccessMemCtrl_io_inst_0_ex_in_flush_req = io_executeStage_inst0_ex_flush_req; // @[ExecuteUnit.scala 62:35]
  assign ExeAccessMemCtrl_io_inst_0_ex_in_eret = io_executeStage_inst0_ex_eret; // @[ExecuteUnit.scala 62:35]
  assign ExeAccessMemCtrl_io_inst_0_ex_in_badvaddr = io_executeStage_inst0_ex_badvaddr; // @[ExecuteUnit.scala 62:35]
  assign ExeAccessMemCtrl_io_inst_0_ex_in_bd = io_executeStage_inst0_ex_bd; // @[ExecuteUnit.scala 62:35]
  assign ExeAccessMemCtrl_io_inst_0_ex_in_excode = io_executeStage_inst0_ex_excode; // @[ExecuteUnit.scala 62:35]
  assign ExeAccessMemCtrl_io_inst_1_inst_info_fusel = io_executeStage_inst1_inst_info_fusel; // @[ExecuteUnit.scala 63:35]
  assign ExeAccessMemCtrl_io_inst_1_inst_info_op = io_executeStage_inst1_inst_info_op; // @[ExecuteUnit.scala 63:35]
  assign ExeAccessMemCtrl_io_inst_1_inst_info_inst = io_executeStage_inst1_inst_info_inst; // @[ExecuteUnit.scala 63:35]
  assign ExeAccessMemCtrl_io_inst_1_src_info_src1_data = io_executeStage_inst1_src_info_src1_data; // @[ExecuteUnit.scala 64:35]
  assign ExeAccessMemCtrl_io_inst_1_src_info_src2_data = io_executeStage_inst1_src_info_src2_data; // @[ExecuteUnit.scala 64:35]
  assign ExeAccessMemCtrl_io_inst_1_ex_in_flush_req = io_executeStage_inst1_ex_flush_req; // @[ExecuteUnit.scala 65:35]
  assign ExeAccessMemCtrl_io_inst_1_ex_in_eret = io_executeStage_inst1_ex_eret; // @[ExecuteUnit.scala 65:35]
  assign ExeAccessMemCtrl_io_inst_1_ex_in_badvaddr = io_executeStage_inst1_ex_badvaddr; // @[ExecuteUnit.scala 65:35]
  assign ExeAccessMemCtrl_io_inst_1_ex_in_bd = io_executeStage_inst1_ex_bd; // @[ExecuteUnit.scala 65:35]
  assign ExeAccessMemCtrl_io_inst_1_ex_in_excode = io_executeStage_inst1_ex_excode; // @[ExecuteUnit.scala 65:35]
endmodule
module TlbL2(
  input         clock,
  input         reset,
  input         io_in_write_en,
  input  [2:0]  io_in_write_index,
  input  [18:0] io_in_write_entry_vpn2,
  input  [7:0]  io_in_write_entry_asid,
  input         io_in_write_entry_g,
  input  [19:0] io_in_write_entry_pfn_0,
  input  [19:0] io_in_write_entry_pfn_1,
  input         io_in_write_entry_c_0,
  input         io_in_write_entry_c_1,
  input         io_in_write_entry_d_0,
  input         io_in_write_entry_d_1,
  input         io_in_write_entry_v_0,
  input         io_in_write_entry_v_1,
  input  [2:0]  io_in_read_index,
  input  [18:0] io_in_entry_hi_vpn2,
  input  [7:0]  io_in_entry_hi_asid,
  input  [18:0] io_in_tlb1_vpn2,
  input  [18:0] io_in_tlb2_vpn2,
  output        io_out_read_entry_g,
  output [19:0] io_out_read_entry_pfn_0,
  output [19:0] io_out_read_entry_pfn_1,
  output        io_out_read_entry_c_0,
  output        io_out_read_entry_c_1,
  output        io_out_read_entry_d_0,
  output        io_out_read_entry_d_1,
  output        io_out_read_entry_v_0,
  output        io_out_read_entry_v_1,
  output        io_out_tlb1_found,
  output        io_out_tlb2_found,
  output [19:0] io_out_tlb1_entry_pfn_0,
  output [19:0] io_out_tlb1_entry_pfn_1,
  output        io_out_tlb1_entry_c_0,
  output        io_out_tlb1_entry_c_1,
  output        io_out_tlb1_entry_v_0,
  output        io_out_tlb1_entry_v_1,
  output [19:0] io_out_tlb2_entry_pfn_0,
  output [19:0] io_out_tlb2_entry_pfn_1,
  output        io_out_tlb2_entry_c_0,
  output        io_out_tlb2_entry_c_1,
  output        io_out_tlb2_entry_d_0,
  output        io_out_tlb2_entry_d_1,
  output        io_out_tlb2_entry_v_0,
  output        io_out_tlb2_entry_v_1,
  output        io_out_tlb_found,
  output [2:0]  io_out_tlb_match_index
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
`endif // RANDOMIZE_REG_INIT
  reg [18:0] tlb_l2_0_vpn2; // @[TlbL2.scala 39:23]
  reg [7:0] tlb_l2_0_asid; // @[TlbL2.scala 39:23]
  reg  tlb_l2_0_g; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_0_pfn_0; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_0_pfn_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_0_c_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_0_c_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_0_d_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_0_d_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_0_v_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_0_v_1; // @[TlbL2.scala 39:23]
  reg [18:0] tlb_l2_1_vpn2; // @[TlbL2.scala 39:23]
  reg [7:0] tlb_l2_1_asid; // @[TlbL2.scala 39:23]
  reg  tlb_l2_1_g; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_1_pfn_0; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_1_pfn_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_1_c_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_1_c_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_1_d_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_1_d_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_1_v_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_1_v_1; // @[TlbL2.scala 39:23]
  reg [18:0] tlb_l2_2_vpn2; // @[TlbL2.scala 39:23]
  reg [7:0] tlb_l2_2_asid; // @[TlbL2.scala 39:23]
  reg  tlb_l2_2_g; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_2_pfn_0; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_2_pfn_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_2_c_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_2_c_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_2_d_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_2_d_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_2_v_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_2_v_1; // @[TlbL2.scala 39:23]
  reg [18:0] tlb_l2_3_vpn2; // @[TlbL2.scala 39:23]
  reg [7:0] tlb_l2_3_asid; // @[TlbL2.scala 39:23]
  reg  tlb_l2_3_g; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_3_pfn_0; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_3_pfn_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_3_c_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_3_c_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_3_d_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_3_d_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_3_v_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_3_v_1; // @[TlbL2.scala 39:23]
  reg [18:0] tlb_l2_4_vpn2; // @[TlbL2.scala 39:23]
  reg [7:0] tlb_l2_4_asid; // @[TlbL2.scala 39:23]
  reg  tlb_l2_4_g; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_4_pfn_0; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_4_pfn_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_4_c_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_4_c_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_4_d_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_4_d_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_4_v_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_4_v_1; // @[TlbL2.scala 39:23]
  reg [18:0] tlb_l2_5_vpn2; // @[TlbL2.scala 39:23]
  reg [7:0] tlb_l2_5_asid; // @[TlbL2.scala 39:23]
  reg  tlb_l2_5_g; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_5_pfn_0; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_5_pfn_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_5_c_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_5_c_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_5_d_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_5_d_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_5_v_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_5_v_1; // @[TlbL2.scala 39:23]
  reg [18:0] tlb_l2_6_vpn2; // @[TlbL2.scala 39:23]
  reg [7:0] tlb_l2_6_asid; // @[TlbL2.scala 39:23]
  reg  tlb_l2_6_g; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_6_pfn_0; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_6_pfn_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_6_c_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_6_c_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_6_d_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_6_d_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_6_v_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_6_v_1; // @[TlbL2.scala 39:23]
  reg [18:0] tlb_l2_7_vpn2; // @[TlbL2.scala 39:23]
  reg [7:0] tlb_l2_7_asid; // @[TlbL2.scala 39:23]
  reg  tlb_l2_7_g; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_7_pfn_0; // @[TlbL2.scala 39:23]
  reg [19:0] tlb_l2_7_pfn_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_7_c_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_7_c_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_7_d_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_7_d_1; // @[TlbL2.scala 39:23]
  reg  tlb_l2_7_v_0; // @[TlbL2.scala 39:23]
  reg  tlb_l2_7_v_1; // @[TlbL2.scala 39:23]
  wire  _tlb_match_1_1_T_2 = tlb_l2_1_vpn2 == io_in_tlb1_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_1_1 = (tlb_l2_1_g | tlb_l2_1_asid == io_in_entry_hi_asid) & _tlb_match_1_1_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_1_0_T_2 = tlb_l2_0_vpn2 == io_in_tlb1_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_1_0 = (tlb_l2_0_g | tlb_l2_0_asid == io_in_entry_hi_asid) & _tlb_match_1_0_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_1_3_T_2 = tlb_l2_3_vpn2 == io_in_tlb1_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_1_3 = (tlb_l2_3_g | tlb_l2_3_asid == io_in_entry_hi_asid) & _tlb_match_1_3_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_1_2_T_2 = tlb_l2_2_vpn2 == io_in_tlb1_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_1_2 = (tlb_l2_2_g | tlb_l2_2_asid == io_in_entry_hi_asid) & _tlb_match_1_2_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_1_5_T_2 = tlb_l2_5_vpn2 == io_in_tlb1_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_1_5 = (tlb_l2_5_g | tlb_l2_5_asid == io_in_entry_hi_asid) & _tlb_match_1_5_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_1_4_T_2 = tlb_l2_4_vpn2 == io_in_tlb1_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_1_4 = (tlb_l2_4_g | tlb_l2_4_asid == io_in_entry_hi_asid) & _tlb_match_1_4_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_1_7_T_2 = tlb_l2_7_vpn2 == io_in_tlb1_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_1_7 = (tlb_l2_7_g | tlb_l2_7_asid == io_in_entry_hi_asid) & _tlb_match_1_7_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_1_6_T_2 = tlb_l2_6_vpn2 == io_in_tlb1_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_1_6 = (tlb_l2_6_g | tlb_l2_6_asid == io_in_entry_hi_asid) & _tlb_match_1_6_T_2; // @[TlbL2.scala 59:82]
  wire [7:0] _io_out_tlb1_found_T = {tlb_match_1_7,tlb_match_1_6,tlb_match_1_5,tlb_match_1_4,tlb_match_1_3,tlb_match_1_2
    ,tlb_match_1_1,tlb_match_1_0}; // @[TlbL2.scala 49:42]
  wire  _tlb_match_2_1_T_2 = tlb_l2_1_vpn2 == io_in_tlb2_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_2_1 = (tlb_l2_1_g | tlb_l2_1_asid == io_in_entry_hi_asid) & _tlb_match_2_1_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_2_0_T_2 = tlb_l2_0_vpn2 == io_in_tlb2_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_2_0 = (tlb_l2_0_g | tlb_l2_0_asid == io_in_entry_hi_asid) & _tlb_match_2_0_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_2_3_T_2 = tlb_l2_3_vpn2 == io_in_tlb2_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_2_3 = (tlb_l2_3_g | tlb_l2_3_asid == io_in_entry_hi_asid) & _tlb_match_2_3_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_2_2_T_2 = tlb_l2_2_vpn2 == io_in_tlb2_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_2_2 = (tlb_l2_2_g | tlb_l2_2_asid == io_in_entry_hi_asid) & _tlb_match_2_2_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_2_5_T_2 = tlb_l2_5_vpn2 == io_in_tlb2_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_2_5 = (tlb_l2_5_g | tlb_l2_5_asid == io_in_entry_hi_asid) & _tlb_match_2_5_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_2_4_T_2 = tlb_l2_4_vpn2 == io_in_tlb2_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_2_4 = (tlb_l2_4_g | tlb_l2_4_asid == io_in_entry_hi_asid) & _tlb_match_2_4_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_2_7_T_2 = tlb_l2_7_vpn2 == io_in_tlb2_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_2_7 = (tlb_l2_7_g | tlb_l2_7_asid == io_in_entry_hi_asid) & _tlb_match_2_7_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_2_6_T_2 = tlb_l2_6_vpn2 == io_in_tlb2_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_2_6 = (tlb_l2_6_g | tlb_l2_6_asid == io_in_entry_hi_asid) & _tlb_match_2_6_T_2; // @[TlbL2.scala 59:82]
  wire [7:0] _io_out_tlb2_found_T = {tlb_match_2_7,tlb_match_2_6,tlb_match_2_5,tlb_match_2_4,tlb_match_2_3,tlb_match_2_2
    ,tlb_match_2_1,tlb_match_2_0}; // @[TlbL2.scala 50:42]
  wire [2:0] _tlb_match_index_1_T = tlb_match_1_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_1_T_1 = tlb_match_1_5 ? 3'h5 : _tlb_match_index_1_T; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_1_T_2 = tlb_match_1_4 ? 3'h4 : _tlb_match_index_1_T_1; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_1_T_3 = tlb_match_1_3 ? 3'h3 : _tlb_match_index_1_T_2; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_1_T_4 = tlb_match_1_2 ? 3'h2 : _tlb_match_index_1_T_3; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_1_T_5 = tlb_match_1_1 ? 3'h1 : _tlb_match_index_1_T_4; // @[Mux.scala 47:70]
  wire [2:0] tlb_match_index_1 = tlb_match_1_0 ? 3'h0 : _tlb_match_index_1_T_5; // @[Mux.scala 47:70]
  wire [19:0] _GEN_25 = 3'h1 == tlb_match_index_1 ? tlb_l2_1_pfn_0 : tlb_l2_0_pfn_0; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_26 = 3'h2 == tlb_match_index_1 ? tlb_l2_2_pfn_0 : _GEN_25; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_27 = 3'h3 == tlb_match_index_1 ? tlb_l2_3_pfn_0 : _GEN_26; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_28 = 3'h4 == tlb_match_index_1 ? tlb_l2_4_pfn_0 : _GEN_27; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_29 = 3'h5 == tlb_match_index_1 ? tlb_l2_5_pfn_0 : _GEN_28; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_30 = 3'h6 == tlb_match_index_1 ? tlb_l2_6_pfn_0 : _GEN_29; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_33 = 3'h1 == tlb_match_index_1 ? tlb_l2_1_pfn_1 : tlb_l2_0_pfn_1; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_34 = 3'h2 == tlb_match_index_1 ? tlb_l2_2_pfn_1 : _GEN_33; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_35 = 3'h3 == tlb_match_index_1 ? tlb_l2_3_pfn_1 : _GEN_34; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_36 = 3'h4 == tlb_match_index_1 ? tlb_l2_4_pfn_1 : _GEN_35; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_37 = 3'h5 == tlb_match_index_1 ? tlb_l2_5_pfn_1 : _GEN_36; // @[TlbL2.scala 51:{26,26}]
  wire [19:0] _GEN_38 = 3'h6 == tlb_match_index_1 ? tlb_l2_6_pfn_1 : _GEN_37; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_41 = 3'h1 == tlb_match_index_1 ? tlb_l2_1_c_0 : tlb_l2_0_c_0; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_42 = 3'h2 == tlb_match_index_1 ? tlb_l2_2_c_0 : _GEN_41; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_43 = 3'h3 == tlb_match_index_1 ? tlb_l2_3_c_0 : _GEN_42; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_44 = 3'h4 == tlb_match_index_1 ? tlb_l2_4_c_0 : _GEN_43; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_45 = 3'h5 == tlb_match_index_1 ? tlb_l2_5_c_0 : _GEN_44; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_46 = 3'h6 == tlb_match_index_1 ? tlb_l2_6_c_0 : _GEN_45; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_49 = 3'h1 == tlb_match_index_1 ? tlb_l2_1_c_1 : tlb_l2_0_c_1; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_50 = 3'h2 == tlb_match_index_1 ? tlb_l2_2_c_1 : _GEN_49; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_51 = 3'h3 == tlb_match_index_1 ? tlb_l2_3_c_1 : _GEN_50; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_52 = 3'h4 == tlb_match_index_1 ? tlb_l2_4_c_1 : _GEN_51; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_53 = 3'h5 == tlb_match_index_1 ? tlb_l2_5_c_1 : _GEN_52; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_54 = 3'h6 == tlb_match_index_1 ? tlb_l2_6_c_1 : _GEN_53; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_73 = 3'h1 == tlb_match_index_1 ? tlb_l2_1_v_0 : tlb_l2_0_v_0; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_74 = 3'h2 == tlb_match_index_1 ? tlb_l2_2_v_0 : _GEN_73; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_75 = 3'h3 == tlb_match_index_1 ? tlb_l2_3_v_0 : _GEN_74; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_76 = 3'h4 == tlb_match_index_1 ? tlb_l2_4_v_0 : _GEN_75; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_77 = 3'h5 == tlb_match_index_1 ? tlb_l2_5_v_0 : _GEN_76; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_78 = 3'h6 == tlb_match_index_1 ? tlb_l2_6_v_0 : _GEN_77; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_81 = 3'h1 == tlb_match_index_1 ? tlb_l2_1_v_1 : tlb_l2_0_v_1; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_82 = 3'h2 == tlb_match_index_1 ? tlb_l2_2_v_1 : _GEN_81; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_83 = 3'h3 == tlb_match_index_1 ? tlb_l2_3_v_1 : _GEN_82; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_84 = 3'h4 == tlb_match_index_1 ? tlb_l2_4_v_1 : _GEN_83; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_85 = 3'h5 == tlb_match_index_1 ? tlb_l2_5_v_1 : _GEN_84; // @[TlbL2.scala 51:{26,26}]
  wire  _GEN_86 = 3'h6 == tlb_match_index_1 ? tlb_l2_6_v_1 : _GEN_85; // @[TlbL2.scala 51:{26,26}]
  wire [2:0] _tlb_match_index_2_T = tlb_match_2_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_2_T_1 = tlb_match_2_5 ? 3'h5 : _tlb_match_index_2_T; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_2_T_2 = tlb_match_2_4 ? 3'h4 : _tlb_match_index_2_T_1; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_2_T_3 = tlb_match_2_3 ? 3'h3 : _tlb_match_index_2_T_2; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_2_T_4 = tlb_match_2_2 ? 3'h2 : _tlb_match_index_2_T_3; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_2_T_5 = tlb_match_2_1 ? 3'h1 : _tlb_match_index_2_T_4; // @[Mux.scala 47:70]
  wire [2:0] tlb_match_index_2 = tlb_match_2_0 ? 3'h0 : _tlb_match_index_2_T_5; // @[Mux.scala 47:70]
  wire [19:0] _GEN_113 = 3'h1 == tlb_match_index_2 ? tlb_l2_1_pfn_0 : tlb_l2_0_pfn_0; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_114 = 3'h2 == tlb_match_index_2 ? tlb_l2_2_pfn_0 : _GEN_113; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_115 = 3'h3 == tlb_match_index_2 ? tlb_l2_3_pfn_0 : _GEN_114; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_116 = 3'h4 == tlb_match_index_2 ? tlb_l2_4_pfn_0 : _GEN_115; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_117 = 3'h5 == tlb_match_index_2 ? tlb_l2_5_pfn_0 : _GEN_116; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_118 = 3'h6 == tlb_match_index_2 ? tlb_l2_6_pfn_0 : _GEN_117; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_121 = 3'h1 == tlb_match_index_2 ? tlb_l2_1_pfn_1 : tlb_l2_0_pfn_1; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_122 = 3'h2 == tlb_match_index_2 ? tlb_l2_2_pfn_1 : _GEN_121; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_123 = 3'h3 == tlb_match_index_2 ? tlb_l2_3_pfn_1 : _GEN_122; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_124 = 3'h4 == tlb_match_index_2 ? tlb_l2_4_pfn_1 : _GEN_123; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_125 = 3'h5 == tlb_match_index_2 ? tlb_l2_5_pfn_1 : _GEN_124; // @[TlbL2.scala 52:{26,26}]
  wire [19:0] _GEN_126 = 3'h6 == tlb_match_index_2 ? tlb_l2_6_pfn_1 : _GEN_125; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_129 = 3'h1 == tlb_match_index_2 ? tlb_l2_1_c_0 : tlb_l2_0_c_0; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_130 = 3'h2 == tlb_match_index_2 ? tlb_l2_2_c_0 : _GEN_129; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_131 = 3'h3 == tlb_match_index_2 ? tlb_l2_3_c_0 : _GEN_130; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_132 = 3'h4 == tlb_match_index_2 ? tlb_l2_4_c_0 : _GEN_131; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_133 = 3'h5 == tlb_match_index_2 ? tlb_l2_5_c_0 : _GEN_132; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_134 = 3'h6 == tlb_match_index_2 ? tlb_l2_6_c_0 : _GEN_133; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_137 = 3'h1 == tlb_match_index_2 ? tlb_l2_1_c_1 : tlb_l2_0_c_1; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_138 = 3'h2 == tlb_match_index_2 ? tlb_l2_2_c_1 : _GEN_137; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_139 = 3'h3 == tlb_match_index_2 ? tlb_l2_3_c_1 : _GEN_138; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_140 = 3'h4 == tlb_match_index_2 ? tlb_l2_4_c_1 : _GEN_139; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_141 = 3'h5 == tlb_match_index_2 ? tlb_l2_5_c_1 : _GEN_140; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_142 = 3'h6 == tlb_match_index_2 ? tlb_l2_6_c_1 : _GEN_141; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_145 = 3'h1 == tlb_match_index_2 ? tlb_l2_1_d_0 : tlb_l2_0_d_0; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_146 = 3'h2 == tlb_match_index_2 ? tlb_l2_2_d_0 : _GEN_145; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_147 = 3'h3 == tlb_match_index_2 ? tlb_l2_3_d_0 : _GEN_146; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_148 = 3'h4 == tlb_match_index_2 ? tlb_l2_4_d_0 : _GEN_147; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_149 = 3'h5 == tlb_match_index_2 ? tlb_l2_5_d_0 : _GEN_148; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_150 = 3'h6 == tlb_match_index_2 ? tlb_l2_6_d_0 : _GEN_149; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_153 = 3'h1 == tlb_match_index_2 ? tlb_l2_1_d_1 : tlb_l2_0_d_1; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_154 = 3'h2 == tlb_match_index_2 ? tlb_l2_2_d_1 : _GEN_153; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_155 = 3'h3 == tlb_match_index_2 ? tlb_l2_3_d_1 : _GEN_154; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_156 = 3'h4 == tlb_match_index_2 ? tlb_l2_4_d_1 : _GEN_155; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_157 = 3'h5 == tlb_match_index_2 ? tlb_l2_5_d_1 : _GEN_156; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_158 = 3'h6 == tlb_match_index_2 ? tlb_l2_6_d_1 : _GEN_157; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_161 = 3'h1 == tlb_match_index_2 ? tlb_l2_1_v_0 : tlb_l2_0_v_0; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_162 = 3'h2 == tlb_match_index_2 ? tlb_l2_2_v_0 : _GEN_161; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_163 = 3'h3 == tlb_match_index_2 ? tlb_l2_3_v_0 : _GEN_162; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_164 = 3'h4 == tlb_match_index_2 ? tlb_l2_4_v_0 : _GEN_163; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_165 = 3'h5 == tlb_match_index_2 ? tlb_l2_5_v_0 : _GEN_164; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_166 = 3'h6 == tlb_match_index_2 ? tlb_l2_6_v_0 : _GEN_165; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_169 = 3'h1 == tlb_match_index_2 ? tlb_l2_1_v_1 : tlb_l2_0_v_1; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_170 = 3'h2 == tlb_match_index_2 ? tlb_l2_2_v_1 : _GEN_169; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_171 = 3'h3 == tlb_match_index_2 ? tlb_l2_3_v_1 : _GEN_170; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_172 = 3'h4 == tlb_match_index_2 ? tlb_l2_4_v_1 : _GEN_171; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_173 = 3'h5 == tlb_match_index_2 ? tlb_l2_5_v_1 : _GEN_172; // @[TlbL2.scala 52:{26,26}]
  wire  _GEN_174 = 3'h6 == tlb_match_index_2 ? tlb_l2_6_v_1 : _GEN_173; // @[TlbL2.scala 52:{26,26}]
  wire  _tlb_match_0_1_T_2 = tlb_l2_1_vpn2 == io_in_entry_hi_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_0_1 = (tlb_l2_1_g | tlb_l2_1_asid == io_in_entry_hi_asid) & _tlb_match_0_1_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_0_0_T_2 = tlb_l2_0_vpn2 == io_in_entry_hi_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_0_0 = (tlb_l2_0_g | tlb_l2_0_asid == io_in_entry_hi_asid) & _tlb_match_0_0_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_0_3_T_2 = tlb_l2_3_vpn2 == io_in_entry_hi_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_0_3 = (tlb_l2_3_g | tlb_l2_3_asid == io_in_entry_hi_asid) & _tlb_match_0_3_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_0_2_T_2 = tlb_l2_2_vpn2 == io_in_entry_hi_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_0_2 = (tlb_l2_2_g | tlb_l2_2_asid == io_in_entry_hi_asid) & _tlb_match_0_2_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_0_5_T_2 = tlb_l2_5_vpn2 == io_in_entry_hi_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_0_5 = (tlb_l2_5_g | tlb_l2_5_asid == io_in_entry_hi_asid) & _tlb_match_0_5_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_0_4_T_2 = tlb_l2_4_vpn2 == io_in_entry_hi_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_0_4 = (tlb_l2_4_g | tlb_l2_4_asid == io_in_entry_hi_asid) & _tlb_match_0_4_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_0_7_T_2 = tlb_l2_7_vpn2 == io_in_entry_hi_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_0_7 = (tlb_l2_7_g | tlb_l2_7_asid == io_in_entry_hi_asid) & _tlb_match_0_7_T_2; // @[TlbL2.scala 59:82]
  wire  _tlb_match_0_6_T_2 = tlb_l2_6_vpn2 == io_in_entry_hi_vpn2; // @[TlbL2.scala 60:25]
  wire  tlb_match_0_6 = (tlb_l2_6_g | tlb_l2_6_asid == io_in_entry_hi_asid) & _tlb_match_0_6_T_2; // @[TlbL2.scala 59:82]
  wire [7:0] _io_out_tlb_found_T = {tlb_match_0_7,tlb_match_0_6,tlb_match_0_5,tlb_match_0_4,tlb_match_0_3,tlb_match_0_2,
    tlb_match_0_1,tlb_match_0_0}; // @[TlbL2.scala 53:42]
  wire  _GEN_193 = 3'h1 == io_in_read_index ? tlb_l2_1_g : tlb_l2_0_g; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_194 = 3'h2 == io_in_read_index ? tlb_l2_2_g : _GEN_193; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_195 = 3'h3 == io_in_read_index ? tlb_l2_3_g : _GEN_194; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_196 = 3'h4 == io_in_read_index ? tlb_l2_4_g : _GEN_195; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_197 = 3'h5 == io_in_read_index ? tlb_l2_5_g : _GEN_196; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_198 = 3'h6 == io_in_read_index ? tlb_l2_6_g : _GEN_197; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_201 = 3'h1 == io_in_read_index ? tlb_l2_1_pfn_0 : tlb_l2_0_pfn_0; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_202 = 3'h2 == io_in_read_index ? tlb_l2_2_pfn_0 : _GEN_201; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_203 = 3'h3 == io_in_read_index ? tlb_l2_3_pfn_0 : _GEN_202; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_204 = 3'h4 == io_in_read_index ? tlb_l2_4_pfn_0 : _GEN_203; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_205 = 3'h5 == io_in_read_index ? tlb_l2_5_pfn_0 : _GEN_204; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_206 = 3'h6 == io_in_read_index ? tlb_l2_6_pfn_0 : _GEN_205; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_209 = 3'h1 == io_in_read_index ? tlb_l2_1_pfn_1 : tlb_l2_0_pfn_1; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_210 = 3'h2 == io_in_read_index ? tlb_l2_2_pfn_1 : _GEN_209; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_211 = 3'h3 == io_in_read_index ? tlb_l2_3_pfn_1 : _GEN_210; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_212 = 3'h4 == io_in_read_index ? tlb_l2_4_pfn_1 : _GEN_211; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_213 = 3'h5 == io_in_read_index ? tlb_l2_5_pfn_1 : _GEN_212; // @[TlbL2.scala 55:{26,26}]
  wire [19:0] _GEN_214 = 3'h6 == io_in_read_index ? tlb_l2_6_pfn_1 : _GEN_213; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_217 = 3'h1 == io_in_read_index ? tlb_l2_1_c_0 : tlb_l2_0_c_0; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_218 = 3'h2 == io_in_read_index ? tlb_l2_2_c_0 : _GEN_217; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_219 = 3'h3 == io_in_read_index ? tlb_l2_3_c_0 : _GEN_218; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_220 = 3'h4 == io_in_read_index ? tlb_l2_4_c_0 : _GEN_219; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_221 = 3'h5 == io_in_read_index ? tlb_l2_5_c_0 : _GEN_220; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_222 = 3'h6 == io_in_read_index ? tlb_l2_6_c_0 : _GEN_221; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_225 = 3'h1 == io_in_read_index ? tlb_l2_1_c_1 : tlb_l2_0_c_1; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_226 = 3'h2 == io_in_read_index ? tlb_l2_2_c_1 : _GEN_225; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_227 = 3'h3 == io_in_read_index ? tlb_l2_3_c_1 : _GEN_226; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_228 = 3'h4 == io_in_read_index ? tlb_l2_4_c_1 : _GEN_227; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_229 = 3'h5 == io_in_read_index ? tlb_l2_5_c_1 : _GEN_228; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_230 = 3'h6 == io_in_read_index ? tlb_l2_6_c_1 : _GEN_229; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_233 = 3'h1 == io_in_read_index ? tlb_l2_1_d_0 : tlb_l2_0_d_0; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_234 = 3'h2 == io_in_read_index ? tlb_l2_2_d_0 : _GEN_233; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_235 = 3'h3 == io_in_read_index ? tlb_l2_3_d_0 : _GEN_234; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_236 = 3'h4 == io_in_read_index ? tlb_l2_4_d_0 : _GEN_235; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_237 = 3'h5 == io_in_read_index ? tlb_l2_5_d_0 : _GEN_236; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_238 = 3'h6 == io_in_read_index ? tlb_l2_6_d_0 : _GEN_237; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_241 = 3'h1 == io_in_read_index ? tlb_l2_1_d_1 : tlb_l2_0_d_1; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_242 = 3'h2 == io_in_read_index ? tlb_l2_2_d_1 : _GEN_241; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_243 = 3'h3 == io_in_read_index ? tlb_l2_3_d_1 : _GEN_242; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_244 = 3'h4 == io_in_read_index ? tlb_l2_4_d_1 : _GEN_243; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_245 = 3'h5 == io_in_read_index ? tlb_l2_5_d_1 : _GEN_244; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_246 = 3'h6 == io_in_read_index ? tlb_l2_6_d_1 : _GEN_245; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_249 = 3'h1 == io_in_read_index ? tlb_l2_1_v_0 : tlb_l2_0_v_0; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_250 = 3'h2 == io_in_read_index ? tlb_l2_2_v_0 : _GEN_249; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_251 = 3'h3 == io_in_read_index ? tlb_l2_3_v_0 : _GEN_250; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_252 = 3'h4 == io_in_read_index ? tlb_l2_4_v_0 : _GEN_251; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_253 = 3'h5 == io_in_read_index ? tlb_l2_5_v_0 : _GEN_252; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_254 = 3'h6 == io_in_read_index ? tlb_l2_6_v_0 : _GEN_253; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_257 = 3'h1 == io_in_read_index ? tlb_l2_1_v_1 : tlb_l2_0_v_1; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_258 = 3'h2 == io_in_read_index ? tlb_l2_2_v_1 : _GEN_257; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_259 = 3'h3 == io_in_read_index ? tlb_l2_3_v_1 : _GEN_258; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_260 = 3'h4 == io_in_read_index ? tlb_l2_4_v_1 : _GEN_259; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_261 = 3'h5 == io_in_read_index ? tlb_l2_5_v_1 : _GEN_260; // @[TlbL2.scala 55:{26,26}]
  wire  _GEN_262 = 3'h6 == io_in_read_index ? tlb_l2_6_v_1 : _GEN_261; // @[TlbL2.scala 55:{26,26}]
  wire [2:0] _tlb_match_index_0_T = tlb_match_0_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_0_T_1 = tlb_match_0_5 ? 3'h5 : _tlb_match_index_0_T; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_0_T_2 = tlb_match_0_4 ? 3'h4 : _tlb_match_index_0_T_1; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_0_T_3 = tlb_match_0_3 ? 3'h3 : _tlb_match_index_0_T_2; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_0_T_4 = tlb_match_0_2 ? 3'h2 : _tlb_match_index_0_T_3; // @[Mux.scala 47:70]
  wire [2:0] _tlb_match_index_0_T_5 = tlb_match_0_1 ? 3'h1 : _tlb_match_index_0_T_4; // @[Mux.scala 47:70]
  assign io_out_read_entry_g = 3'h7 == io_in_read_index ? tlb_l2_7_g : _GEN_198; // @[TlbL2.scala 55:{26,26}]
  assign io_out_read_entry_pfn_0 = 3'h7 == io_in_read_index ? tlb_l2_7_pfn_0 : _GEN_206; // @[TlbL2.scala 55:{26,26}]
  assign io_out_read_entry_pfn_1 = 3'h7 == io_in_read_index ? tlb_l2_7_pfn_1 : _GEN_214; // @[TlbL2.scala 55:{26,26}]
  assign io_out_read_entry_c_0 = 3'h7 == io_in_read_index ? tlb_l2_7_c_0 : _GEN_222; // @[TlbL2.scala 55:{26,26}]
  assign io_out_read_entry_c_1 = 3'h7 == io_in_read_index ? tlb_l2_7_c_1 : _GEN_230; // @[TlbL2.scala 55:{26,26}]
  assign io_out_read_entry_d_0 = 3'h7 == io_in_read_index ? tlb_l2_7_d_0 : _GEN_238; // @[TlbL2.scala 55:{26,26}]
  assign io_out_read_entry_d_1 = 3'h7 == io_in_read_index ? tlb_l2_7_d_1 : _GEN_246; // @[TlbL2.scala 55:{26,26}]
  assign io_out_read_entry_v_0 = 3'h7 == io_in_read_index ? tlb_l2_7_v_0 : _GEN_254; // @[TlbL2.scala 55:{26,26}]
  assign io_out_read_entry_v_1 = 3'h7 == io_in_read_index ? tlb_l2_7_v_1 : _GEN_262; // @[TlbL2.scala 55:{26,26}]
  assign io_out_tlb1_found = |_io_out_tlb1_found_T; // @[TlbL2.scala 49:49]
  assign io_out_tlb2_found = |_io_out_tlb2_found_T; // @[TlbL2.scala 50:49]
  assign io_out_tlb1_entry_pfn_0 = 3'h7 == tlb_match_index_1 ? tlb_l2_7_pfn_0 : _GEN_30; // @[TlbL2.scala 51:{26,26}]
  assign io_out_tlb1_entry_pfn_1 = 3'h7 == tlb_match_index_1 ? tlb_l2_7_pfn_1 : _GEN_38; // @[TlbL2.scala 51:{26,26}]
  assign io_out_tlb1_entry_c_0 = 3'h7 == tlb_match_index_1 ? tlb_l2_7_c_0 : _GEN_46; // @[TlbL2.scala 51:{26,26}]
  assign io_out_tlb1_entry_c_1 = 3'h7 == tlb_match_index_1 ? tlb_l2_7_c_1 : _GEN_54; // @[TlbL2.scala 51:{26,26}]
  assign io_out_tlb1_entry_v_0 = 3'h7 == tlb_match_index_1 ? tlb_l2_7_v_0 : _GEN_78; // @[TlbL2.scala 51:{26,26}]
  assign io_out_tlb1_entry_v_1 = 3'h7 == tlb_match_index_1 ? tlb_l2_7_v_1 : _GEN_86; // @[TlbL2.scala 51:{26,26}]
  assign io_out_tlb2_entry_pfn_0 = 3'h7 == tlb_match_index_2 ? tlb_l2_7_pfn_0 : _GEN_118; // @[TlbL2.scala 52:{26,26}]
  assign io_out_tlb2_entry_pfn_1 = 3'h7 == tlb_match_index_2 ? tlb_l2_7_pfn_1 : _GEN_126; // @[TlbL2.scala 52:{26,26}]
  assign io_out_tlb2_entry_c_0 = 3'h7 == tlb_match_index_2 ? tlb_l2_7_c_0 : _GEN_134; // @[TlbL2.scala 52:{26,26}]
  assign io_out_tlb2_entry_c_1 = 3'h7 == tlb_match_index_2 ? tlb_l2_7_c_1 : _GEN_142; // @[TlbL2.scala 52:{26,26}]
  assign io_out_tlb2_entry_d_0 = 3'h7 == tlb_match_index_2 ? tlb_l2_7_d_0 : _GEN_150; // @[TlbL2.scala 52:{26,26}]
  assign io_out_tlb2_entry_d_1 = 3'h7 == tlb_match_index_2 ? tlb_l2_7_d_1 : _GEN_158; // @[TlbL2.scala 52:{26,26}]
  assign io_out_tlb2_entry_v_0 = 3'h7 == tlb_match_index_2 ? tlb_l2_7_v_0 : _GEN_166; // @[TlbL2.scala 52:{26,26}]
  assign io_out_tlb2_entry_v_1 = 3'h7 == tlb_match_index_2 ? tlb_l2_7_v_1 : _GEN_174; // @[TlbL2.scala 52:{26,26}]
  assign io_out_tlb_found = |_io_out_tlb_found_T; // @[TlbL2.scala 53:49]
  assign io_out_tlb_match_index = tlb_match_0_0 ? 3'h0 : _tlb_match_index_0_T_5; // @[Mux.scala 47:70]
  always @(posedge clock) begin
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_vpn2 <= 19'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_vpn2 <= io_in_write_entry_vpn2; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_asid <= 8'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_asid <= io_in_write_entry_asid; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_g <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_g <= io_in_write_entry_g; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_pfn_0 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_pfn_0 <= io_in_write_entry_pfn_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_pfn_1 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_pfn_1 <= io_in_write_entry_pfn_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_c_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_c_0 <= io_in_write_entry_c_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_c_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_c_1 <= io_in_write_entry_c_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_d_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_d_0 <= io_in_write_entry_d_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_d_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_d_1 <= io_in_write_entry_d_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_v_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_v_0 <= io_in_write_entry_v_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_0_v_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h0 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_0_v_1 <= io_in_write_entry_v_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_vpn2 <= 19'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_vpn2 <= io_in_write_entry_vpn2; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_asid <= 8'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_asid <= io_in_write_entry_asid; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_g <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_g <= io_in_write_entry_g; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_pfn_0 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_pfn_0 <= io_in_write_entry_pfn_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_pfn_1 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_pfn_1 <= io_in_write_entry_pfn_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_c_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_c_0 <= io_in_write_entry_c_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_c_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_c_1 <= io_in_write_entry_c_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_d_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_d_0 <= io_in_write_entry_d_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_d_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_d_1 <= io_in_write_entry_d_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_v_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_v_0 <= io_in_write_entry_v_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_1_v_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h1 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_1_v_1 <= io_in_write_entry_v_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_vpn2 <= 19'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_vpn2 <= io_in_write_entry_vpn2; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_asid <= 8'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_asid <= io_in_write_entry_asid; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_g <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_g <= io_in_write_entry_g; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_pfn_0 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_pfn_0 <= io_in_write_entry_pfn_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_pfn_1 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_pfn_1 <= io_in_write_entry_pfn_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_c_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_c_0 <= io_in_write_entry_c_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_c_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_c_1 <= io_in_write_entry_c_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_d_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_d_0 <= io_in_write_entry_d_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_d_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_d_1 <= io_in_write_entry_d_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_v_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_v_0 <= io_in_write_entry_v_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_2_v_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h2 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_2_v_1 <= io_in_write_entry_v_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_vpn2 <= 19'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_vpn2 <= io_in_write_entry_vpn2; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_asid <= 8'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_asid <= io_in_write_entry_asid; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_g <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_g <= io_in_write_entry_g; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_pfn_0 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_pfn_0 <= io_in_write_entry_pfn_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_pfn_1 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_pfn_1 <= io_in_write_entry_pfn_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_c_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_c_0 <= io_in_write_entry_c_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_c_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_c_1 <= io_in_write_entry_c_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_d_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_d_0 <= io_in_write_entry_d_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_d_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_d_1 <= io_in_write_entry_d_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_v_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_v_0 <= io_in_write_entry_v_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_3_v_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h3 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_3_v_1 <= io_in_write_entry_v_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_vpn2 <= 19'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_vpn2 <= io_in_write_entry_vpn2; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_asid <= 8'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_asid <= io_in_write_entry_asid; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_g <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_g <= io_in_write_entry_g; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_pfn_0 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_pfn_0 <= io_in_write_entry_pfn_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_pfn_1 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_pfn_1 <= io_in_write_entry_pfn_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_c_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_c_0 <= io_in_write_entry_c_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_c_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_c_1 <= io_in_write_entry_c_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_d_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_d_0 <= io_in_write_entry_d_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_d_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_d_1 <= io_in_write_entry_d_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_v_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_v_0 <= io_in_write_entry_v_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_4_v_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h4 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_4_v_1 <= io_in_write_entry_v_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_vpn2 <= 19'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_vpn2 <= io_in_write_entry_vpn2; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_asid <= 8'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_asid <= io_in_write_entry_asid; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_g <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_g <= io_in_write_entry_g; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_pfn_0 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_pfn_0 <= io_in_write_entry_pfn_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_pfn_1 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_pfn_1 <= io_in_write_entry_pfn_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_c_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_c_0 <= io_in_write_entry_c_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_c_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_c_1 <= io_in_write_entry_c_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_d_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_d_0 <= io_in_write_entry_d_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_d_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_d_1 <= io_in_write_entry_d_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_v_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_v_0 <= io_in_write_entry_v_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_5_v_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h5 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_5_v_1 <= io_in_write_entry_v_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_vpn2 <= 19'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_vpn2 <= io_in_write_entry_vpn2; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_asid <= 8'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_asid <= io_in_write_entry_asid; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_g <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_g <= io_in_write_entry_g; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_pfn_0 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_pfn_0 <= io_in_write_entry_pfn_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_pfn_1 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_pfn_1 <= io_in_write_entry_pfn_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_c_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_c_0 <= io_in_write_entry_c_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_c_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_c_1 <= io_in_write_entry_c_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_d_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_d_0 <= io_in_write_entry_d_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_d_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_d_1 <= io_in_write_entry_d_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_v_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_v_0 <= io_in_write_entry_v_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_6_v_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h6 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_6_v_1 <= io_in_write_entry_v_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_vpn2 <= 19'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_vpn2 <= io_in_write_entry_vpn2; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_asid <= 8'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_asid <= io_in_write_entry_asid; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_g <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_g <= io_in_write_entry_g; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_pfn_0 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_pfn_0 <= io_in_write_entry_pfn_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_pfn_1 <= 20'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_pfn_1 <= io_in_write_entry_pfn_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_c_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_c_0 <= io_in_write_entry_c_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_c_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_c_1 <= io_in_write_entry_c_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_d_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_d_0 <= io_in_write_entry_d_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_d_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_d_1 <= io_in_write_entry_d_1; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_v_0 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_v_0 <= io_in_write_entry_v_0; // @[TlbL2.scala 66:31]
      end
    end
    if (reset) begin // @[TlbL2.scala 39:23]
      tlb_l2_7_v_1 <= 1'h0; // @[TlbL2.scala 39:23]
    end else if (io_in_write_en) begin // @[TlbL2.scala 65:24]
      if (3'h7 == io_in_write_index) begin // @[TlbL2.scala 66:31]
        tlb_l2_7_v_1 <= io_in_write_entry_v_1; // @[TlbL2.scala 66:31]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlb_l2_0_vpn2 = _RAND_0[18:0];
  _RAND_1 = {1{`RANDOM}};
  tlb_l2_0_asid = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  tlb_l2_0_g = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  tlb_l2_0_pfn_0 = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  tlb_l2_0_pfn_1 = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  tlb_l2_0_c_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  tlb_l2_0_c_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  tlb_l2_0_d_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tlb_l2_0_d_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  tlb_l2_0_v_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  tlb_l2_0_v_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tlb_l2_1_vpn2 = _RAND_11[18:0];
  _RAND_12 = {1{`RANDOM}};
  tlb_l2_1_asid = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  tlb_l2_1_g = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  tlb_l2_1_pfn_0 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  tlb_l2_1_pfn_1 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  tlb_l2_1_c_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  tlb_l2_1_c_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  tlb_l2_1_d_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  tlb_l2_1_d_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  tlb_l2_1_v_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  tlb_l2_1_v_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  tlb_l2_2_vpn2 = _RAND_22[18:0];
  _RAND_23 = {1{`RANDOM}};
  tlb_l2_2_asid = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  tlb_l2_2_g = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  tlb_l2_2_pfn_0 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  tlb_l2_2_pfn_1 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  tlb_l2_2_c_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  tlb_l2_2_c_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  tlb_l2_2_d_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  tlb_l2_2_d_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  tlb_l2_2_v_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  tlb_l2_2_v_1 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  tlb_l2_3_vpn2 = _RAND_33[18:0];
  _RAND_34 = {1{`RANDOM}};
  tlb_l2_3_asid = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  tlb_l2_3_g = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  tlb_l2_3_pfn_0 = _RAND_36[19:0];
  _RAND_37 = {1{`RANDOM}};
  tlb_l2_3_pfn_1 = _RAND_37[19:0];
  _RAND_38 = {1{`RANDOM}};
  tlb_l2_3_c_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  tlb_l2_3_c_1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  tlb_l2_3_d_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  tlb_l2_3_d_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  tlb_l2_3_v_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  tlb_l2_3_v_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tlb_l2_4_vpn2 = _RAND_44[18:0];
  _RAND_45 = {1{`RANDOM}};
  tlb_l2_4_asid = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  tlb_l2_4_g = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  tlb_l2_4_pfn_0 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  tlb_l2_4_pfn_1 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  tlb_l2_4_c_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  tlb_l2_4_c_1 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  tlb_l2_4_d_0 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  tlb_l2_4_d_1 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  tlb_l2_4_v_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  tlb_l2_4_v_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  tlb_l2_5_vpn2 = _RAND_55[18:0];
  _RAND_56 = {1{`RANDOM}};
  tlb_l2_5_asid = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  tlb_l2_5_g = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  tlb_l2_5_pfn_0 = _RAND_58[19:0];
  _RAND_59 = {1{`RANDOM}};
  tlb_l2_5_pfn_1 = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  tlb_l2_5_c_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  tlb_l2_5_c_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  tlb_l2_5_d_0 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  tlb_l2_5_d_1 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  tlb_l2_5_v_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tlb_l2_5_v_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  tlb_l2_6_vpn2 = _RAND_66[18:0];
  _RAND_67 = {1{`RANDOM}};
  tlb_l2_6_asid = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  tlb_l2_6_g = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  tlb_l2_6_pfn_0 = _RAND_69[19:0];
  _RAND_70 = {1{`RANDOM}};
  tlb_l2_6_pfn_1 = _RAND_70[19:0];
  _RAND_71 = {1{`RANDOM}};
  tlb_l2_6_c_0 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  tlb_l2_6_c_1 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  tlb_l2_6_d_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  tlb_l2_6_d_1 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  tlb_l2_6_v_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  tlb_l2_6_v_1 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  tlb_l2_7_vpn2 = _RAND_77[18:0];
  _RAND_78 = {1{`RANDOM}};
  tlb_l2_7_asid = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  tlb_l2_7_g = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  tlb_l2_7_pfn_0 = _RAND_80[19:0];
  _RAND_81 = {1{`RANDOM}};
  tlb_l2_7_pfn_1 = _RAND_81[19:0];
  _RAND_82 = {1{`RANDOM}};
  tlb_l2_7_c_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  tlb_l2_7_c_1 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  tlb_l2_7_d_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  tlb_l2_7_d_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  tlb_l2_7_v_0 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  tlb_l2_7_v_1 = _RAND_87[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cp0(
  input         clock,
  input         reset,
  input  [5:0]  io_ext_int,
  input         io_ctrl_exe_stall,
  input         io_ctrl_mem_stall,
  output        io_decoderUnit_access_allowed,
  output        io_decoderUnit_kernel_mode,
  output        io_decoderUnit_intterupt_allowed,
  output [7:0]  io_decoderUnit_cause_ip,
  output [7:0]  io_decoderUnit_status_im,
  input  [6:0]  io_executeUnit_in_inst_info_op,
  input  [7:0]  io_executeUnit_in_inst_info_cp0_addr,
  input  [31:0] io_executeUnit_in_mtc0_wdata,
  output [31:0] io_executeUnit_out_cp0_rdata,
  output [31:0] io_executeUnit_out_debug_cp0_count,
  output [31:0] io_executeUnit_out_debug_cp0_random,
  output [31:0] io_executeUnit_out_debug_cp0_cause,
  input  [31:0] io_memoryUnit_in_inst_0_pc,
  input         io_memoryUnit_in_inst_0_ex_flush_req,
  input         io_memoryUnit_in_inst_0_ex_tlb_refill,
  input         io_memoryUnit_in_inst_0_ex_eret,
  input  [31:0] io_memoryUnit_in_inst_0_ex_badvaddr,
  input         io_memoryUnit_in_inst_0_ex_bd,
  input  [4:0]  io_memoryUnit_in_inst_0_ex_excode,
  input  [31:0] io_memoryUnit_in_inst_1_pc,
  input         io_memoryUnit_in_inst_1_ex_flush_req,
  input         io_memoryUnit_in_inst_1_ex_tlb_refill,
  input         io_memoryUnit_in_inst_1_ex_eret,
  input  [31:0] io_memoryUnit_in_inst_1_ex_badvaddr,
  input         io_memoryUnit_in_inst_1_ex_bd,
  input  [4:0]  io_memoryUnit_in_inst_1_ex_excode,
  output        io_memoryUnit_out_flush,
  output [31:0] io_memoryUnit_out_flush_pc,
  input  [18:0] io_tlb_0_vpn2,
  output        io_tlb_0_found,
  output [19:0] io_tlb_0_info_pfn_0,
  output [19:0] io_tlb_0_info_pfn_1,
  output        io_tlb_0_info_c_0,
  output        io_tlb_0_info_c_1,
  output        io_tlb_0_info_v_0,
  output        io_tlb_0_info_v_1,
  input  [18:0] io_tlb_1_vpn2,
  output        io_tlb_1_found,
  output [19:0] io_tlb_1_info_pfn_0,
  output [19:0] io_tlb_1_info_pfn_1,
  output        io_tlb_1_info_c_0,
  output        io_tlb_1_info_c_1,
  output        io_tlb_1_info_d_0,
  output        io_tlb_1_info_d_1,
  output        io_tlb_1_info_v_0,
  output        io_tlb_1_info_v_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  wire  TlbL2_clock; // @[Cp0.scala 78:22]
  wire  TlbL2_reset; // @[Cp0.scala 78:22]
  wire  TlbL2_io_in_write_en; // @[Cp0.scala 78:22]
  wire [2:0] TlbL2_io_in_write_index; // @[Cp0.scala 78:22]
  wire [18:0] TlbL2_io_in_write_entry_vpn2; // @[Cp0.scala 78:22]
  wire [7:0] TlbL2_io_in_write_entry_asid; // @[Cp0.scala 78:22]
  wire  TlbL2_io_in_write_entry_g; // @[Cp0.scala 78:22]
  wire [19:0] TlbL2_io_in_write_entry_pfn_0; // @[Cp0.scala 78:22]
  wire [19:0] TlbL2_io_in_write_entry_pfn_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_in_write_entry_c_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_in_write_entry_c_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_in_write_entry_d_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_in_write_entry_d_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_in_write_entry_v_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_in_write_entry_v_1; // @[Cp0.scala 78:22]
  wire [2:0] TlbL2_io_in_read_index; // @[Cp0.scala 78:22]
  wire [18:0] TlbL2_io_in_entry_hi_vpn2; // @[Cp0.scala 78:22]
  wire [7:0] TlbL2_io_in_entry_hi_asid; // @[Cp0.scala 78:22]
  wire [18:0] TlbL2_io_in_tlb1_vpn2; // @[Cp0.scala 78:22]
  wire [18:0] TlbL2_io_in_tlb2_vpn2; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_read_entry_g; // @[Cp0.scala 78:22]
  wire [19:0] TlbL2_io_out_read_entry_pfn_0; // @[Cp0.scala 78:22]
  wire [19:0] TlbL2_io_out_read_entry_pfn_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_read_entry_c_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_read_entry_c_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_read_entry_d_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_read_entry_d_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_read_entry_v_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_read_entry_v_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb1_found; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb2_found; // @[Cp0.scala 78:22]
  wire [19:0] TlbL2_io_out_tlb1_entry_pfn_0; // @[Cp0.scala 78:22]
  wire [19:0] TlbL2_io_out_tlb1_entry_pfn_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb1_entry_c_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb1_entry_c_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb1_entry_v_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb1_entry_v_1; // @[Cp0.scala 78:22]
  wire [19:0] TlbL2_io_out_tlb2_entry_pfn_0; // @[Cp0.scala 78:22]
  wire [19:0] TlbL2_io_out_tlb2_entry_pfn_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb2_entry_c_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb2_entry_c_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb2_entry_d_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb2_entry_d_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb2_entry_v_0; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb2_entry_v_1; // @[Cp0.scala 78:22]
  wire  TlbL2_io_out_tlb_found; // @[Cp0.scala 78:22]
  wire [2:0] TlbL2_io_out_tlb_match_index; // @[Cp0.scala 78:22]
  wire [31:0] pc = io_memoryUnit_in_inst_0_ex_flush_req ? io_memoryUnit_in_inst_0_pc : io_memoryUnit_in_inst_1_pc; // @[Cp0.scala 69:23]
  wire  ex_flush_req = io_memoryUnit_in_inst_0_ex_flush_req ? io_memoryUnit_in_inst_0_ex_flush_req :
    io_memoryUnit_in_inst_1_ex_flush_req; // @[Cp0.scala 70:23]
  wire  ex_tlb_refill = io_memoryUnit_in_inst_0_ex_flush_req ? io_memoryUnit_in_inst_0_ex_tlb_refill :
    io_memoryUnit_in_inst_1_ex_tlb_refill; // @[Cp0.scala 70:23]
  wire  ex_eret = io_memoryUnit_in_inst_0_ex_flush_req ? io_memoryUnit_in_inst_0_ex_eret :
    io_memoryUnit_in_inst_1_ex_eret; // @[Cp0.scala 70:23]
  wire [31:0] ex_badvaddr = io_memoryUnit_in_inst_0_ex_flush_req ? io_memoryUnit_in_inst_0_ex_badvaddr :
    io_memoryUnit_in_inst_1_ex_badvaddr; // @[Cp0.scala 70:23]
  wire  ex_bd = io_memoryUnit_in_inst_0_ex_flush_req ? io_memoryUnit_in_inst_0_ex_bd : io_memoryUnit_in_inst_1_ex_bd; // @[Cp0.scala 70:23]
  wire [4:0] ex_excode = io_memoryUnit_in_inst_0_ex_flush_req ? io_memoryUnit_in_inst_0_ex_excode :
    io_memoryUnit_in_inst_1_ex_excode; // @[Cp0.scala 70:23]
  wire  mtc0_wen = io_executeUnit_in_inst_info_op == 7'h12; // @[Cp0.scala 71:51]
  reg  cp0_index_p; // @[Cp0.scala 90:26]
  reg [2:0] cp0_index_index; // @[Cp0.scala 90:26]
  reg [2:0] cp0_random_random; // @[Cp0.scala 96:27]
  reg [19:0] cp0_entrylo0_pfn; // @[Cp0.scala 99:29]
  reg [2:0] cp0_entrylo0_c; // @[Cp0.scala 99:29]
  reg  cp0_entrylo0_d; // @[Cp0.scala 99:29]
  reg  cp0_entrylo0_v; // @[Cp0.scala 99:29]
  reg  cp0_entrylo0_g; // @[Cp0.scala 99:29]
  reg [19:0] cp0_entrylo1_pfn; // @[Cp0.scala 102:29]
  reg [2:0] cp0_entrylo1_c; // @[Cp0.scala 102:29]
  reg  cp0_entrylo1_d; // @[Cp0.scala 102:29]
  reg  cp0_entrylo1_v; // @[Cp0.scala 102:29]
  reg  cp0_entrylo1_g; // @[Cp0.scala 102:29]
  reg [8:0] cp0_context_ptebase; // @[Cp0.scala 105:28]
  reg [18:0] cp0_context_badvpn2; // @[Cp0.scala 105:28]
  reg [2:0] cp0_wired_wired; // @[Cp0.scala 111:26]
  reg [31:0] cp0_badvaddr_badvaddr; // @[Cp0.scala 114:29]
  reg [31:0] cp0_count_count; // @[Cp0.scala 120:26]
  reg [18:0] cp0_entryhi_vpn2; // @[Cp0.scala 123:28]
  reg [7:0] cp0_entryhi_asid; // @[Cp0.scala 123:28]
  reg [31:0] cp0_compare_compare; // @[Cp0.scala 126:28]
  reg  cp0_status_cu0; // @[Cp0.scala 132:27]
  reg  cp0_status_bev; // @[Cp0.scala 132:27]
  reg [7:0] cp0_status_im; // @[Cp0.scala 132:27]
  reg  cp0_status_um; // @[Cp0.scala 132:27]
  reg  cp0_status_erl; // @[Cp0.scala 132:27]
  reg  cp0_status_exl; // @[Cp0.scala 132:27]
  reg  cp0_status_ie; // @[Cp0.scala 132:27]
  reg  cp0_cause_bd; // @[Cp0.scala 135:26]
  reg  cp0_cause_iv; // @[Cp0.scala 135:26]
  reg [7:0] cp0_cause_ip; // @[Cp0.scala 135:26]
  reg [4:0] cp0_cause_excode; // @[Cp0.scala 135:26]
  reg [31:0] cp0_epc_epc; // @[Cp0.scala 138:24]
  reg [17:0] cp0_ebase_ebase; // @[Cp0.scala 147:26]
  reg [31:0] cp0_taglo; // @[Cp0.scala 166:26]
  reg [31:0] cp0_taghi; // @[Cp0.scala 169:26]
  reg [31:0] cp0_error_epc_epc; // @[Cp0.scala 172:30]
  wire  _T = ~io_ctrl_exe_stall; // @[Cp0.scala 174:35]
  wire  _T_1 = io_executeUnit_in_inst_info_op == 7'h4a; // @[Cp0.scala 174:57]
  wire [2:0] _cp0_index_index_T_1 = TlbL2_io_out_tlb_found ? TlbL2_io_out_tlb_match_index : cp0_index_index; // @[Cp0.scala 196:29]
  wire [2:0] _cp0_random_random_T_2 = cp0_random_random - 3'h1; // @[Cp0.scala 202:103]
  wire [2:0] _cp0_random_random_T_3 = cp0_random_random == cp0_wired_wired ? 3'h7 : _cp0_random_random_T_2; // @[Cp0.scala 202:27]
  wire  wdata_g = io_executeUnit_in_mtc0_wdata[0]; // @[Cp0.scala 207:38]
  wire  wdata_v = io_executeUnit_in_mtc0_wdata[1]; // @[Cp0.scala 207:38]
  wire  wdata_d = io_executeUnit_in_mtc0_wdata[2]; // @[Cp0.scala 207:38]
  wire [2:0] wdata_c = io_executeUnit_in_mtc0_wdata[5:3]; // @[Cp0.scala 207:38]
  wire [19:0] wdata_pfn = io_executeUnit_in_mtc0_wdata[25:6]; // @[Cp0.scala 207:38]
  wire  _T_15 = io_executeUnit_in_inst_info_op == 7'h49; // @[Cp0.scala 213:23]
  wire [2:0] _cp0_entrylo0_c_T = {2'h1,TlbL2_io_out_read_entry_c_0}; // @[Cat.scala 33:92]
  wire [2:0] _cp0_entrylo1_c_T = {2'h1,TlbL2_io_out_read_entry_c_1}; // @[Cat.scala 33:92]
  wire  _T_20 = ~io_ctrl_mem_stall; // @[Cp0.scala 241:8]
  wire  _T_21 = ~io_ctrl_mem_stall & ex_flush_req; // @[Cp0.scala 241:19]
  wire  _T_22 = 5'h3 == ex_excode; // @[Cp0.scala 242:52]
  wire  _T_23 = 5'h4 == ex_excode; // @[Cp0.scala 242:52]
  wire  _T_24 = 5'h2 == ex_excode; // @[Cp0.scala 242:52]
  wire  _T_27 = 5'h3 == ex_excode | 5'h4 == ex_excode | 5'h2 == ex_excode; // @[Cp0.scala 242:52]
  wire  _T_36 = 5'h5 == ex_excode; // @[Cp0.scala 261:70]
  wire  _T_38 = 5'h6 == ex_excode; // @[Cp0.scala 261:70]
  reg  tick; // @[Cp0.scala 267:21]
  wire [31:0] _cp0_count_count_T_1 = cp0_count_count + 32'h1; // @[Cp0.scala 270:40]
  wire [31:0] _GEN_47 = tick ? _cp0_count_count_T_1 : cp0_count_count; // @[Cp0.scala 269:14 270:21 120:26]
  wire [7:0] wdata_2_asid = io_executeUnit_in_mtc0_wdata[7:0]; // @[Cp0.scala 285:38]
  wire [18:0] wdata_2_vpn2 = io_executeUnit_in_mtc0_wdata[31:13]; // @[Cp0.scala 285:38]
  wire  _T_61 = io_executeUnit_in_inst_info_cp0_addr == 8'h58; // @[Cp0.scala 293:32]
  wire  _GEN_60 = cp0_status_erl & cp0_status_exl; // @[Cp0.scala 300:26 132:27 303:22]
  wire  wdata_3_um = io_executeUnit_in_mtc0_wdata[4]; // @[Cp0.scala 309:38]
  wire [7:0] wdata_3_im = io_executeUnit_in_mtc0_wdata[15:8]; // @[Cp0.scala 309:38]
  wire  wdata_3_bev = io_executeUnit_in_mtc0_wdata[22]; // @[Cp0.scala 309:38]
  wire  wdata_3_cu0 = io_executeUnit_in_mtc0_wdata[28]; // @[Cp0.scala 309:38]
  wire  _GEN_61 = mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h60 ? wdata_3_cu0 : cp0_status_cu0; // @[Cp0.scala 308:53 310:22 132:27]
  wire  _GEN_62 = mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h60 ? wdata_g : cp0_status_ie; // @[Cp0.scala 308:53 311:22 132:27]
  wire  _GEN_63 = mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h60 ? wdata_v : cp0_status_exl; // @[Cp0.scala 308:53 312:22 132:27]
  wire  _GEN_64 = mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h60 ? wdata_d : cp0_status_erl; // @[Cp0.scala 308:53 313:22 132:27]
  wire  _GEN_65 = mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h60 ? wdata_3_um : cp0_status_um; // @[Cp0.scala 308:53 314:22 132:27]
  wire [7:0] _GEN_66 = mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h60 ? wdata_3_im : cp0_status_im; // @[Cp0.scala 308:53 315:22 132:27]
  wire  _GEN_67 = mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h60 ? wdata_3_bev : cp0_status_bev; // @[Cp0.scala 308:53 316:22 132:27]
  wire  _GEN_70 = _T ? _GEN_63 : cp0_status_exl; // @[Cp0.scala 307:26 132:27]
  wire  _GEN_74 = _T ? _GEN_67 : cp0_status_bev; // @[Cp0.scala 307:26 132:27]
  wire  _GEN_75 = _T_21 | _GEN_70; // @[Cp0.scala 305:42 306:20]
  wire  _GEN_81 = _T_21 ? cp0_status_bev : _GEN_74; // @[Cp0.scala 132:27 305:42]
  wire  _GEN_88 = _T_20 & ex_eret ? cp0_status_bev : _GEN_81; // @[Cp0.scala 132:27 299:31]
  wire  _cp0_cause_ip_T_4 = cp0_cause_ip[7] | cp0_compare_compare == cp0_count_count | io_ext_int[5]; // @[Cp0.scala 322:64]
  wire [7:0] _cp0_cause_ip_T_7 = {_cp0_cause_ip_T_4,io_ext_int[4:0],cp0_cause_ip[1:0]}; // @[Cat.scala 33:92]
  wire  _T_72 = ~cp0_status_exl; // @[Cp0.scala 327:10]
  wire [4:0] _cp0_cause_excode_T_1 = 5'h0 == ex_excode ? 5'h1f : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_3 = 5'h1 == ex_excode ? 5'h0 : _cp0_cause_excode_T_1; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_5 = _T_24 ? 5'h1 : _cp0_cause_excode_T_3; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_7 = _T_22 ? 5'h2 : _cp0_cause_excode_T_5; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_9 = _T_23 ? 5'h3 : _cp0_cause_excode_T_7; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_11 = _T_36 ? 5'h4 : _cp0_cause_excode_T_9; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_13 = _T_38 ? 5'h5 : _cp0_cause_excode_T_11; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_15 = 5'h7 == ex_excode ? 5'h8 : _cp0_cause_excode_T_13; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_17 = 5'h8 == ex_excode ? 5'h9 : _cp0_cause_excode_T_15; // @[Mux.scala 81:58]
  wire [4:0] _cp0_cause_excode_T_19 = 5'h9 == ex_excode ? 5'ha : _cp0_cause_excode_T_17; // @[Mux.scala 81:58]
  wire [7:0] _cp0_cause_ip_T_9 = {1'h0,cp0_cause_ip[6:0]}; // @[Cat.scala 33:92]
  wire  wdata_4_iv = io_executeUnit_in_mtc0_wdata[23]; // @[Cp0.scala 353:40]
  wire [7:0] _cp0_cause_ip_T_12 = {cp0_cause_ip[7:2],wdata_3_im[1:0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_90 = io_executeUnit_in_inst_info_cp0_addr == 8'h68 ? _cp0_cause_ip_T_12 : _cp0_cause_ip_T_7; // @[Cp0.scala 321:16 352:48 354:22]
  wire  _GEN_91 = io_executeUnit_in_inst_info_cp0_addr == 8'h68 ? wdata_4_iv : cp0_cause_iv; // @[Cp0.scala 352:48 358:22 135:26]
  wire [7:0] _GEN_92 = _T_61 ? _cp0_cause_ip_T_9 : _GEN_90; // @[Cp0.scala 350:44 351:22]
  wire  _GEN_93 = _T_61 ? cp0_cause_iv : _GEN_91; // @[Cp0.scala 135:26 350:44]
  wire [31:0] _cp0_epc_epc_T_1 = pc - 32'h4; // @[Cp0.scala 366:36]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T = {cp0_index_p,28'h0,cp0_index_index}; // @[Cp0.scala 406:45]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_1 = {29'h0,cp0_random_random}; // @[Cp0.scala 407:46]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_2 = {6'h0,cp0_entrylo0_pfn,cp0_entrylo0_c,cp0_entrylo0_d,cp0_entrylo0_v,
    cp0_entrylo0_g}; // @[Cp0.scala 408:48]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_3 = {6'h0,cp0_entrylo1_pfn,cp0_entrylo1_c,cp0_entrylo1_d,cp0_entrylo1_v,
    cp0_entrylo1_g}; // @[Cp0.scala 409:48]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_4 = {cp0_context_ptebase,cp0_context_badvpn2,4'h0}; // @[Cp0.scala 410:47]
  wire [30:0] _io_executeUnit_out_cp0_rdata_T_5 = {28'h0,cp0_wired_wired}; // @[Cp0.scala 412:45]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_6 = {cp0_entryhi_vpn2,5'h0,cp0_entryhi_asid}; // @[Cp0.scala 415:47]
  wire [7:0] io_executeUnit_out_cp0_rdata_lo_2 = {3'h0,cp0_status_um,1'h0,cp0_status_erl,cp0_status_exl,cp0_status_ie}; // @[Cp0.scala 417:46]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_7 = {3'h0,cp0_status_cu0,5'h0,cp0_status_bev,6'h0,cp0_status_im,
    io_executeUnit_out_cp0_rdata_lo_2}; // @[Cp0.scala 417:46]
  wire [15:0] io_executeUnit_out_cp0_rdata_lo_3 = {cp0_cause_ip,1'h0,cp0_cause_excode,2'h0}; // @[Cp0.scala 418:45]
  wire [15:0] io_executeUnit_out_cp0_rdata_hi_6 = {cp0_cause_bd,7'h0,cp0_cause_iv,7'h0}; // @[Cp0.scala 418:45]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_8 = {cp0_cause_bd,7'h0,cp0_cause_iv,7'h0,cp0_cause_ip,1'h0,
    cp0_cause_excode,2'h0}; // @[Cp0.scala 418:45]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_9 = {2'h2,cp0_ebase_ebase,12'h0}; // @[Cp0.scala 421:45]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_13 = 8'h0 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_15 = 8'h8 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T_1 : _io_executeUnit_out_cp0_rdata_T_13; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_17 = 8'h10 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T_2 : _io_executeUnit_out_cp0_rdata_T_15; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_19 = 8'h18 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T_3 : _io_executeUnit_out_cp0_rdata_T_17; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_21 = 8'h20 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T_4 : _io_executeUnit_out_cp0_rdata_T_19; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_23 = 8'h28 == io_executeUnit_in_inst_info_cp0_addr ? 32'h0 :
    _io_executeUnit_out_cp0_rdata_T_21; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_25 = 8'h30 == io_executeUnit_in_inst_info_cp0_addr ? {{1'd0},
    _io_executeUnit_out_cp0_rdata_T_5} : _io_executeUnit_out_cp0_rdata_T_23; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_27 = 8'h40 == io_executeUnit_in_inst_info_cp0_addr ? cp0_badvaddr_badvaddr
     : _io_executeUnit_out_cp0_rdata_T_25; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_29 = 8'h48 == io_executeUnit_in_inst_info_cp0_addr ? cp0_count_count :
    _io_executeUnit_out_cp0_rdata_T_27; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_31 = 8'h50 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T_6 : _io_executeUnit_out_cp0_rdata_T_29; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_33 = 8'h58 == io_executeUnit_in_inst_info_cp0_addr ? cp0_compare_compare
     : _io_executeUnit_out_cp0_rdata_T_31; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_35 = 8'h60 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T_7 : _io_executeUnit_out_cp0_rdata_T_33; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_37 = 8'h68 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T_8 : _io_executeUnit_out_cp0_rdata_T_35; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_39 = 8'h70 == io_executeUnit_in_inst_info_cp0_addr ? cp0_epc_epc :
    _io_executeUnit_out_cp0_rdata_T_37; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_41 = 8'h78 == io_executeUnit_in_inst_info_cp0_addr ? 32'h18003 :
    _io_executeUnit_out_cp0_rdata_T_39; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_43 = 8'h79 == io_executeUnit_in_inst_info_cp0_addr ?
    _io_executeUnit_out_cp0_rdata_T_9 : _io_executeUnit_out_cp0_rdata_T_41; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_45 = 8'h80 == io_executeUnit_in_inst_info_cp0_addr ? 32'h80000083 :
    _io_executeUnit_out_cp0_rdata_T_43; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_47 = 8'h81 == io_executeUnit_in_inst_info_cp0_addr ? 32'he291480 :
    _io_executeUnit_out_cp0_rdata_T_45; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_49 = 8'he0 == io_executeUnit_in_inst_info_cp0_addr ? cp0_taglo :
    _io_executeUnit_out_cp0_rdata_T_47; // @[Mux.scala 81:58]
  wire [31:0] _io_executeUnit_out_cp0_rdata_T_51 = 8'he8 == io_executeUnit_in_inst_info_cp0_addr ? cp0_taghi :
    _io_executeUnit_out_cp0_rdata_T_49; // @[Mux.scala 81:58]
  wire  _io_decoderUnit_kernel_mode_T_3 = ~ex_eret; // @[Cp0.scala 433:24]
  wire  _io_decoderUnit_kernel_mode_T_4 = cp0_status_erl & ~ex_eret; // @[Cp0.scala 433:21]
  wire  _io_decoderUnit_kernel_mode_T_5 = cp0_status_exl & ~(ex_eret & cp0_status_erl) | _io_decoderUnit_kernel_mode_T_4
    ; // @[Cp0.scala 432:82]
  wire  _io_decoderUnit_kernel_mode_T_6 = ~cp0_status_um; // @[Cp0.scala 434:5]
  wire  _io_decoderUnit_kernel_mode_T_7 = _io_decoderUnit_kernel_mode_T_5 | _io_decoderUnit_kernel_mode_T_6; // @[Cp0.scala 433:34]
  wire  _io_decoderUnit_kernel_mode_T_9 = ex_flush_req & _io_decoderUnit_kernel_mode_T_3; // @[Cp0.scala 435:19]
  wire [31:0] trap_base = cp0_status_bev ? 32'hbfc00200 : _io_executeUnit_out_cp0_rdata_T_9; // @[Cp0.scala 443:22]
  wire [31:0] _io_memoryUnit_out_flush_pc_T = cp0_status_erl ? cp0_error_epc_epc : cp0_epc_epc; // @[Cp0.scala 452:38]
  wire [31:0] _io_memoryUnit_out_flush_pc_T_2 = trap_base + 32'h180; // @[Cp0.scala 457:17]
  wire  _io_memoryUnit_out_flush_pc_T_6 = ex_excode == 5'h1 & cp0_cause_iv & ~cp0_status_bev; // @[Cp0.scala 459:46]
  wire [8:0] _io_memoryUnit_out_flush_pc_T_9 = ex_tlb_refill & ex_excode != 5'h1 ? 9'h0 : 9'h180; // @[Cp0.scala 461:12]
  wire [9:0] _io_memoryUnit_out_flush_pc_T_10 = _io_memoryUnit_out_flush_pc_T_6 ? 10'h200 : {{1'd0},
    _io_memoryUnit_out_flush_pc_T_9}; // @[Cp0.scala 458:22]
  wire [31:0] _GEN_118 = {{22'd0}, _io_memoryUnit_out_flush_pc_T_10}; // @[Cp0.scala 458:17]
  wire [31:0] _io_memoryUnit_out_flush_pc_T_12 = trap_base + _GEN_118; // @[Cp0.scala 458:17]
  wire [31:0] _io_memoryUnit_out_flush_pc_T_13 = cp0_status_exl ? _io_memoryUnit_out_flush_pc_T_2 :
    _io_memoryUnit_out_flush_pc_T_12; // @[Cp0.scala 455:38]
  wire  _GEN_114 = ex_flush_req & _T_20; // @[Cp0.scala 453:28 454:29 448:30]
  wire [31:0] _GEN_115 = ex_flush_req ? _io_memoryUnit_out_flush_pc_T_13 : 32'h0; // @[Cp0.scala 453:28 449:30 455:32]
  TlbL2 TlbL2 ( // @[Cp0.scala 78:22]
    .clock(TlbL2_clock),
    .reset(TlbL2_reset),
    .io_in_write_en(TlbL2_io_in_write_en),
    .io_in_write_index(TlbL2_io_in_write_index),
    .io_in_write_entry_vpn2(TlbL2_io_in_write_entry_vpn2),
    .io_in_write_entry_asid(TlbL2_io_in_write_entry_asid),
    .io_in_write_entry_g(TlbL2_io_in_write_entry_g),
    .io_in_write_entry_pfn_0(TlbL2_io_in_write_entry_pfn_0),
    .io_in_write_entry_pfn_1(TlbL2_io_in_write_entry_pfn_1),
    .io_in_write_entry_c_0(TlbL2_io_in_write_entry_c_0),
    .io_in_write_entry_c_1(TlbL2_io_in_write_entry_c_1),
    .io_in_write_entry_d_0(TlbL2_io_in_write_entry_d_0),
    .io_in_write_entry_d_1(TlbL2_io_in_write_entry_d_1),
    .io_in_write_entry_v_0(TlbL2_io_in_write_entry_v_0),
    .io_in_write_entry_v_1(TlbL2_io_in_write_entry_v_1),
    .io_in_read_index(TlbL2_io_in_read_index),
    .io_in_entry_hi_vpn2(TlbL2_io_in_entry_hi_vpn2),
    .io_in_entry_hi_asid(TlbL2_io_in_entry_hi_asid),
    .io_in_tlb1_vpn2(TlbL2_io_in_tlb1_vpn2),
    .io_in_tlb2_vpn2(TlbL2_io_in_tlb2_vpn2),
    .io_out_read_entry_g(TlbL2_io_out_read_entry_g),
    .io_out_read_entry_pfn_0(TlbL2_io_out_read_entry_pfn_0),
    .io_out_read_entry_pfn_1(TlbL2_io_out_read_entry_pfn_1),
    .io_out_read_entry_c_0(TlbL2_io_out_read_entry_c_0),
    .io_out_read_entry_c_1(TlbL2_io_out_read_entry_c_1),
    .io_out_read_entry_d_0(TlbL2_io_out_read_entry_d_0),
    .io_out_read_entry_d_1(TlbL2_io_out_read_entry_d_1),
    .io_out_read_entry_v_0(TlbL2_io_out_read_entry_v_0),
    .io_out_read_entry_v_1(TlbL2_io_out_read_entry_v_1),
    .io_out_tlb1_found(TlbL2_io_out_tlb1_found),
    .io_out_tlb2_found(TlbL2_io_out_tlb2_found),
    .io_out_tlb1_entry_pfn_0(TlbL2_io_out_tlb1_entry_pfn_0),
    .io_out_tlb1_entry_pfn_1(TlbL2_io_out_tlb1_entry_pfn_1),
    .io_out_tlb1_entry_c_0(TlbL2_io_out_tlb1_entry_c_0),
    .io_out_tlb1_entry_c_1(TlbL2_io_out_tlb1_entry_c_1),
    .io_out_tlb1_entry_v_0(TlbL2_io_out_tlb1_entry_v_0),
    .io_out_tlb1_entry_v_1(TlbL2_io_out_tlb1_entry_v_1),
    .io_out_tlb2_entry_pfn_0(TlbL2_io_out_tlb2_entry_pfn_0),
    .io_out_tlb2_entry_pfn_1(TlbL2_io_out_tlb2_entry_pfn_1),
    .io_out_tlb2_entry_c_0(TlbL2_io_out_tlb2_entry_c_0),
    .io_out_tlb2_entry_c_1(TlbL2_io_out_tlb2_entry_c_1),
    .io_out_tlb2_entry_d_0(TlbL2_io_out_tlb2_entry_d_0),
    .io_out_tlb2_entry_d_1(TlbL2_io_out_tlb2_entry_d_1),
    .io_out_tlb2_entry_v_0(TlbL2_io_out_tlb2_entry_v_0),
    .io_out_tlb2_entry_v_1(TlbL2_io_out_tlb2_entry_v_1),
    .io_out_tlb_found(TlbL2_io_out_tlb_found),
    .io_out_tlb_match_index(TlbL2_io_out_tlb_match_index)
  );
  assign io_decoderUnit_access_allowed = io_decoderUnit_kernel_mode | cp0_status_cu0; // @[Cp0.scala 436:66]
  assign io_decoderUnit_kernel_mode = _io_decoderUnit_kernel_mode_T_7 | _io_decoderUnit_kernel_mode_T_9; // @[Cp0.scala 434:20]
  assign io_decoderUnit_intterupt_allowed = cp0_status_ie & _T_72 & ~cp0_status_erl; // @[Cp0.scala 437:72]
  assign io_decoderUnit_cause_ip = cp0_cause_ip; // @[Cp0.scala 430:28]
  assign io_decoderUnit_status_im = cp0_status_im; // @[Cp0.scala 431:28]
  assign io_executeUnit_out_cp0_rdata = 8'hf0 == io_executeUnit_in_inst_info_cp0_addr ? cp0_error_epc_epc :
    _io_executeUnit_out_cp0_rdata_T_51; // @[Mux.scala 81:58]
  assign io_executeUnit_out_debug_cp0_count = cp0_count_count; // @[Cp0.scala 440:39]
  assign io_executeUnit_out_debug_cp0_random = {29'h0,cp0_random_random}; // @[Cp0.scala 441:59]
  assign io_executeUnit_out_debug_cp0_cause = {io_executeUnit_out_cp0_rdata_hi_6,io_executeUnit_out_cp0_rdata_lo_3}; // @[Cp0.scala 439:58]
  assign io_memoryUnit_out_flush = ex_eret ? _T_20 : _GEN_114; // @[Cp0.scala 450:17 451:32]
  assign io_memoryUnit_out_flush_pc = ex_eret ? _io_memoryUnit_out_flush_pc_T : _GEN_115; // @[Cp0.scala 450:17 452:32]
  assign io_tlb_0_found = TlbL2_io_out_tlb1_found; // @[Cp0.scala 82:23]
  assign io_tlb_0_info_pfn_0 = TlbL2_io_out_tlb1_entry_pfn_0; // @[Cp0.scala 84:23]
  assign io_tlb_0_info_pfn_1 = TlbL2_io_out_tlb1_entry_pfn_1; // @[Cp0.scala 84:23]
  assign io_tlb_0_info_c_0 = TlbL2_io_out_tlb1_entry_c_0; // @[Cp0.scala 84:23]
  assign io_tlb_0_info_c_1 = TlbL2_io_out_tlb1_entry_c_1; // @[Cp0.scala 84:23]
  assign io_tlb_0_info_v_0 = TlbL2_io_out_tlb1_entry_v_0; // @[Cp0.scala 84:23]
  assign io_tlb_0_info_v_1 = TlbL2_io_out_tlb1_entry_v_1; // @[Cp0.scala 84:23]
  assign io_tlb_1_found = TlbL2_io_out_tlb2_found; // @[Cp0.scala 83:23]
  assign io_tlb_1_info_pfn_0 = TlbL2_io_out_tlb2_entry_pfn_0; // @[Cp0.scala 85:23]
  assign io_tlb_1_info_pfn_1 = TlbL2_io_out_tlb2_entry_pfn_1; // @[Cp0.scala 85:23]
  assign io_tlb_1_info_c_0 = TlbL2_io_out_tlb2_entry_c_0; // @[Cp0.scala 85:23]
  assign io_tlb_1_info_c_1 = TlbL2_io_out_tlb2_entry_c_1; // @[Cp0.scala 85:23]
  assign io_tlb_1_info_d_0 = TlbL2_io_out_tlb2_entry_d_0; // @[Cp0.scala 85:23]
  assign io_tlb_1_info_d_1 = TlbL2_io_out_tlb2_entry_d_1; // @[Cp0.scala 85:23]
  assign io_tlb_1_info_v_0 = TlbL2_io_out_tlb2_entry_v_0; // @[Cp0.scala 85:23]
  assign io_tlb_1_info_v_1 = TlbL2_io_out_tlb2_entry_v_1; // @[Cp0.scala 85:23]
  assign TlbL2_clock = clock;
  assign TlbL2_reset = reset;
  assign TlbL2_io_in_write_en = ~io_ctrl_exe_stall & (io_executeUnit_in_inst_info_op == 7'h4a |
    io_executeUnit_in_inst_info_op == 7'h4b); // @[Cp0.scala 174:46]
  assign TlbL2_io_in_write_index = _T_1 ? cp0_index_index : cp0_random_random; // @[Cp0.scala 175:38]
  assign TlbL2_io_in_write_entry_vpn2 = cp0_entryhi_vpn2; // @[Cp0.scala 177:32]
  assign TlbL2_io_in_write_entry_asid = cp0_entryhi_asid; // @[Cp0.scala 176:32]
  assign TlbL2_io_in_write_entry_g = cp0_entrylo0_g | cp0_entrylo1_g; // @[Cp0.scala 178:50]
  assign TlbL2_io_in_write_entry_pfn_0 = cp0_entrylo0_pfn; // @[Cp0.scala 179:32]
  assign TlbL2_io_in_write_entry_pfn_1 = cp0_entrylo1_pfn; // @[Cp0.scala 180:32]
  assign TlbL2_io_in_write_entry_c_0 = cp0_entrylo0_c[0]; // @[Cp0.scala 181:32]
  assign TlbL2_io_in_write_entry_c_1 = cp0_entrylo1_c[0]; // @[Cp0.scala 182:32]
  assign TlbL2_io_in_write_entry_d_0 = cp0_entrylo0_d; // @[Cp0.scala 183:32]
  assign TlbL2_io_in_write_entry_d_1 = cp0_entrylo1_d; // @[Cp0.scala 184:32]
  assign TlbL2_io_in_write_entry_v_0 = cp0_entrylo0_v; // @[Cp0.scala 185:32]
  assign TlbL2_io_in_write_entry_v_1 = cp0_entrylo1_v; // @[Cp0.scala 186:32]
  assign TlbL2_io_in_read_index = cp0_index_index; // @[Cp0.scala 189:32]
  assign TlbL2_io_in_entry_hi_vpn2 = cp0_entryhi_vpn2; // @[Cp0.scala 188:32]
  assign TlbL2_io_in_entry_hi_asid = cp0_entryhi_asid; // @[Cp0.scala 187:32]
  assign TlbL2_io_in_tlb1_vpn2 = io_tlb_0_vpn2; // @[Cp0.scala 80:23]
  assign TlbL2_io_in_tlb2_vpn2 = io_tlb_1_vpn2; // @[Cp0.scala 81:23]
  always @(posedge clock) begin
    if (reset) begin // @[Cp0.scala 90:26]
      cp0_index_p <= 1'h0; // @[Cp0.scala 90:26]
    end else if (_T) begin // @[Cp0.scala 192:20]
      if (!(mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h0)) begin // @[Cp0.scala 193:52]
        if (io_executeUnit_in_inst_info_op == 7'h48) begin // @[Cp0.scala 195:37]
          cp0_index_p <= ~TlbL2_io_out_tlb_found; // @[Cp0.scala 197:23]
        end
      end
    end
    if (reset) begin // @[Cp0.scala 90:26]
      cp0_index_index <= 3'h0; // @[Cp0.scala 90:26]
    end else if (_T) begin // @[Cp0.scala 192:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h0) begin // @[Cp0.scala 193:52]
        cp0_index_index <= io_executeUnit_in_mtc0_wdata[2:0]; // @[Cp0.scala 194:23]
      end else if (io_executeUnit_in_inst_info_op == 7'h48) begin // @[Cp0.scala 195:37]
        cp0_index_index <= _cp0_index_index_T_1; // @[Cp0.scala 196:23]
      end
    end
    if (reset) begin // @[Cp0.scala 96:27]
      cp0_random_random <= 3'h7; // @[Cp0.scala 96:27]
    end else if (_T) begin // @[Cp0.scala 252:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h30) begin // @[Cp0.scala 253:52]
        cp0_random_random <= 3'h7; // @[Cp0.scala 255:25]
      end else begin
        cp0_random_random <= _cp0_random_random_T_3; // @[Cp0.scala 202:21]
      end
    end else begin
      cp0_random_random <= _cp0_random_random_T_3; // @[Cp0.scala 202:21]
    end
    if (reset) begin // @[Cp0.scala 99:29]
      cp0_entrylo0_pfn <= 20'h0; // @[Cp0.scala 99:29]
    end else if (_T) begin // @[Cp0.scala 205:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h10) begin // @[Cp0.scala 206:55]
        cp0_entrylo0_pfn <= wdata_pfn; // @[Cp0.scala 208:24]
      end else if (io_executeUnit_in_inst_info_op == 7'h49) begin // @[Cp0.scala 213:37]
        cp0_entrylo0_pfn <= TlbL2_io_out_read_entry_pfn_0; // @[Cp0.scala 214:24]
      end
    end
    if (reset) begin // @[Cp0.scala 99:29]
      cp0_entrylo0_c <= 3'h0; // @[Cp0.scala 99:29]
    end else if (_T) begin // @[Cp0.scala 205:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h10) begin // @[Cp0.scala 206:55]
        cp0_entrylo0_c <= wdata_c; // @[Cp0.scala 209:24]
      end else if (io_executeUnit_in_inst_info_op == 7'h49) begin // @[Cp0.scala 213:37]
        cp0_entrylo0_c <= _cp0_entrylo0_c_T; // @[Cp0.scala 216:24]
      end
    end
    if (reset) begin // @[Cp0.scala 99:29]
      cp0_entrylo0_d <= 1'h0; // @[Cp0.scala 99:29]
    end else if (_T) begin // @[Cp0.scala 205:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h10) begin // @[Cp0.scala 206:55]
        cp0_entrylo0_d <= wdata_d; // @[Cp0.scala 210:24]
      end else if (io_executeUnit_in_inst_info_op == 7'h49) begin // @[Cp0.scala 213:37]
        cp0_entrylo0_d <= TlbL2_io_out_read_entry_d_0; // @[Cp0.scala 217:24]
      end
    end
    if (reset) begin // @[Cp0.scala 99:29]
      cp0_entrylo0_v <= 1'h0; // @[Cp0.scala 99:29]
    end else if (_T) begin // @[Cp0.scala 205:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h10) begin // @[Cp0.scala 206:55]
        cp0_entrylo0_v <= wdata_v; // @[Cp0.scala 211:24]
      end else if (io_executeUnit_in_inst_info_op == 7'h49) begin // @[Cp0.scala 213:37]
        cp0_entrylo0_v <= TlbL2_io_out_read_entry_v_0; // @[Cp0.scala 218:24]
      end
    end
    if (reset) begin // @[Cp0.scala 99:29]
      cp0_entrylo0_g <= 1'h0; // @[Cp0.scala 99:29]
    end else if (_T) begin // @[Cp0.scala 205:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h10) begin // @[Cp0.scala 206:55]
        cp0_entrylo0_g <= wdata_g; // @[Cp0.scala 212:24]
      end else if (io_executeUnit_in_inst_info_op == 7'h49) begin // @[Cp0.scala 213:37]
        cp0_entrylo0_g <= TlbL2_io_out_read_entry_g; // @[Cp0.scala 215:24]
      end
    end
    if (reset) begin // @[Cp0.scala 102:29]
      cp0_entrylo1_pfn <= 20'h0; // @[Cp0.scala 102:29]
    end else if (_T) begin // @[Cp0.scala 223:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h18) begin // @[Cp0.scala 224:55]
        cp0_entrylo1_pfn <= wdata_pfn; // @[Cp0.scala 226:24]
      end else if (_T_15) begin // @[Cp0.scala 231:37]
        cp0_entrylo1_pfn <= TlbL2_io_out_read_entry_pfn_1; // @[Cp0.scala 232:24]
      end
    end
    if (reset) begin // @[Cp0.scala 102:29]
      cp0_entrylo1_c <= 3'h0; // @[Cp0.scala 102:29]
    end else if (_T) begin // @[Cp0.scala 223:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h18) begin // @[Cp0.scala 224:55]
        cp0_entrylo1_c <= wdata_c; // @[Cp0.scala 227:24]
      end else if (_T_15) begin // @[Cp0.scala 231:37]
        cp0_entrylo1_c <= _cp0_entrylo1_c_T; // @[Cp0.scala 234:24]
      end
    end
    if (reset) begin // @[Cp0.scala 102:29]
      cp0_entrylo1_d <= 1'h0; // @[Cp0.scala 102:29]
    end else if (_T) begin // @[Cp0.scala 223:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h18) begin // @[Cp0.scala 224:55]
        cp0_entrylo1_d <= wdata_d; // @[Cp0.scala 228:24]
      end else if (_T_15) begin // @[Cp0.scala 231:37]
        cp0_entrylo1_d <= TlbL2_io_out_read_entry_d_1; // @[Cp0.scala 235:24]
      end
    end
    if (reset) begin // @[Cp0.scala 102:29]
      cp0_entrylo1_v <= 1'h0; // @[Cp0.scala 102:29]
    end else if (_T) begin // @[Cp0.scala 223:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h18) begin // @[Cp0.scala 224:55]
        cp0_entrylo1_v <= wdata_v; // @[Cp0.scala 229:24]
      end else if (_T_15) begin // @[Cp0.scala 231:37]
        cp0_entrylo1_v <= TlbL2_io_out_read_entry_v_1; // @[Cp0.scala 236:24]
      end
    end
    if (reset) begin // @[Cp0.scala 102:29]
      cp0_entrylo1_g <= 1'h0; // @[Cp0.scala 102:29]
    end else if (_T) begin // @[Cp0.scala 223:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h18) begin // @[Cp0.scala 224:55]
        cp0_entrylo1_g <= wdata_g; // @[Cp0.scala 230:24]
      end else if (_T_15) begin // @[Cp0.scala 231:37]
        cp0_entrylo1_g <= TlbL2_io_out_read_entry_g; // @[Cp0.scala 233:24]
      end
    end
    if (reset) begin // @[Cp0.scala 105:28]
      cp0_context_ptebase <= 9'h0; // @[Cp0.scala 105:28]
    end else if (!(~io_ctrl_mem_stall & ex_flush_req)) begin // @[Cp0.scala 241:36]
      if (_T) begin // @[Cp0.scala 245:26]
        if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h20) begin // @[Cp0.scala 246:54]
          cp0_context_ptebase <= io_executeUnit_in_mtc0_wdata[31:23]; // @[Cp0.scala 247:27]
        end
      end
    end
    if (reset) begin // @[Cp0.scala 105:28]
      cp0_context_badvpn2 <= 19'h0; // @[Cp0.scala 105:28]
    end else if (~io_ctrl_mem_stall & ex_flush_req) begin // @[Cp0.scala 241:36]
      if (5'h3 == ex_excode | 5'h4 == ex_excode | 5'h2 == ex_excode) begin // @[Cp0.scala 242:65]
        cp0_context_badvpn2 <= ex_badvaddr[31:13]; // @[Cp0.scala 243:27]
      end
    end
    if (reset) begin // @[Cp0.scala 111:26]
      cp0_wired_wired <= 3'h0; // @[Cp0.scala 111:26]
    end else if (_T) begin // @[Cp0.scala 252:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h30) begin // @[Cp0.scala 253:52]
        cp0_wired_wired <= io_executeUnit_in_mtc0_wdata[2:0]; // @[Cp0.scala 254:25]
      end
    end
    if (reset) begin // @[Cp0.scala 114:29]
      cp0_badvaddr_badvaddr <= 32'h0; // @[Cp0.scala 114:29]
    end else if (_T_21) begin // @[Cp0.scala 260:36]
      if (5'h5 == ex_excode | _T_22 | 5'h6 == ex_excode | _T_23 | _T_24) begin // @[Cp0.scala 261:83]
        if (io_memoryUnit_in_inst_0_ex_flush_req) begin // @[Cp0.scala 70:23]
          cp0_badvaddr_badvaddr <= io_memoryUnit_in_inst_0_ex_badvaddr;
        end else begin
          cp0_badvaddr_badvaddr <= io_memoryUnit_in_inst_1_ex_badvaddr;
        end
      end
    end
    if (reset) begin // @[Cp0.scala 120:26]
      cp0_count_count <= 32'h1; // @[Cp0.scala 120:26]
    end else if (_T) begin // @[Cp0.scala 272:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h48) begin // @[Cp0.scala 273:52]
        cp0_count_count <= io_executeUnit_in_mtc0_wdata; // @[Cp0.scala 274:23]
      end else begin
        cp0_count_count <= _GEN_47;
      end
    end else begin
      cp0_count_count <= _GEN_47;
    end
    if (reset) begin // @[Cp0.scala 123:28]
      cp0_entryhi_vpn2 <= 19'h0; // @[Cp0.scala 123:28]
    end else if (_T_21) begin // @[Cp0.scala 279:36]
      if (_T_27) begin // @[Cp0.scala 280:65]
        cp0_entryhi_vpn2 <= ex_badvaddr[31:13]; // @[Cp0.scala 281:24]
      end
    end else if (_T) begin // @[Cp0.scala 283:26]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h50) begin // @[Cp0.scala 284:54]
        cp0_entryhi_vpn2 <= wdata_2_vpn2; // @[Cp0.scala 287:24]
      end
    end
    if (reset) begin // @[Cp0.scala 123:28]
      cp0_entryhi_asid <= 8'h0; // @[Cp0.scala 123:28]
    end else if (!(_T_21)) begin // @[Cp0.scala 279:36]
      if (_T) begin // @[Cp0.scala 283:26]
        if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h50) begin // @[Cp0.scala 284:54]
          cp0_entryhi_asid <= wdata_2_asid; // @[Cp0.scala 286:24]
        end
      end
    end
    if (reset) begin // @[Cp0.scala 126:28]
      cp0_compare_compare <= 32'h0; // @[Cp0.scala 126:28]
    end else if (_T) begin // @[Cp0.scala 292:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h58) begin // @[Cp0.scala 293:54]
        cp0_compare_compare <= io_executeUnit_in_mtc0_wdata; // @[Cp0.scala 294:27]
      end
    end
    if (reset) begin // @[Cp0.scala 132:27]
      cp0_status_cu0 <= 1'h0; // @[Cp0.scala 132:27]
    end else if (!(_T_20 & ex_eret)) begin // @[Cp0.scala 299:31]
      if (!(_T_21)) begin // @[Cp0.scala 305:42]
        if (_T) begin // @[Cp0.scala 307:26]
          cp0_status_cu0 <= _GEN_61;
        end
      end
    end
    cp0_status_bev <= reset | _GEN_88; // @[Cp0.scala 132:{27,27}]
    if (reset) begin // @[Cp0.scala 132:27]
      cp0_status_im <= 8'h0; // @[Cp0.scala 132:27]
    end else if (!(_T_20 & ex_eret)) begin // @[Cp0.scala 299:31]
      if (!(_T_21)) begin // @[Cp0.scala 305:42]
        if (_T) begin // @[Cp0.scala 307:26]
          cp0_status_im <= _GEN_66;
        end
      end
    end
    if (reset) begin // @[Cp0.scala 132:27]
      cp0_status_um <= 1'h0; // @[Cp0.scala 132:27]
    end else if (!(_T_20 & ex_eret)) begin // @[Cp0.scala 299:31]
      if (!(_T_21)) begin // @[Cp0.scala 305:42]
        if (_T) begin // @[Cp0.scala 307:26]
          cp0_status_um <= _GEN_65;
        end
      end
    end
    if (reset) begin // @[Cp0.scala 132:27]
      cp0_status_erl <= 1'h0; // @[Cp0.scala 132:27]
    end else if (_T_20 & ex_eret) begin // @[Cp0.scala 299:31]
      if (cp0_status_erl) begin // @[Cp0.scala 300:26]
        cp0_status_erl <= 1'h0; // @[Cp0.scala 301:22]
      end
    end else if (!(_T_21)) begin // @[Cp0.scala 305:42]
      if (_T) begin // @[Cp0.scala 307:26]
        cp0_status_erl <= _GEN_64;
      end
    end
    if (reset) begin // @[Cp0.scala 132:27]
      cp0_status_exl <= 1'h0; // @[Cp0.scala 132:27]
    end else if (_T_20 & ex_eret) begin // @[Cp0.scala 299:31]
      cp0_status_exl <= _GEN_60;
    end else begin
      cp0_status_exl <= _GEN_75;
    end
    if (reset) begin // @[Cp0.scala 132:27]
      cp0_status_ie <= 1'h0; // @[Cp0.scala 132:27]
    end else if (!(_T_20 & ex_eret)) begin // @[Cp0.scala 299:31]
      if (!(_T_21)) begin // @[Cp0.scala 305:42]
        if (_T) begin // @[Cp0.scala 307:26]
          cp0_status_ie <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[Cp0.scala 135:26]
      cp0_cause_bd <= 1'h0; // @[Cp0.scala 135:26]
    end else if (_T_21) begin // @[Cp0.scala 326:36]
      if (~cp0_status_exl) begin // @[Cp0.scala 327:27]
        if (io_memoryUnit_in_inst_0_ex_flush_req) begin // @[Cp0.scala 70:23]
          cp0_cause_bd <= io_memoryUnit_in_inst_0_ex_bd;
        end else begin
          cp0_cause_bd <= io_memoryUnit_in_inst_1_ex_bd;
        end
      end
    end
    if (reset) begin // @[Cp0.scala 135:26]
      cp0_cause_iv <= 1'h0; // @[Cp0.scala 135:26]
    end else if (!(_T_21)) begin // @[Cp0.scala 326:36]
      if (_T) begin // @[Cp0.scala 348:26]
        if (mtc0_wen) begin // @[Cp0.scala 349:20]
          cp0_cause_iv <= _GEN_93;
        end
      end
    end
    if (reset) begin // @[Cp0.scala 135:26]
      cp0_cause_ip <= 8'h0; // @[Cp0.scala 135:26]
    end else if (_T_21) begin // @[Cp0.scala 326:36]
      cp0_cause_ip <= _cp0_cause_ip_T_7; // @[Cp0.scala 321:16]
    end else if (_T) begin // @[Cp0.scala 348:26]
      if (mtc0_wen) begin // @[Cp0.scala 349:20]
        cp0_cause_ip <= _GEN_92;
      end else begin
        cp0_cause_ip <= _cp0_cause_ip_T_7; // @[Cp0.scala 321:16]
      end
    end else begin
      cp0_cause_ip <= _cp0_cause_ip_T_7; // @[Cp0.scala 321:16]
    end
    if (reset) begin // @[Cp0.scala 135:26]
      cp0_cause_excode <= 5'h0; // @[Cp0.scala 135:26]
    end else if (_T_21) begin // @[Cp0.scala 326:36]
      if (5'hb == ex_excode) begin // @[Mux.scala 81:58]
        cp0_cause_excode <= 5'hc;
      end else if (5'ha == ex_excode) begin // @[Mux.scala 81:58]
        cp0_cause_excode <= 5'hb;
      end else begin
        cp0_cause_excode <= _cp0_cause_excode_T_19;
      end
    end
    if (reset) begin // @[Cp0.scala 138:24]
      cp0_epc_epc <= 32'h0; // @[Cp0.scala 138:24]
    end else if (_T_21) begin // @[Cp0.scala 364:36]
      if (_T_72) begin // @[Cp0.scala 365:27]
        if (ex_bd) begin // @[Cp0.scala 366:25]
          cp0_epc_epc <= _cp0_epc_epc_T_1;
        end else begin
          cp0_epc_epc <= pc;
        end
      end
    end else if (_T) begin // @[Cp0.scala 368:26]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h70) begin // @[Cp0.scala 369:50]
        cp0_epc_epc <= io_executeUnit_in_mtc0_wdata; // @[Cp0.scala 370:19]
      end
    end
    if (reset) begin // @[Cp0.scala 147:26]
      cp0_ebase_ebase <= 18'h0; // @[Cp0.scala 147:26]
    end else if (_T) begin // @[Cp0.scala 375:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'h79) begin // @[Cp0.scala 376:52]
        cp0_ebase_ebase <= io_executeUnit_in_mtc0_wdata[29:12]; // @[Cp0.scala 377:23]
      end
    end
    if (reset) begin // @[Cp0.scala 166:26]
      cp0_taglo <= 32'h0; // @[Cp0.scala 166:26]
    end else if (_T) begin // @[Cp0.scala 382:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'he0) begin // @[Cp0.scala 383:52]
        cp0_taglo <= io_executeUnit_in_mtc0_wdata; // @[Cp0.scala 384:17]
      end
    end
    if (reset) begin // @[Cp0.scala 169:26]
      cp0_taghi <= 32'h0; // @[Cp0.scala 169:26]
    end else if (_T) begin // @[Cp0.scala 389:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'he8) begin // @[Cp0.scala 390:52]
        cp0_taghi <= io_executeUnit_in_mtc0_wdata; // @[Cp0.scala 391:17]
      end
    end
    if (reset) begin // @[Cp0.scala 172:30]
      cp0_error_epc_epc <= 32'h0; // @[Cp0.scala 172:30]
    end else if (_T) begin // @[Cp0.scala 396:20]
      if (mtc0_wen & io_executeUnit_in_inst_info_cp0_addr == 8'hf0) begin // @[Cp0.scala 397:56]
        cp0_error_epc_epc <= io_executeUnit_in_mtc0_wdata; // @[Cp0.scala 398:25]
      end
    end
    if (reset) begin // @[Cp0.scala 267:21]
      tick <= 1'h0; // @[Cp0.scala 267:21]
    end else begin
      tick <= ~tick; // @[Cp0.scala 268:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cp0_index_p = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cp0_index_index = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  cp0_random_random = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  cp0_entrylo0_pfn = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  cp0_entrylo0_c = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  cp0_entrylo0_d = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  cp0_entrylo0_v = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cp0_entrylo0_g = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cp0_entrylo1_pfn = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  cp0_entrylo1_c = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  cp0_entrylo1_d = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cp0_entrylo1_v = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  cp0_entrylo1_g = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  cp0_context_ptebase = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  cp0_context_badvpn2 = _RAND_14[18:0];
  _RAND_15 = {1{`RANDOM}};
  cp0_wired_wired = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  cp0_badvaddr_badvaddr = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  cp0_count_count = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  cp0_entryhi_vpn2 = _RAND_18[18:0];
  _RAND_19 = {1{`RANDOM}};
  cp0_entryhi_asid = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  cp0_compare_compare = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  cp0_status_cu0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  cp0_status_bev = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  cp0_status_im = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  cp0_status_um = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  cp0_status_erl = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  cp0_status_exl = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  cp0_status_ie = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  cp0_cause_bd = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  cp0_cause_iv = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  cp0_cause_ip = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  cp0_cause_excode = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  cp0_epc_epc = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  cp0_ebase_ebase = _RAND_33[17:0];
  _RAND_34 = {1{`RANDOM}};
  cp0_taglo = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  cp0_taghi = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  cp0_error_epc_epc = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  tick = _RAND_37[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemoryStage(
  input         clock,
  input         reset,
  input         io_ctrl_allow_to_go,
  input         io_ctrl_clear_0,
  input         io_ctrl_clear_1,
  input  [31:0] io_executeUnit_inst0_pc,
  input  [3:0]  io_executeUnit_inst0_inst_info_fusel,
  input  [6:0]  io_executeUnit_inst0_inst_info_op,
  input         io_executeUnit_inst0_inst_info_reg_wen,
  input  [4:0]  io_executeUnit_inst0_inst_info_reg_waddr,
  input  [31:0] io_executeUnit_inst0_inst_info_inst,
  input  [31:0] io_executeUnit_inst0_rd_info_wdata,
  input         io_executeUnit_inst0_ex_flush_req,
  input         io_executeUnit_inst0_ex_eret,
  input  [31:0] io_executeUnit_inst0_ex_badvaddr,
  input         io_executeUnit_inst0_ex_bd,
  input  [4:0]  io_executeUnit_inst0_ex_excode,
  input  [31:0] io_executeUnit_inst0_cp0_cp0_count,
  input  [31:0] io_executeUnit_inst0_cp0_cp0_random,
  input  [31:0] io_executeUnit_inst0_cp0_cp0_cause,
  input         io_executeUnit_inst0_mem_en,
  input  [6:0]  io_executeUnit_inst0_mem_inst_info_op,
  input  [31:0] io_executeUnit_inst0_mem_addr,
  input  [31:0] io_executeUnit_inst0_mem_wdata,
  input         io_executeUnit_inst0_mem_sel_0,
  input         io_executeUnit_inst0_mem_sel_1,
  input  [31:0] io_executeUnit_inst1_pc,
  input  [3:0]  io_executeUnit_inst1_inst_info_fusel,
  input         io_executeUnit_inst1_inst_info_reg_wen,
  input  [4:0]  io_executeUnit_inst1_inst_info_reg_waddr,
  input  [31:0] io_executeUnit_inst1_rd_info_wdata,
  input         io_executeUnit_inst1_ex_flush_req,
  input         io_executeUnit_inst1_ex_eret,
  input  [31:0] io_executeUnit_inst1_ex_badvaddr,
  input         io_executeUnit_inst1_ex_bd,
  input  [4:0]  io_executeUnit_inst1_ex_excode,
  output [31:0] io_memoryUnit_inst0_pc,
  output [3:0]  io_memoryUnit_inst0_inst_info_fusel,
  output [6:0]  io_memoryUnit_inst0_inst_info_op,
  output        io_memoryUnit_inst0_inst_info_reg_wen,
  output [4:0]  io_memoryUnit_inst0_inst_info_reg_waddr,
  output [31:0] io_memoryUnit_inst0_inst_info_inst,
  output [31:0] io_memoryUnit_inst0_rd_info_wdata,
  output        io_memoryUnit_inst0_ex_flush_req,
  output        io_memoryUnit_inst0_ex_eret,
  output [31:0] io_memoryUnit_inst0_ex_badvaddr,
  output        io_memoryUnit_inst0_ex_bd,
  output [4:0]  io_memoryUnit_inst0_ex_excode,
  output [31:0] io_memoryUnit_inst0_cp0_cp0_count,
  output [31:0] io_memoryUnit_inst0_cp0_cp0_random,
  output [31:0] io_memoryUnit_inst0_cp0_cp0_cause,
  output        io_memoryUnit_inst0_mem_en,
  output [6:0]  io_memoryUnit_inst0_mem_inst_info_op,
  output [31:0] io_memoryUnit_inst0_mem_addr,
  output [31:0] io_memoryUnit_inst0_mem_wdata,
  output        io_memoryUnit_inst0_mem_sel_0,
  output        io_memoryUnit_inst0_mem_sel_1,
  output [31:0] io_memoryUnit_inst1_pc,
  output [3:0]  io_memoryUnit_inst1_inst_info_fusel,
  output        io_memoryUnit_inst1_inst_info_reg_wen,
  output [4:0]  io_memoryUnit_inst1_inst_info_reg_waddr,
  output [31:0] io_memoryUnit_inst1_rd_info_wdata,
  output        io_memoryUnit_inst1_ex_flush_req,
  output        io_memoryUnit_inst1_ex_eret,
  output [31:0] io_memoryUnit_inst1_ex_badvaddr,
  output        io_memoryUnit_inst1_ex_bd,
  output [4:0]  io_memoryUnit_inst1_ex_excode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] inst0_pc; // @[MemoryStage.scala 50:22]
  reg [3:0] inst0_inst_info_fusel; // @[MemoryStage.scala 50:22]
  reg [6:0] inst0_inst_info_op; // @[MemoryStage.scala 50:22]
  reg  inst0_inst_info_reg_wen; // @[MemoryStage.scala 50:22]
  reg [4:0] inst0_inst_info_reg_waddr; // @[MemoryStage.scala 50:22]
  reg [31:0] inst0_inst_info_inst; // @[MemoryStage.scala 50:22]
  reg [31:0] inst0_rd_info_wdata; // @[MemoryStage.scala 50:22]
  reg  inst0_ex_flush_req; // @[MemoryStage.scala 50:22]
  reg  inst0_ex_eret; // @[MemoryStage.scala 50:22]
  reg [31:0] inst0_ex_badvaddr; // @[MemoryStage.scala 50:22]
  reg  inst0_ex_bd; // @[MemoryStage.scala 50:22]
  reg [4:0] inst0_ex_excode; // @[MemoryStage.scala 50:22]
  reg [31:0] inst0_cp0_cp0_count; // @[MemoryStage.scala 50:22]
  reg [31:0] inst0_cp0_cp0_random; // @[MemoryStage.scala 50:22]
  reg [31:0] inst0_cp0_cp0_cause; // @[MemoryStage.scala 50:22]
  reg  inst0_mem_en; // @[MemoryStage.scala 50:22]
  reg [6:0] inst0_mem_inst_info_op; // @[MemoryStage.scala 50:22]
  reg [31:0] inst0_mem_addr; // @[MemoryStage.scala 50:22]
  reg [31:0] inst0_mem_wdata; // @[MemoryStage.scala 50:22]
  reg  inst0_mem_sel_0; // @[MemoryStage.scala 50:22]
  reg  inst0_mem_sel_1; // @[MemoryStage.scala 50:22]
  reg [31:0] inst1_pc; // @[MemoryStage.scala 51:22]
  reg [3:0] inst1_inst_info_fusel; // @[MemoryStage.scala 51:22]
  reg  inst1_inst_info_reg_wen; // @[MemoryStage.scala 51:22]
  reg [4:0] inst1_inst_info_reg_waddr; // @[MemoryStage.scala 51:22]
  reg [31:0] inst1_rd_info_wdata; // @[MemoryStage.scala 51:22]
  reg  inst1_ex_flush_req; // @[MemoryStage.scala 51:22]
  reg  inst1_ex_eret; // @[MemoryStage.scala 51:22]
  reg [31:0] inst1_ex_badvaddr; // @[MemoryStage.scala 51:22]
  reg  inst1_ex_bd; // @[MemoryStage.scala 51:22]
  reg [4:0] inst1_ex_excode; // @[MemoryStage.scala 51:22]
  assign io_memoryUnit_inst0_pc = inst0_pc; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_inst_info_fusel = inst0_inst_info_fusel; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_inst_info_op = inst0_inst_info_op; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_inst_info_reg_wen = inst0_inst_info_reg_wen; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_inst_info_reg_waddr = inst0_inst_info_reg_waddr; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_inst_info_inst = inst0_inst_info_inst; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_rd_info_wdata = inst0_rd_info_wdata; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_ex_flush_req = inst0_ex_flush_req; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_ex_eret = inst0_ex_eret; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_ex_badvaddr = inst0_ex_badvaddr; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_ex_bd = inst0_ex_bd; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_ex_excode = inst0_ex_excode; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_cp0_cp0_count = inst0_cp0_cp0_count; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_cp0_cp0_random = inst0_cp0_cp0_random; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_cp0_cp0_cause = inst0_cp0_cp0_cause; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_mem_en = inst0_mem_en; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_mem_inst_info_op = inst0_mem_inst_info_op; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_mem_addr = inst0_mem_addr; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_mem_wdata = inst0_mem_wdata; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_mem_sel_0 = inst0_mem_sel_0; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst0_mem_sel_1 = inst0_mem_sel_1; // @[MemoryStage.scala 65:23]
  assign io_memoryUnit_inst1_pc = inst1_pc; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_inst_info_fusel = inst1_inst_info_fusel; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_inst_info_reg_wen = inst1_inst_info_reg_wen; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_inst_info_reg_waddr = inst1_inst_info_reg_waddr; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_rd_info_wdata = inst1_rd_info_wdata; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_ex_flush_req = inst1_ex_flush_req; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_ex_eret = inst1_ex_eret; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_ex_badvaddr = inst1_ex_badvaddr; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_ex_bd = inst1_ex_bd; // @[MemoryStage.scala 66:23]
  assign io_memoryUnit_inst1_ex_excode = inst1_ex_excode; // @[MemoryStage.scala 66:23]
  always @(posedge clock) begin
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_pc <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_pc <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_pc <= io_executeUnit_inst0_pc; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_inst_info_fusel <= 4'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_inst_info_fusel <= 4'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_inst_info_fusel <= io_executeUnit_inst0_inst_info_fusel; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_inst_info_op <= 7'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_inst_info_op <= 7'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_inst_info_op <= io_executeUnit_inst0_inst_info_op; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_inst_info_reg_wen <= 1'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_inst_info_reg_wen <= 1'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_inst_info_reg_wen <= io_executeUnit_inst0_inst_info_reg_wen; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_inst_info_reg_waddr <= 5'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_inst_info_reg_waddr <= 5'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_inst_info_reg_waddr <= io_executeUnit_inst0_inst_info_reg_waddr; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_inst_info_inst <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_inst_info_inst <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_inst_info_inst <= io_executeUnit_inst0_inst_info_inst; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_rd_info_wdata <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_rd_info_wdata <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_rd_info_wdata <= io_executeUnit_inst0_rd_info_wdata; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_ex_flush_req <= 1'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_ex_flush_req <= 1'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_ex_flush_req <= io_executeUnit_inst0_ex_flush_req; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_ex_eret <= 1'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_ex_eret <= 1'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_ex_eret <= io_executeUnit_inst0_ex_eret; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_ex_badvaddr <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_ex_badvaddr <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_ex_badvaddr <= io_executeUnit_inst0_ex_badvaddr; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_ex_bd <= 1'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_ex_bd <= 1'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_ex_bd <= io_executeUnit_inst0_ex_bd; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_ex_excode <= 5'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_ex_excode <= 5'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_ex_excode <= io_executeUnit_inst0_ex_excode; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_cp0_cp0_count <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_cp0_cp0_count <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_cp0_cp0_count <= io_executeUnit_inst0_cp0_cp0_count; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_cp0_cp0_random <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_cp0_cp0_random <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_cp0_cp0_random <= io_executeUnit_inst0_cp0_cp0_random; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_cp0_cp0_cause <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_cp0_cp0_cause <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_cp0_cp0_cause <= io_executeUnit_inst0_cp0_cp0_cause; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_mem_en <= 1'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_mem_en <= 1'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_mem_en <= io_executeUnit_inst0_mem_en; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_mem_inst_info_op <= 7'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_mem_inst_info_op <= 7'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_mem_inst_info_op <= io_executeUnit_inst0_mem_inst_info_op; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_mem_addr <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_mem_addr <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_mem_addr <= io_executeUnit_inst0_mem_addr; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_mem_wdata <= 32'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_mem_wdata <= 32'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_mem_wdata <= io_executeUnit_inst0_mem_wdata; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_mem_sel_0 <= 1'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_mem_sel_0 <= 1'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_mem_sel_0 <= io_executeUnit_inst0_mem_sel_0; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 50:22]
      inst0_mem_sel_1 <= 1'h0; // @[MemoryStage.scala 50:22]
    end else if (io_ctrl_clear_0) begin // @[MemoryStage.scala 53:26]
      inst0_mem_sel_1 <= 1'h0; // @[MemoryStage.scala 54:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 55:35]
      inst0_mem_sel_1 <= io_executeUnit_inst0_mem_sel_1; // @[MemoryStage.scala 56:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_pc <= 32'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_pc <= 32'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_pc <= io_executeUnit_inst1_pc; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_inst_info_fusel <= 4'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_inst_info_fusel <= 4'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_inst_info_fusel <= io_executeUnit_inst1_inst_info_fusel; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_inst_info_reg_wen <= 1'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_inst_info_reg_wen <= 1'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_inst_info_reg_wen <= io_executeUnit_inst1_inst_info_reg_wen; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_inst_info_reg_waddr <= 5'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_inst_info_reg_waddr <= 5'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_inst_info_reg_waddr <= io_executeUnit_inst1_inst_info_reg_waddr; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_rd_info_wdata <= 32'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_rd_info_wdata <= 32'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_rd_info_wdata <= io_executeUnit_inst1_rd_info_wdata; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_ex_flush_req <= 1'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_ex_flush_req <= 1'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_ex_flush_req <= io_executeUnit_inst1_ex_flush_req; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_ex_eret <= 1'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_ex_eret <= 1'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_ex_eret <= io_executeUnit_inst1_ex_eret; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_ex_badvaddr <= 32'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_ex_badvaddr <= 32'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_ex_badvaddr <= io_executeUnit_inst1_ex_badvaddr; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_ex_bd <= 1'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_ex_bd <= 1'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_ex_bd <= io_executeUnit_inst1_ex_bd; // @[MemoryStage.scala 62:11]
    end
    if (reset) begin // @[MemoryStage.scala 51:22]
      inst1_ex_excode <= 5'h0; // @[MemoryStage.scala 51:22]
    end else if (io_ctrl_clear_1) begin // @[MemoryStage.scala 59:26]
      inst1_ex_excode <= 5'h0; // @[MemoryStage.scala 60:11]
    end else if (io_ctrl_allow_to_go) begin // @[MemoryStage.scala 61:35]
      inst1_ex_excode <= io_executeUnit_inst1_ex_excode; // @[MemoryStage.scala 62:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst0_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  inst0_inst_info_fusel = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  inst0_inst_info_op = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  inst0_inst_info_reg_wen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  inst0_inst_info_reg_waddr = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  inst0_inst_info_inst = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  inst0_rd_info_wdata = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  inst0_ex_flush_req = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  inst0_ex_eret = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  inst0_ex_badvaddr = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  inst0_ex_bd = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inst0_ex_excode = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  inst0_cp0_cp0_count = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  inst0_cp0_cp0_random = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  inst0_cp0_cp0_cause = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  inst0_mem_en = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  inst0_mem_inst_info_op = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  inst0_mem_addr = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  inst0_mem_wdata = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inst0_mem_sel_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  inst0_mem_sel_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  inst1_pc = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  inst1_inst_info_fusel = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  inst1_inst_info_reg_wen = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  inst1_inst_info_reg_waddr = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  inst1_rd_info_wdata = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  inst1_ex_flush_req = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  inst1_ex_eret = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  inst1_ex_badvaddr = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inst1_ex_bd = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  inst1_ex_excode = _RAND_30[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DataMemoryAccess(
  input         io_memoryUnit_in_mem_en,
  input  [6:0]  io_memoryUnit_in_inst_info_op,
  input  [31:0] io_memoryUnit_in_mem_wdata,
  input  [31:0] io_memoryUnit_in_mem_addr,
  input         io_memoryUnit_in_mem_sel_0,
  input         io_memoryUnit_in_mem_sel_1,
  input         io_memoryUnit_in_ex_0_flush_req,
  input         io_memoryUnit_in_ex_1_flush_req,
  output [31:0] io_memoryUnit_out_rdata,
  input  [31:0] io_dataMemory_in_rdata,
  output        io_dataMemory_out_en,
  output [1:0]  io_dataMemory_out_rlen,
  output [3:0]  io_dataMemory_out_wen,
  output [31:0] io_dataMemory_out_wdata
);
  wire [1:0] mem_addr2 = io_memoryUnit_in_mem_addr[1:0]; // @[DataMemoryAccess.scala 39:27]
  wire  _io_dataMemory_out_en_T = ~io_memoryUnit_in_ex_0_flush_req; // @[DataMemoryAccess.scala 44:37]
  wire  _io_dataMemory_out_en_T_5 = io_memoryUnit_in_mem_sel_1 & _io_dataMemory_out_en_T & ~
    io_memoryUnit_in_ex_1_flush_req; // @[DataMemoryAccess.scala 45:72]
  wire  _io_dataMemory_out_en_T_6 = io_memoryUnit_in_mem_sel_0 & ~io_memoryUnit_in_ex_0_flush_req |
    _io_dataMemory_out_en_T_5; // @[DataMemoryAccess.scala 44:71]
  wire [23:0] _io_memoryUnit_out_rdata_T_3 = io_dataMemory_in_rdata[31] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_memoryUnit_out_rdata_T_4 = {_io_memoryUnit_out_rdata_T_3,io_dataMemory_in_rdata[31:24]}; // @[Cat.scala 33:92]
  wire [23:0] _io_memoryUnit_out_rdata_T_8 = io_dataMemory_in_rdata[23] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_memoryUnit_out_rdata_T_9 = {_io_memoryUnit_out_rdata_T_8,io_dataMemory_in_rdata[23:16]}; // @[Cat.scala 33:92]
  wire [23:0] _io_memoryUnit_out_rdata_T_13 = io_dataMemory_in_rdata[15] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_memoryUnit_out_rdata_T_14 = {_io_memoryUnit_out_rdata_T_13,io_dataMemory_in_rdata[15:8]}; // @[Cat.scala 33:92]
  wire [23:0] _io_memoryUnit_out_rdata_T_18 = io_dataMemory_in_rdata[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_memoryUnit_out_rdata_T_19 = {_io_memoryUnit_out_rdata_T_18,io_dataMemory_in_rdata[7:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_21 = 2'h2 == mem_addr2 ? _io_memoryUnit_out_rdata_T_9 :
    _io_memoryUnit_out_rdata_T_4; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_23 = 2'h1 == mem_addr2 ? _io_memoryUnit_out_rdata_T_14 :
    _io_memoryUnit_out_rdata_T_21; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_25 = 2'h0 == mem_addr2 ? _io_memoryUnit_out_rdata_T_19 :
    _io_memoryUnit_out_rdata_T_23; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_28 = {24'h0,io_dataMemory_in_rdata[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_31 = {24'h0,io_dataMemory_in_rdata[23:16]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_34 = {24'h0,io_dataMemory_in_rdata[15:8]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_37 = {24'h0,io_dataMemory_in_rdata[7:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_39 = 2'h2 == mem_addr2 ? _io_memoryUnit_out_rdata_T_31 :
    _io_memoryUnit_out_rdata_T_28; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_41 = 2'h1 == mem_addr2 ? _io_memoryUnit_out_rdata_T_34 :
    _io_memoryUnit_out_rdata_T_39; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_43 = 2'h0 == mem_addr2 ? _io_memoryUnit_out_rdata_T_37 :
    _io_memoryUnit_out_rdata_T_41; // @[Mux.scala 81:58]
  wire [15:0] _io_memoryUnit_out_rdata_T_48 = io_dataMemory_in_rdata[31] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_memoryUnit_out_rdata_T_49 = {_io_memoryUnit_out_rdata_T_48,io_dataMemory_in_rdata[31:16]}; // @[Cat.scala 33:92]
  wire [15:0] _io_memoryUnit_out_rdata_T_53 = io_dataMemory_in_rdata[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_memoryUnit_out_rdata_T_54 = {_io_memoryUnit_out_rdata_T_53,io_dataMemory_in_rdata[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_55 = mem_addr2[1] ? _io_memoryUnit_out_rdata_T_49 :
    _io_memoryUnit_out_rdata_T_54; // @[DataMemoryAccess.scala 72:20]
  wire [31:0] _io_memoryUnit_out_rdata_T_59 = {16'h0,io_dataMemory_in_rdata[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_62 = {16'h0,io_dataMemory_in_rdata[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_63 = mem_addr2[1] ? _io_memoryUnit_out_rdata_T_59 :
    _io_memoryUnit_out_rdata_T_62; // @[DataMemoryAccess.scala 77:21]
  wire [31:0] _io_memoryUnit_out_rdata_T_66 = {io_dataMemory_in_rdata[23:0],io_memoryUnit_in_mem_wdata[7:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_69 = {io_dataMemory_in_rdata[15:0],io_memoryUnit_in_mem_wdata[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_72 = {io_dataMemory_in_rdata[7:0],io_memoryUnit_in_mem_wdata[23:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_74 = 2'h2 == mem_addr2 ? _io_memoryUnit_out_rdata_T_66 : io_dataMemory_in_rdata
    ; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_76 = 2'h1 == mem_addr2 ? _io_memoryUnit_out_rdata_T_69 :
    _io_memoryUnit_out_rdata_T_74; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_78 = 2'h0 == mem_addr2 ? _io_memoryUnit_out_rdata_T_72 :
    _io_memoryUnit_out_rdata_T_76; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_81 = {io_memoryUnit_in_mem_wdata[31:8],io_dataMemory_in_rdata[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_84 = {io_memoryUnit_in_mem_wdata[31:16],io_dataMemory_in_rdata[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_87 = {io_memoryUnit_in_mem_wdata[31:24],io_dataMemory_in_rdata[31:8]}; // @[Cat.scala 33:92]
  wire [31:0] _io_memoryUnit_out_rdata_T_89 = 2'h2 == mem_addr2 ? _io_memoryUnit_out_rdata_T_84 :
    _io_memoryUnit_out_rdata_T_81; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_91 = 2'h1 == mem_addr2 ? _io_memoryUnit_out_rdata_T_87 :
    _io_memoryUnit_out_rdata_T_89; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_93 = 2'h0 == mem_addr2 ? io_dataMemory_in_rdata : _io_memoryUnit_out_rdata_T_91
    ; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_95 = 7'h30 == io_memoryUnit_in_inst_info_op ? _io_memoryUnit_out_rdata_T_25 : 32'h0
    ; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_97 = 7'h31 == io_memoryUnit_in_inst_info_op ? _io_memoryUnit_out_rdata_T_43 :
    _io_memoryUnit_out_rdata_T_95; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_99 = 7'h32 == io_memoryUnit_in_inst_info_op ? _io_memoryUnit_out_rdata_T_55 :
    _io_memoryUnit_out_rdata_T_97; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_101 = 7'h33 == io_memoryUnit_in_inst_info_op ? _io_memoryUnit_out_rdata_T_63 :
    _io_memoryUnit_out_rdata_T_99; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_103 = 7'h35 == io_memoryUnit_in_inst_info_op ? io_dataMemory_in_rdata :
    _io_memoryUnit_out_rdata_T_101; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_105 = 7'h34 == io_memoryUnit_in_inst_info_op ? io_dataMemory_in_rdata :
    _io_memoryUnit_out_rdata_T_103; // @[Mux.scala 81:58]
  wire [31:0] _io_memoryUnit_out_rdata_T_107 = 7'h36 == io_memoryUnit_in_inst_info_op ? _io_memoryUnit_out_rdata_T_78 :
    _io_memoryUnit_out_rdata_T_105; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_2 = {io_memoryUnit_in_mem_wdata[7:0],io_memoryUnit_in_mem_wdata[7:0],
    io_memoryUnit_in_mem_wdata[7:0],io_memoryUnit_in_mem_wdata[7:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataMemory_out_wdata_T_4 = {io_memoryUnit_in_mem_wdata[15:0],io_memoryUnit_in_mem_wdata[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataMemory_out_wdata_T_6 = {8'h0,io_memoryUnit_in_mem_wdata[31:8]}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataMemory_out_wdata_T_8 = {16'h0,io_memoryUnit_in_mem_wdata[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataMemory_out_wdata_T_10 = {24'h0,io_memoryUnit_in_mem_wdata[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataMemory_out_wdata_T_12 = 2'h2 == mem_addr2 ? _io_dataMemory_out_wdata_T_6 :
    io_memoryUnit_in_mem_wdata; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_14 = 2'h1 == mem_addr2 ? _io_dataMemory_out_wdata_T_8 :
    _io_dataMemory_out_wdata_T_12; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_16 = 2'h0 == mem_addr2 ? _io_dataMemory_out_wdata_T_10 :
    _io_dataMemory_out_wdata_T_14; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_18 = {io_memoryUnit_in_mem_wdata[7:0],24'h0}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataMemory_out_wdata_T_20 = {io_memoryUnit_in_mem_wdata[15:0],16'h0}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataMemory_out_wdata_T_22 = {io_memoryUnit_in_mem_wdata[23:0],8'h0}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataMemory_out_wdata_T_24 = 2'h2 == mem_addr2 ? _io_dataMemory_out_wdata_T_20 :
    _io_dataMemory_out_wdata_T_18; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_26 = 2'h1 == mem_addr2 ? _io_dataMemory_out_wdata_T_22 :
    _io_dataMemory_out_wdata_T_24; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_28 = 2'h0 == mem_addr2 ? io_memoryUnit_in_mem_wdata :
    _io_dataMemory_out_wdata_T_26; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_30 = 7'h38 == io_memoryUnit_in_inst_info_op ? _io_dataMemory_out_wdata_T_2 :
    io_memoryUnit_in_mem_wdata; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_32 = 7'h3a == io_memoryUnit_in_inst_info_op ? _io_dataMemory_out_wdata_T_4 :
    _io_dataMemory_out_wdata_T_30; // @[Mux.scala 81:58]
  wire [31:0] _io_dataMemory_out_wdata_T_34 = 7'h3c == io_memoryUnit_in_inst_info_op ? _io_dataMemory_out_wdata_T_16 :
    _io_dataMemory_out_wdata_T_32; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_1 = 2'h2 == mem_addr2 ? 4'h4 : 4'h8; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_3 = 2'h1 == mem_addr2 ? 4'h2 : _io_dataMemory_out_wen_T_1; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_5 = 2'h0 == mem_addr2 ? 4'h1 : _io_dataMemory_out_wen_T_3; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_7 = mem_addr2[1] ? 4'hc : 4'h3; // @[DataMemoryAccess.scala 148:20]
  wire [3:0] _io_dataMemory_out_wen_T_9 = 2'h2 == mem_addr2 ? 4'h7 : 4'hf; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_11 = 2'h1 == mem_addr2 ? 4'h3 : _io_dataMemory_out_wen_T_9; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_13 = 2'h0 == mem_addr2 ? 4'h1 : _io_dataMemory_out_wen_T_11; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_15 = 2'h2 == mem_addr2 ? 4'hc : 4'h8; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_17 = 2'h1 == mem_addr2 ? 4'he : _io_dataMemory_out_wen_T_15; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_19 = 2'h0 == mem_addr2 ? 4'hf : _io_dataMemory_out_wen_T_17; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_21 = 7'h38 == io_memoryUnit_in_inst_info_op ? _io_dataMemory_out_wen_T_5 : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_23 = 7'h3a == io_memoryUnit_in_inst_info_op ? _io_dataMemory_out_wen_T_7 :
    _io_dataMemory_out_wen_T_21; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_25 = 7'h3b == io_memoryUnit_in_inst_info_op ? 4'hf : _io_dataMemory_out_wen_T_23; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_27 = 7'h39 == io_memoryUnit_in_inst_info_op ? 4'hf : _io_dataMemory_out_wen_T_25; // @[Mux.scala 81:58]
  wire [3:0] _io_dataMemory_out_wen_T_29 = 7'h3c == io_memoryUnit_in_inst_info_op ? _io_dataMemory_out_wen_T_13 :
    _io_dataMemory_out_wen_T_27; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_1 = 7'h35 == io_memoryUnit_in_inst_info_op ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_3 = 7'h34 == io_memoryUnit_in_inst_info_op ? 2'h2 : _io_dataMemory_out_rlen_T_1; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_5 = 7'h32 == io_memoryUnit_in_inst_info_op ? 2'h1 : _io_dataMemory_out_rlen_T_3; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_7 = 7'h33 == io_memoryUnit_in_inst_info_op ? 2'h1 : _io_dataMemory_out_rlen_T_5; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_9 = 7'h30 == io_memoryUnit_in_inst_info_op ? 2'h0 : _io_dataMemory_out_rlen_T_7; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_11 = 7'h31 == io_memoryUnit_in_inst_info_op ? 2'h0 : _io_dataMemory_out_rlen_T_9; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_13 = 7'h36 == io_memoryUnit_in_inst_info_op ? 2'h2 : _io_dataMemory_out_rlen_T_11
    ; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_15 = 7'h37 == io_memoryUnit_in_inst_info_op ? 2'h2 : _io_dataMemory_out_rlen_T_13
    ; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_17 = 7'h3b == io_memoryUnit_in_inst_info_op ? 2'h2 : _io_dataMemory_out_rlen_T_15
    ; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_19 = 7'h3c == io_memoryUnit_in_inst_info_op ? 2'h2 : _io_dataMemory_out_rlen_T_17
    ; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_21 = 7'h3d == io_memoryUnit_in_inst_info_op ? 2'h2 : _io_dataMemory_out_rlen_T_19
    ; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_23 = 7'h39 == io_memoryUnit_in_inst_info_op ? 2'h2 : _io_dataMemory_out_rlen_T_21
    ; // @[Mux.scala 81:58]
  wire [1:0] _io_dataMemory_out_rlen_T_25 = 7'h3a == io_memoryUnit_in_inst_info_op ? 2'h1 : _io_dataMemory_out_rlen_T_23
    ; // @[Mux.scala 81:58]
  assign io_memoryUnit_out_rdata = 7'h37 == io_memoryUnit_in_inst_info_op ? _io_memoryUnit_out_rdata_T_93 :
    _io_memoryUnit_out_rdata_T_107; // @[Mux.scala 81:58]
  assign io_dataMemory_out_en = io_memoryUnit_in_mem_en & _io_dataMemory_out_en_T_6; // @[DataMemoryAccess.scala 43:51]
  assign io_dataMemory_out_rlen = 7'h38 == io_memoryUnit_in_inst_info_op ? 2'h0 : _io_dataMemory_out_rlen_T_25; // @[Mux.scala 81:58]
  assign io_dataMemory_out_wen = 7'h3d == io_memoryUnit_in_inst_info_op ? _io_dataMemory_out_wen_T_19 :
    _io_dataMemory_out_wen_T_29; // @[Mux.scala 81:58]
  assign io_dataMemory_out_wdata = 7'h3d == io_memoryUnit_in_inst_info_op ? _io_dataMemory_out_wdata_T_28 :
    _io_dataMemory_out_wdata_T_34; // @[Mux.scala 81:58]
endmodule
module MemoryUnit(
  output        io_ctrl_flush_req,
  input         io_ctrl_allow_to_go,
  input  [31:0] io_memoryStage_inst0_pc,
  input  [3:0]  io_memoryStage_inst0_inst_info_fusel,
  input  [6:0]  io_memoryStage_inst0_inst_info_op,
  input         io_memoryStage_inst0_inst_info_reg_wen,
  input  [4:0]  io_memoryStage_inst0_inst_info_reg_waddr,
  input  [31:0] io_memoryStage_inst0_inst_info_inst,
  input  [31:0] io_memoryStage_inst0_rd_info_wdata,
  input         io_memoryStage_inst0_ex_flush_req,
  input         io_memoryStage_inst0_ex_eret,
  input  [31:0] io_memoryStage_inst0_ex_badvaddr,
  input         io_memoryStage_inst0_ex_bd,
  input  [4:0]  io_memoryStage_inst0_ex_excode,
  input  [31:0] io_memoryStage_inst0_cp0_cp0_count,
  input  [31:0] io_memoryStage_inst0_cp0_cp0_random,
  input  [31:0] io_memoryStage_inst0_cp0_cp0_cause,
  input         io_memoryStage_inst0_mem_en,
  input  [6:0]  io_memoryStage_inst0_mem_inst_info_op,
  input  [31:0] io_memoryStage_inst0_mem_addr,
  input  [31:0] io_memoryStage_inst0_mem_wdata,
  input         io_memoryStage_inst0_mem_sel_0,
  input         io_memoryStage_inst0_mem_sel_1,
  input  [31:0] io_memoryStage_inst1_pc,
  input  [3:0]  io_memoryStage_inst1_inst_info_fusel,
  input         io_memoryStage_inst1_inst_info_reg_wen,
  input  [4:0]  io_memoryStage_inst1_inst_info_reg_waddr,
  input  [31:0] io_memoryStage_inst1_rd_info_wdata,
  input         io_memoryStage_inst1_ex_flush_req,
  input         io_memoryStage_inst1_ex_eret,
  input  [31:0] io_memoryStage_inst1_ex_badvaddr,
  input         io_memoryStage_inst1_ex_bd,
  input  [4:0]  io_memoryStage_inst1_ex_excode,
  output        io_fetchUnit_flush,
  output [31:0] io_fetchUnit_flush_pc,
  output        io_fetchUnit_ex_flush,
  output [31:0] io_fetchUnit_ex_flush_pc,
  output        io_decoderUnit_0_wen,
  output [4:0]  io_decoderUnit_0_waddr,
  output [31:0] io_decoderUnit_0_wdata,
  output        io_decoderUnit_1_wen,
  output [4:0]  io_decoderUnit_1_waddr,
  output [31:0] io_decoderUnit_1_wdata,
  output [31:0] io_cp0_in_inst_0_pc,
  output        io_cp0_in_inst_0_ex_flush_req,
  output        io_cp0_in_inst_0_ex_tlb_refill,
  output        io_cp0_in_inst_0_ex_eret,
  output [31:0] io_cp0_in_inst_0_ex_badvaddr,
  output        io_cp0_in_inst_0_ex_bd,
  output [4:0]  io_cp0_in_inst_0_ex_excode,
  output [31:0] io_cp0_in_inst_1_pc,
  output        io_cp0_in_inst_1_ex_flush_req,
  output        io_cp0_in_inst_1_ex_tlb_refill,
  output        io_cp0_in_inst_1_ex_eret,
  output [31:0] io_cp0_in_inst_1_ex_badvaddr,
  output        io_cp0_in_inst_1_ex_bd,
  output [4:0]  io_cp0_in_inst_1_ex_excode,
  input         io_cp0_out_flush,
  input  [31:0] io_cp0_out_flush_pc,
  output [31:0] io_writeBackStage_inst0_pc,
  output [3:0]  io_writeBackStage_inst0_inst_info_fusel,
  output [6:0]  io_writeBackStage_inst0_inst_info_op,
  output        io_writeBackStage_inst0_inst_info_reg_wen,
  output [4:0]  io_writeBackStage_inst0_inst_info_reg_waddr,
  output [31:0] io_writeBackStage_inst0_inst_info_inst,
  output [31:0] io_writeBackStage_inst0_rd_info_wdata,
  output        io_writeBackStage_inst0_ex_flush_req,
  output        io_writeBackStage_inst0_ex_tlb_refill,
  output        io_writeBackStage_inst0_ex_eret,
  output [31:0] io_writeBackStage_inst0_ex_badvaddr,
  output        io_writeBackStage_inst0_ex_bd,
  output [4:0]  io_writeBackStage_inst0_ex_excode,
  output [31:0] io_writeBackStage_inst0_cp0_cp0_count,
  output [31:0] io_writeBackStage_inst0_cp0_cp0_random,
  output [31:0] io_writeBackStage_inst0_cp0_cp0_cause,
  output [31:0] io_writeBackStage_inst1_pc,
  output [3:0]  io_writeBackStage_inst1_inst_info_fusel,
  output        io_writeBackStage_inst1_inst_info_reg_wen,
  output [4:0]  io_writeBackStage_inst1_inst_info_reg_waddr,
  output [31:0] io_writeBackStage_inst1_rd_info_wdata,
  output        io_writeBackStage_inst1_ex_flush_req,
  output        io_writeBackStage_inst1_ex_tlb_refill,
  output        io_writeBackStage_inst1_ex_eret,
  output [31:0] io_writeBackStage_inst1_ex_badvaddr,
  output        io_writeBackStage_inst1_ex_bd,
  output [4:0]  io_writeBackStage_inst1_ex_excode,
  input         io_dataMemory_in_tlb_invalid,
  input         io_dataMemory_in_tlb_refill,
  input         io_dataMemory_in_tlb_modify,
  input  [31:0] io_dataMemory_in_rdata,
  output        io_dataMemory_out_en,
  output [1:0]  io_dataMemory_out_rlen,
  output [3:0]  io_dataMemory_out_wen,
  output [31:0] io_dataMemory_out_wdata
);
  wire  DataMemoryAccess_io_memoryUnit_in_mem_en; // @[MemoryUnit.scala 44:32]
  wire [6:0] DataMemoryAccess_io_memoryUnit_in_inst_info_op; // @[MemoryUnit.scala 44:32]
  wire [31:0] DataMemoryAccess_io_memoryUnit_in_mem_wdata; // @[MemoryUnit.scala 44:32]
  wire [31:0] DataMemoryAccess_io_memoryUnit_in_mem_addr; // @[MemoryUnit.scala 44:32]
  wire  DataMemoryAccess_io_memoryUnit_in_mem_sel_0; // @[MemoryUnit.scala 44:32]
  wire  DataMemoryAccess_io_memoryUnit_in_mem_sel_1; // @[MemoryUnit.scala 44:32]
  wire  DataMemoryAccess_io_memoryUnit_in_ex_0_flush_req; // @[MemoryUnit.scala 44:32]
  wire  DataMemoryAccess_io_memoryUnit_in_ex_1_flush_req; // @[MemoryUnit.scala 44:32]
  wire [31:0] DataMemoryAccess_io_memoryUnit_out_rdata; // @[MemoryUnit.scala 44:32]
  wire [31:0] DataMemoryAccess_io_dataMemory_in_rdata; // @[MemoryUnit.scala 44:32]
  wire  DataMemoryAccess_io_dataMemory_out_en; // @[MemoryUnit.scala 44:32]
  wire [1:0] DataMemoryAccess_io_dataMemory_out_rlen; // @[MemoryUnit.scala 44:32]
  wire [3:0] DataMemoryAccess_io_dataMemory_out_wen; // @[MemoryUnit.scala 44:32]
  wire [31:0] DataMemoryAccess_io_dataMemory_out_wdata; // @[MemoryUnit.scala 44:32]
  wire  _io_writeBackStage_inst0_rd_info_wdata_T_1 = io_writeBackStage_inst0_inst_info_fusel == 4'h4 &
    io_memoryStage_inst0_inst_info_reg_wen; // @[MemoryUnit.scala 65:56]
  wire  _inst0_access_mem_T_1 = io_dataMemory_out_en & (io_dataMemory_in_tlb_invalid | io_dataMemory_in_tlb_refill); // @[MemoryUnit.scala 71:27]
  wire  _inst0_access_mem_T_2 = io_memoryStage_inst0_inst_info_fusel == 4'h4; // @[MemoryUnit.scala 71:132]
  wire  inst0_access_mem = io_dataMemory_out_en & (io_dataMemory_in_tlb_invalid | io_dataMemory_in_tlb_refill) &
    io_memoryStage_inst0_inst_info_fusel == 4'h4; // @[MemoryUnit.scala 71:92]
  wire  _inst0_tlbmod_T = |io_dataMemory_out_wen; // @[MemoryUnit.scala 73:59]
  wire  _inst0_tlbmod_T_1 = io_dataMemory_in_tlb_modify & |io_dataMemory_out_wen; // @[MemoryUnit.scala 73:34]
  wire  inst0_tlbmod = io_dataMemory_in_tlb_modify & |io_dataMemory_out_wen & _inst0_access_mem_T_2; // @[MemoryUnit.scala 73:63]
  wire  _io_writeBackStage_inst0_ex_excode_T = io_memoryStage_inst0_ex_excode != 5'h0; // @[MemoryUnit.scala 77:39]
  wire [4:0] _io_writeBackStage_inst0_ex_excode_T_2 = _inst0_tlbmod_T ? 5'h4 : 5'h3; // @[MemoryUnit.scala 78:56]
  wire [4:0] _io_writeBackStage_inst0_ex_excode_T_3 = inst0_tlbmod ? 5'h2 : io_memoryStage_inst0_ex_excode; // @[Mux.scala 101:16]
  wire [4:0] _io_writeBackStage_inst0_ex_excode_T_4 = inst0_access_mem ? _io_writeBackStage_inst0_ex_excode_T_2 :
    _io_writeBackStage_inst0_ex_excode_T_3; // @[Mux.scala 101:16]
  wire  _io_writeBackStage_inst1_rd_info_wdata_T_1 = io_writeBackStage_inst1_inst_info_fusel == 4'h4 &
    io_memoryStage_inst1_inst_info_reg_wen; // @[MemoryUnit.scala 89:56]
  wire  _inst1_access_mem_T_2 = io_memoryStage_inst1_inst_info_fusel == 4'h4; // @[MemoryUnit.scala 95:132]
  wire  inst1_access_mem = _inst0_access_mem_T_1 & io_memoryStage_inst1_inst_info_fusel == 4'h4; // @[MemoryUnit.scala 95:92]
  wire  inst1_tlbmod = _inst0_tlbmod_T_1 & _inst1_access_mem_T_2; // @[MemoryUnit.scala 97:63]
  wire  _io_writeBackStage_inst1_ex_excode_T = io_memoryStage_inst1_ex_excode != 5'h0; // @[MemoryUnit.scala 101:39]
  wire [4:0] _io_writeBackStage_inst1_ex_excode_T_3 = inst1_tlbmod ? 5'h2 : io_memoryStage_inst1_ex_excode; // @[Mux.scala 101:16]
  wire [4:0] _io_writeBackStage_inst1_ex_excode_T_4 = inst1_access_mem ? _io_writeBackStage_inst0_ex_excode_T_2 :
    _io_writeBackStage_inst1_ex_excode_T_3; // @[Mux.scala 101:16]
  DataMemoryAccess DataMemoryAccess ( // @[MemoryUnit.scala 44:32]
    .io_memoryUnit_in_mem_en(DataMemoryAccess_io_memoryUnit_in_mem_en),
    .io_memoryUnit_in_inst_info_op(DataMemoryAccess_io_memoryUnit_in_inst_info_op),
    .io_memoryUnit_in_mem_wdata(DataMemoryAccess_io_memoryUnit_in_mem_wdata),
    .io_memoryUnit_in_mem_addr(DataMemoryAccess_io_memoryUnit_in_mem_addr),
    .io_memoryUnit_in_mem_sel_0(DataMemoryAccess_io_memoryUnit_in_mem_sel_0),
    .io_memoryUnit_in_mem_sel_1(DataMemoryAccess_io_memoryUnit_in_mem_sel_1),
    .io_memoryUnit_in_ex_0_flush_req(DataMemoryAccess_io_memoryUnit_in_ex_0_flush_req),
    .io_memoryUnit_in_ex_1_flush_req(DataMemoryAccess_io_memoryUnit_in_ex_1_flush_req),
    .io_memoryUnit_out_rdata(DataMemoryAccess_io_memoryUnit_out_rdata),
    .io_dataMemory_in_rdata(DataMemoryAccess_io_dataMemory_in_rdata),
    .io_dataMemory_out_en(DataMemoryAccess_io_dataMemory_out_en),
    .io_dataMemory_out_rlen(DataMemoryAccess_io_dataMemory_out_rlen),
    .io_dataMemory_out_wen(DataMemoryAccess_io_dataMemory_out_wen),
    .io_dataMemory_out_wdata(DataMemoryAccess_io_dataMemory_out_wdata)
  );
  assign io_ctrl_flush_req = io_fetchUnit_ex_flush | io_fetchUnit_flush; // @[MemoryUnit.scala 119:46]
  assign io_fetchUnit_flush = io_writeBackStage_inst0_inst_info_op == 7'h12 & io_ctrl_allow_to_go; // @[MemoryUnit.scala 114:81]
  assign io_fetchUnit_flush_pc = io_writeBackStage_inst0_pc + 32'h4; // @[MemoryUnit.scala 115:58]
  assign io_fetchUnit_ex_flush = io_cp0_out_flush; // @[MemoryUnit.scala 116:28]
  assign io_fetchUnit_ex_flush_pc = io_cp0_out_flush_pc; // @[MemoryUnit.scala 117:28]
  assign io_decoderUnit_0_wen = io_writeBackStage_inst0_inst_info_reg_wen; // @[MemoryUnit.scala 55:27]
  assign io_decoderUnit_0_waddr = io_writeBackStage_inst0_inst_info_reg_waddr; // @[MemoryUnit.scala 56:27]
  assign io_decoderUnit_0_wdata = io_writeBackStage_inst0_rd_info_wdata; // @[MemoryUnit.scala 57:27]
  assign io_decoderUnit_1_wen = io_writeBackStage_inst1_inst_info_reg_wen; // @[MemoryUnit.scala 58:27]
  assign io_decoderUnit_1_waddr = io_writeBackStage_inst1_inst_info_reg_waddr; // @[MemoryUnit.scala 59:27]
  assign io_decoderUnit_1_wdata = io_writeBackStage_inst1_rd_info_wdata; // @[MemoryUnit.scala 60:27]
  assign io_cp0_in_inst_0_pc = io_writeBackStage_inst0_pc; // @[MemoryUnit.scala 109:24]
  assign io_cp0_in_inst_0_ex_flush_req = io_writeBackStage_inst0_ex_flush_req; // @[MemoryUnit.scala 110:24]
  assign io_cp0_in_inst_0_ex_tlb_refill = io_writeBackStage_inst0_ex_tlb_refill; // @[MemoryUnit.scala 110:24]
  assign io_cp0_in_inst_0_ex_eret = io_writeBackStage_inst0_ex_eret; // @[MemoryUnit.scala 110:24]
  assign io_cp0_in_inst_0_ex_badvaddr = io_writeBackStage_inst0_ex_badvaddr; // @[MemoryUnit.scala 110:24]
  assign io_cp0_in_inst_0_ex_bd = io_writeBackStage_inst0_ex_bd; // @[MemoryUnit.scala 110:24]
  assign io_cp0_in_inst_0_ex_excode = io_writeBackStage_inst0_ex_excode; // @[MemoryUnit.scala 110:24]
  assign io_cp0_in_inst_1_pc = io_writeBackStage_inst1_pc; // @[MemoryUnit.scala 111:24]
  assign io_cp0_in_inst_1_ex_flush_req = io_writeBackStage_inst1_ex_flush_req; // @[MemoryUnit.scala 112:24]
  assign io_cp0_in_inst_1_ex_tlb_refill = io_writeBackStage_inst1_ex_tlb_refill; // @[MemoryUnit.scala 112:24]
  assign io_cp0_in_inst_1_ex_eret = io_writeBackStage_inst1_ex_eret; // @[MemoryUnit.scala 112:24]
  assign io_cp0_in_inst_1_ex_badvaddr = io_writeBackStage_inst1_ex_badvaddr; // @[MemoryUnit.scala 112:24]
  assign io_cp0_in_inst_1_ex_bd = io_writeBackStage_inst1_ex_bd; // @[MemoryUnit.scala 112:24]
  assign io_cp0_in_inst_1_ex_excode = io_writeBackStage_inst1_ex_excode; // @[MemoryUnit.scala 112:24]
  assign io_writeBackStage_inst0_pc = io_memoryStage_inst0_pc; // @[MemoryUnit.scala 62:37]
  assign io_writeBackStage_inst0_inst_info_fusel = io_memoryStage_inst0_inst_info_fusel; // @[MemoryUnit.scala 63:37]
  assign io_writeBackStage_inst0_inst_info_op = io_memoryStage_inst0_inst_info_op; // @[MemoryUnit.scala 63:37]
  assign io_writeBackStage_inst0_inst_info_reg_wen = io_memoryStage_inst0_inst_info_reg_wen; // @[MemoryUnit.scala 63:37]
  assign io_writeBackStage_inst0_inst_info_reg_waddr = io_memoryStage_inst0_inst_info_reg_waddr; // @[MemoryUnit.scala 63:37]
  assign io_writeBackStage_inst0_inst_info_inst = io_memoryStage_inst0_inst_info_inst; // @[MemoryUnit.scala 63:37]
  assign io_writeBackStage_inst0_rd_info_wdata = _io_writeBackStage_inst0_rd_info_wdata_T_1 ?
    DataMemoryAccess_io_memoryUnit_out_rdata : io_memoryStage_inst0_rd_info_wdata; // @[MemoryUnit.scala 64:47]
  assign io_writeBackStage_inst0_ex_flush_req = io_memoryStage_inst0_ex_flush_req | io_writeBackStage_inst0_ex_excode
     != 5'h0 | io_writeBackStage_inst0_ex_tlb_refill; // @[MemoryUnit.scala 83:124]
  assign io_writeBackStage_inst0_ex_tlb_refill = io_dataMemory_in_tlb_refill & _inst0_access_mem_T_2; // @[MemoryUnit.scala 82:72]
  assign io_writeBackStage_inst0_ex_eret = io_memoryStage_inst0_ex_eret; // @[MemoryUnit.scala 69:30]
  assign io_writeBackStage_inst0_ex_badvaddr = io_memoryStage_inst0_ex_badvaddr; // @[MemoryUnit.scala 69:30]
  assign io_writeBackStage_inst0_ex_bd = io_memoryStage_inst0_ex_bd; // @[MemoryUnit.scala 69:30]
  assign io_writeBackStage_inst0_ex_excode = _io_writeBackStage_inst0_ex_excode_T ? io_memoryStage_inst0_ex_excode :
    _io_writeBackStage_inst0_ex_excode_T_4; // @[Mux.scala 101:16]
  assign io_writeBackStage_inst0_cp0_cp0_count = io_memoryStage_inst0_cp0_cp0_count; // @[MemoryUnit.scala 84:31]
  assign io_writeBackStage_inst0_cp0_cp0_random = io_memoryStage_inst0_cp0_cp0_random; // @[MemoryUnit.scala 84:31]
  assign io_writeBackStage_inst0_cp0_cp0_cause = io_memoryStage_inst0_cp0_cp0_cause; // @[MemoryUnit.scala 84:31]
  assign io_writeBackStage_inst1_pc = io_memoryStage_inst1_pc; // @[MemoryUnit.scala 86:37]
  assign io_writeBackStage_inst1_inst_info_fusel = io_memoryStage_inst1_inst_info_fusel; // @[MemoryUnit.scala 87:37]
  assign io_writeBackStage_inst1_inst_info_reg_wen = io_memoryStage_inst1_inst_info_reg_wen; // @[MemoryUnit.scala 87:37]
  assign io_writeBackStage_inst1_inst_info_reg_waddr = io_memoryStage_inst1_inst_info_reg_waddr; // @[MemoryUnit.scala 87:37]
  assign io_writeBackStage_inst1_rd_info_wdata = _io_writeBackStage_inst1_rd_info_wdata_T_1 ?
    DataMemoryAccess_io_memoryUnit_out_rdata : io_memoryStage_inst1_rd_info_wdata; // @[MemoryUnit.scala 88:47]
  assign io_writeBackStage_inst1_ex_flush_req = io_memoryStage_inst1_ex_flush_req | io_writeBackStage_inst1_ex_excode
     != 5'h0 | io_writeBackStage_inst1_ex_tlb_refill; // @[MemoryUnit.scala 107:124]
  assign io_writeBackStage_inst1_ex_tlb_refill = io_dataMemory_in_tlb_refill & _inst1_access_mem_T_2; // @[MemoryUnit.scala 106:72]
  assign io_writeBackStage_inst1_ex_eret = io_memoryStage_inst1_ex_eret; // @[MemoryUnit.scala 93:30]
  assign io_writeBackStage_inst1_ex_badvaddr = io_memoryStage_inst1_ex_badvaddr; // @[MemoryUnit.scala 93:30]
  assign io_writeBackStage_inst1_ex_bd = io_memoryStage_inst1_ex_bd; // @[MemoryUnit.scala 93:30]
  assign io_writeBackStage_inst1_ex_excode = _io_writeBackStage_inst1_ex_excode_T ? io_memoryStage_inst1_ex_excode :
    _io_writeBackStage_inst1_ex_excode_T_4; // @[Mux.scala 101:16]
  assign io_dataMemory_out_en = DataMemoryAccess_io_dataMemory_out_en; // @[MemoryUnit.scala 53:44]
  assign io_dataMemory_out_rlen = DataMemoryAccess_io_dataMemory_out_rlen; // @[MemoryUnit.scala 53:44]
  assign io_dataMemory_out_wen = DataMemoryAccess_io_dataMemory_out_wen; // @[MemoryUnit.scala 53:44]
  assign io_dataMemory_out_wdata = DataMemoryAccess_io_dataMemory_out_wdata; // @[MemoryUnit.scala 53:44]
  assign DataMemoryAccess_io_memoryUnit_in_mem_en = io_memoryStage_inst0_mem_en; // @[MemoryUnit.scala 45:44]
  assign DataMemoryAccess_io_memoryUnit_in_inst_info_op = io_memoryStage_inst0_mem_inst_info_op; // @[MemoryUnit.scala 46:44]
  assign DataMemoryAccess_io_memoryUnit_in_mem_wdata = io_memoryStage_inst0_mem_wdata; // @[MemoryUnit.scala 47:44]
  assign DataMemoryAccess_io_memoryUnit_in_mem_addr = io_memoryStage_inst0_mem_addr; // @[MemoryUnit.scala 48:44]
  assign DataMemoryAccess_io_memoryUnit_in_mem_sel_0 = io_memoryStage_inst0_mem_sel_0; // @[MemoryUnit.scala 49:44]
  assign DataMemoryAccess_io_memoryUnit_in_mem_sel_1 = io_memoryStage_inst0_mem_sel_1; // @[MemoryUnit.scala 49:44]
  assign DataMemoryAccess_io_memoryUnit_in_ex_0_flush_req = io_memoryStage_inst0_ex_flush_req; // @[MemoryUnit.scala 50:44]
  assign DataMemoryAccess_io_memoryUnit_in_ex_1_flush_req = io_memoryStage_inst1_ex_flush_req; // @[MemoryUnit.scala 51:44]
  assign DataMemoryAccess_io_dataMemory_in_rdata = io_dataMemory_in_rdata; // @[MemoryUnit.scala 52:44]
endmodule
module WriteBackStage(
  input         clock,
  input         reset,
  input         io_ctrl_allow_to_go,
  input  [31:0] io_memoryUnit_inst0_pc,
  input         io_memoryUnit_inst0_inst_info_reg_wen,
  input  [4:0]  io_memoryUnit_inst0_inst_info_reg_waddr,
  input  [31:0] io_memoryUnit_inst0_rd_info_wdata,
  input         io_memoryUnit_inst0_ex_flush_req,
  input  [4:0]  io_memoryUnit_inst0_ex_excode,
  input  [31:0] io_memoryUnit_inst0_cp0_cp0_count,
  input  [31:0] io_memoryUnit_inst0_cp0_cp0_random,
  input  [31:0] io_memoryUnit_inst0_cp0_cp0_cause,
  input  [31:0] io_memoryUnit_inst1_pc,
  input         io_memoryUnit_inst1_inst_info_reg_wen,
  input  [4:0]  io_memoryUnit_inst1_inst_info_reg_waddr,
  input  [31:0] io_memoryUnit_inst1_rd_info_wdata,
  input         io_memoryUnit_inst1_ex_flush_req,
  output [31:0] io_writeBackUnit_inst0_pc,
  output        io_writeBackUnit_inst0_inst_info_reg_wen,
  output [4:0]  io_writeBackUnit_inst0_inst_info_reg_waddr,
  output [31:0] io_writeBackUnit_inst0_rd_info_wdata,
  output        io_writeBackUnit_inst0_ex_flush_req,
  output [4:0]  io_writeBackUnit_inst0_ex_excode,
  output [31:0] io_writeBackUnit_inst0_cp0_cp0_count,
  output [31:0] io_writeBackUnit_inst0_cp0_cp0_random,
  output [31:0] io_writeBackUnit_inst0_cp0_cp0_cause,
  output [31:0] io_writeBackUnit_inst1_pc,
  output        io_writeBackUnit_inst1_inst_info_reg_wen,
  output [4:0]  io_writeBackUnit_inst1_inst_info_reg_waddr,
  output [31:0] io_writeBackUnit_inst1_rd_info_wdata,
  output        io_writeBackUnit_inst1_ex_flush_req
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] inst0_pc; // @[WriteBackStage.scala 33:22]
  reg  inst0_inst_info_reg_wen; // @[WriteBackStage.scala 33:22]
  reg [4:0] inst0_inst_info_reg_waddr; // @[WriteBackStage.scala 33:22]
  reg [31:0] inst0_rd_info_wdata; // @[WriteBackStage.scala 33:22]
  reg  inst0_ex_flush_req; // @[WriteBackStage.scala 33:22]
  reg [4:0] inst0_ex_excode; // @[WriteBackStage.scala 33:22]
  reg [31:0] inst0_cp0_cp0_count; // @[WriteBackStage.scala 33:22]
  reg [31:0] inst0_cp0_cp0_random; // @[WriteBackStage.scala 33:22]
  reg [31:0] inst0_cp0_cp0_cause; // @[WriteBackStage.scala 33:22]
  reg [31:0] inst1_pc; // @[WriteBackStage.scala 34:22]
  reg  inst1_inst_info_reg_wen; // @[WriteBackStage.scala 34:22]
  reg [4:0] inst1_inst_info_reg_waddr; // @[WriteBackStage.scala 34:22]
  reg [31:0] inst1_rd_info_wdata; // @[WriteBackStage.scala 34:22]
  reg  inst1_ex_flush_req; // @[WriteBackStage.scala 34:22]
  assign io_writeBackUnit_inst0_pc = inst0_pc; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst0_inst_info_reg_wen = inst0_inst_info_reg_wen; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst0_inst_info_reg_waddr = inst0_inst_info_reg_waddr; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst0_rd_info_wdata = inst0_rd_info_wdata; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst0_ex_flush_req = inst0_ex_flush_req; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst0_ex_excode = inst0_ex_excode; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst0_cp0_cp0_count = inst0_cp0_cp0_count; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst0_cp0_cp0_random = inst0_cp0_cp0_random; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst0_cp0_cp0_cause = inst0_cp0_cp0_cause; // @[WriteBackStage.scala 48:26]
  assign io_writeBackUnit_inst1_pc = inst1_pc; // @[WriteBackStage.scala 49:26]
  assign io_writeBackUnit_inst1_inst_info_reg_wen = inst1_inst_info_reg_wen; // @[WriteBackStage.scala 49:26]
  assign io_writeBackUnit_inst1_inst_info_reg_waddr = inst1_inst_info_reg_waddr; // @[WriteBackStage.scala 49:26]
  assign io_writeBackUnit_inst1_rd_info_wdata = inst1_rd_info_wdata; // @[WriteBackStage.scala 49:26]
  assign io_writeBackUnit_inst1_ex_flush_req = inst1_ex_flush_req; // @[WriteBackStage.scala 49:26]
  always @(posedge clock) begin
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_pc <= 32'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_pc <= io_memoryUnit_inst0_pc; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_inst_info_reg_wen <= 1'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_inst_info_reg_wen <= io_memoryUnit_inst0_inst_info_reg_wen; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_inst_info_reg_waddr <= 5'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_inst_info_reg_waddr <= io_memoryUnit_inst0_inst_info_reg_waddr; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_rd_info_wdata <= 32'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_rd_info_wdata <= io_memoryUnit_inst0_rd_info_wdata; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_ex_flush_req <= 1'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_ex_flush_req <= io_memoryUnit_inst0_ex_flush_req; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_ex_excode <= 5'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_ex_excode <= io_memoryUnit_inst0_ex_excode; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_cp0_cp0_count <= 32'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_cp0_cp0_count <= io_memoryUnit_inst0_cp0_cp0_count; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_cp0_cp0_random <= 32'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_cp0_cp0_random <= io_memoryUnit_inst0_cp0_cp0_random; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 33:22]
      inst0_cp0_cp0_cause <= 32'h0; // @[WriteBackStage.scala 33:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 38:35]
      inst0_cp0_cp0_cause <= io_memoryUnit_inst0_cp0_cp0_cause; // @[WriteBackStage.scala 39:11]
    end
    if (reset) begin // @[WriteBackStage.scala 34:22]
      inst1_pc <= 32'h0; // @[WriteBackStage.scala 34:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 44:35]
      inst1_pc <= io_memoryUnit_inst1_pc; // @[WriteBackStage.scala 45:11]
    end
    if (reset) begin // @[WriteBackStage.scala 34:22]
      inst1_inst_info_reg_wen <= 1'h0; // @[WriteBackStage.scala 34:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 44:35]
      inst1_inst_info_reg_wen <= io_memoryUnit_inst1_inst_info_reg_wen; // @[WriteBackStage.scala 45:11]
    end
    if (reset) begin // @[WriteBackStage.scala 34:22]
      inst1_inst_info_reg_waddr <= 5'h0; // @[WriteBackStage.scala 34:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 44:35]
      inst1_inst_info_reg_waddr <= io_memoryUnit_inst1_inst_info_reg_waddr; // @[WriteBackStage.scala 45:11]
    end
    if (reset) begin // @[WriteBackStage.scala 34:22]
      inst1_rd_info_wdata <= 32'h0; // @[WriteBackStage.scala 34:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 44:35]
      inst1_rd_info_wdata <= io_memoryUnit_inst1_rd_info_wdata; // @[WriteBackStage.scala 45:11]
    end
    if (reset) begin // @[WriteBackStage.scala 34:22]
      inst1_ex_flush_req <= 1'h0; // @[WriteBackStage.scala 34:22]
    end else if (io_ctrl_allow_to_go) begin // @[WriteBackStage.scala 44:35]
      inst1_ex_flush_req <= io_memoryUnit_inst1_ex_flush_req; // @[WriteBackStage.scala 45:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst0_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  inst0_inst_info_reg_wen = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst0_inst_info_reg_waddr = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  inst0_rd_info_wdata = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  inst0_ex_flush_req = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  inst0_ex_excode = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  inst0_cp0_cp0_count = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  inst0_cp0_cp0_random = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  inst0_cp0_cp0_cause = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  inst1_pc = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  inst1_inst_info_reg_wen = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inst1_inst_info_reg_waddr = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  inst1_rd_info_wdata = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  inst1_ex_flush_req = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBackUnit(
  input         clock,
  input         reset,
  input         io_ctrl_allow_to_go,
  input  [31:0] io_writeBackStage_inst0_pc,
  input         io_writeBackStage_inst0_inst_info_reg_wen,
  input  [4:0]  io_writeBackStage_inst0_inst_info_reg_waddr,
  input  [31:0] io_writeBackStage_inst0_rd_info_wdata,
  input         io_writeBackStage_inst0_ex_flush_req,
  input  [4:0]  io_writeBackStage_inst0_ex_excode,
  input  [31:0] io_writeBackStage_inst0_cp0_cp0_count,
  input  [31:0] io_writeBackStage_inst0_cp0_cp0_random,
  input  [31:0] io_writeBackStage_inst0_cp0_cp0_cause,
  input  [31:0] io_writeBackStage_inst1_pc,
  input         io_writeBackStage_inst1_inst_info_reg_wen,
  input  [4:0]  io_writeBackStage_inst1_inst_info_reg_waddr,
  input  [31:0] io_writeBackStage_inst1_rd_info_wdata,
  input         io_writeBackStage_inst1_ex_flush_req,
  output        io_regfile_0_wen,
  output [4:0]  io_regfile_0_waddr,
  output [31:0] io_regfile_0_wdata,
  output        io_regfile_1_wen,
  output [4:0]  io_regfile_1_waddr,
  output [31:0] io_regfile_1_wdata,
  output [31:0] io_debug_wb_pc,
  output [3:0]  io_debug_wb_rf_wen,
  output [4:0]  io_debug_wb_rf_wnum,
  output [31:0] io_debug_wb_rf_wdata,
  output [31:0] io_debug_cp0_count,
  output [31:0] io_debug_cp0_random,
  output [31:0] io_debug_cp0_cause,
  output        io_debug_int,
  output        io_debug_commit
);
  wire  _io_regfile_0_wen_T_1 = ~io_writeBackStage_inst0_ex_flush_req; // @[WriteBackUnit.scala 19:73]
  wire [31:0] _io_debug_wb_pc_T_2 = io_writeBackStage_inst0_ex_flush_req ? 32'h0 : io_writeBackStage_inst1_pc; // @[WriteBackUnit.scala 31:8]
  wire [3:0] _io_debug_wb_rf_wen_T_4 = io_regfile_0_wen ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _io_debug_wb_rf_wen_T_6 = io_regfile_1_wen ? 4'hf : 4'h0; // @[Bitwise.scala 77:12]
  wire [3:0] _io_debug_wb_rf_wen_T_7 = clock ? _io_debug_wb_rf_wen_T_4 : _io_debug_wb_rf_wen_T_6; // @[WriteBackUnit.scala 36:8]
  assign io_regfile_0_wen = io_writeBackStage_inst0_inst_info_reg_wen & io_ctrl_allow_to_go & ~
    io_writeBackStage_inst0_ex_flush_req; // @[WriteBackUnit.scala 19:70]
  assign io_regfile_0_waddr = io_writeBackStage_inst0_inst_info_reg_waddr; // @[WriteBackUnit.scala 20:23]
  assign io_regfile_0_wdata = io_writeBackStage_inst0_rd_info_wdata; // @[WriteBackUnit.scala 21:23]
  assign io_regfile_1_wen = io_writeBackStage_inst1_inst_info_reg_wen & io_ctrl_allow_to_go & _io_regfile_0_wen_T_1 & ~
    io_writeBackStage_inst1_ex_flush_req; // @[WriteBackUnit.scala 24:111]
  assign io_regfile_1_waddr = io_writeBackStage_inst1_inst_info_reg_waddr; // @[WriteBackUnit.scala 25:23]
  assign io_regfile_1_wdata = io_writeBackStage_inst1_rd_info_wdata; // @[WriteBackUnit.scala 26:23]
  assign io_debug_wb_pc = clock ? io_writeBackStage_inst0_pc : _io_debug_wb_pc_T_2; // @[WriteBackUnit.scala 28:24]
  assign io_debug_wb_rf_wen = reset ? 4'h0 : _io_debug_wb_rf_wen_T_7; // @[WriteBackUnit.scala 33:28]
  assign io_debug_wb_rf_wnum = clock ? io_regfile_0_waddr : io_regfile_1_waddr; // @[WriteBackUnit.scala 42:29]
  assign io_debug_wb_rf_wdata = clock ? io_regfile_0_wdata : io_regfile_1_wdata; // @[WriteBackUnit.scala 47:30]
  assign io_debug_cp0_count = io_writeBackStage_inst0_cp0_cp0_count; // @[WriteBackUnit.scala 53:23]
  assign io_debug_cp0_random = io_writeBackStage_inst0_cp0_cp0_random; // @[WriteBackUnit.scala 54:23]
  assign io_debug_cp0_cause = io_writeBackStage_inst0_cp0_cp0_cause; // @[WriteBackUnit.scala 52:23]
  assign io_debug_int = io_writeBackStage_inst0_ex_excode == 5'h1; // @[WriteBackUnit.scala 55:60]
  assign io_debug_commit = io_ctrl_allow_to_go; // @[WriteBackUnit.scala 56:23]
endmodule
module Core(
  input         clock,
  input         reset,
  input  [5:0]  io_ext_int,
  output        io_inst_req,
  output [31:0] io_inst_addr_0,
  output [31:0] io_inst_addr_1,
  input  [31:0] io_inst_inst_0,
  input  [31:0] io_inst_inst_1,
  input         io_inst_inst_valid_0,
  input         io_inst_inst_valid_1,
  output        io_inst_cpu_stall,
  input         io_inst_icache_stall,
  input         io_inst_tlb1_invalid,
  input  [18:0] io_inst_tlb2_vpn,
  output        io_inst_tlb2_found,
  output [19:0] io_inst_tlb2_entry_pfn_0,
  output [19:0] io_inst_tlb2_entry_pfn_1,
  output        io_inst_tlb2_entry_c_0,
  output        io_inst_tlb2_entry_c_1,
  output        io_inst_tlb2_entry_v_0,
  output        io_inst_tlb2_entry_v_1,
  output        io_inst_fence_value,
  output [31:0] io_inst_fence_addr,
  output        io_inst_fence_tlb,
  output        io_data_stallM,
  input         io_data_dstall,
  output [31:0] io_data_E_mem_va,
  output [31:0] io_data_M_mem_va,
  output [31:0] io_data_M_fence_addr,
  output        io_data_M_fence_d,
  output        io_data_M_mem_en,
  output        io_data_M_mem_write,
  output [3:0]  io_data_M_wmask,
  output [1:0]  io_data_M_mem_size,
  output [31:0] io_data_M_wdata,
  input  [31:0] io_data_M_rdata,
  input  [18:0] io_data_tlb_vpn2,
  output        io_data_tlb_found,
  output [19:0] io_data_tlb_entry_pfn_0,
  output [19:0] io_data_tlb_entry_pfn_1,
  output        io_data_tlb_entry_c_0,
  output        io_data_tlb_entry_c_1,
  output        io_data_tlb_entry_d_0,
  output        io_data_tlb_entry_d_1,
  output        io_data_tlb_entry_v_0,
  output        io_data_tlb_entry_v_1,
  output        io_data_fence_tlb,
  input         io_data_data_tlb_refill,
  input         io_data_data_tlb_invalid,
  input         io_data_data_tlb_mod,
  output [31:0] io_debug_wb_pc,
  output [3:0]  io_debug_wb_rf_wen,
  output [4:0]  io_debug_wb_rf_wnum,
  output [31:0] io_debug_wb_rf_wdata,
  output [31:0] io_debug_cp0_count,
  output [31:0] io_debug_cp0_random,
  output [31:0] io_debug_cp0_cause,
  output        io_debug_int,
  output        io_debug_commit
);
  wire  Ctrl_io_cacheCtrl_iCache_stall; // @[Core.scala 24:30]
  wire  Ctrl_io_cacheCtrl_dCache_stall; // @[Core.scala 24:30]
  wire  Ctrl_io_fetchUnit_allow_to_go; // @[Core.scala 24:30]
  wire  Ctrl_io_instBuffer_delay_slot_do_flush; // @[Core.scala 24:30]
  wire  Ctrl_io_decoderUnit_inst0_src1_ren; // @[Core.scala 24:30]
  wire [4:0] Ctrl_io_decoderUnit_inst0_src1_raddr; // @[Core.scala 24:30]
  wire  Ctrl_io_decoderUnit_inst0_src2_ren; // @[Core.scala 24:30]
  wire [4:0] Ctrl_io_decoderUnit_inst0_src2_raddr; // @[Core.scala 24:30]
  wire  Ctrl_io_decoderUnit_branch_flag; // @[Core.scala 24:30]
  wire  Ctrl_io_decoderUnit_allow_to_go; // @[Core.scala 24:30]
  wire  Ctrl_io_decoderUnit_do_flush; // @[Core.scala 24:30]
  wire  Ctrl_io_executeUnit_inst_0_mem_ren; // @[Core.scala 24:30]
  wire [4:0] Ctrl_io_executeUnit_inst_0_reg_waddr; // @[Core.scala 24:30]
  wire  Ctrl_io_executeUnit_inst_1_mem_ren; // @[Core.scala 24:30]
  wire [4:0] Ctrl_io_executeUnit_inst_1_reg_waddr; // @[Core.scala 24:30]
  wire  Ctrl_io_executeUnit_fu_stall; // @[Core.scala 24:30]
  wire  Ctrl_io_executeUnit_branch_flag; // @[Core.scala 24:30]
  wire  Ctrl_io_executeUnit_allow_to_go; // @[Core.scala 24:30]
  wire  Ctrl_io_executeUnit_do_flush; // @[Core.scala 24:30]
  wire  Ctrl_io_executeUnit_fu_allow_to_go; // @[Core.scala 24:30]
  wire  Ctrl_io_executeUnit_fu_do_flush; // @[Core.scala 24:30]
  wire  Ctrl_io_memoryUnit_flush_req; // @[Core.scala 24:30]
  wire  Ctrl_io_memoryUnit_allow_to_go; // @[Core.scala 24:30]
  wire  Ctrl_io_memoryUnit_do_flush; // @[Core.scala 24:30]
  wire  Ctrl_io_writeBackUnit_allow_to_go; // @[Core.scala 24:30]
  wire  FetchStage_clock; // @[Core.scala 25:30]
  wire  FetchStage_reset; // @[Core.scala 25:30]
  wire  FetchStage_io_memory_ex; // @[Core.scala 25:30]
  wire [31:0] FetchStage_io_memory_ex_pc; // @[Core.scala 25:30]
  wire  FetchStage_io_memory_flush; // @[Core.scala 25:30]
  wire [31:0] FetchStage_io_memory_flush_pc; // @[Core.scala 25:30]
  wire  FetchStage_io_decoder_branch; // @[Core.scala 25:30]
  wire [31:0] FetchStage_io_decoder_target; // @[Core.scala 25:30]
  wire  FetchStage_io_execute_branch; // @[Core.scala 25:30]
  wire [31:0] FetchStage_io_execute_target; // @[Core.scala 25:30]
  wire  FetchStage_io_instBuffer_full; // @[Core.scala 25:30]
  wire  FetchStage_io_iCache_inst_valid_0; // @[Core.scala 25:30]
  wire  FetchStage_io_iCache_inst_valid_1; // @[Core.scala 25:30]
  wire [31:0] FetchStage_io_iCache_pc; // @[Core.scala 25:30]
  wire [31:0] FetchStage_io_iCache_pc_next; // @[Core.scala 25:30]
  wire  BPU_clock; // @[Core.scala 26:30]
  wire  BPU_reset; // @[Core.scala 26:30]
  wire [31:0] BPU_io_instrD; // @[Core.scala 26:30]
  wire  BPU_io_enaD; // @[Core.scala 26:30]
  wire [31:0] BPU_io_pcD; // @[Core.scala 26:30]
  wire [31:0] BPU_io_pc_plus4D; // @[Core.scala 26:30]
  wire [31:0] BPU_io_pcE; // @[Core.scala 26:30]
  wire  BPU_io_branchE; // @[Core.scala 26:30]
  wire  BPU_io_actual_takeE; // @[Core.scala 26:30]
  wire  BPU_io_branchD; // @[Core.scala 26:30]
  wire  BPU_io_pred_takeD; // @[Core.scala 26:30]
  wire [31:0] BPU_io_branch_targetD; // @[Core.scala 26:30]
  wire  InstBuffer_clock; // @[Core.scala 27:30]
  wire  InstBuffer_reset; // @[Core.scala 27:30]
  wire  InstBuffer_io_fifo_rst; // @[Core.scala 27:30]
  wire  InstBuffer_io_flush_delay_slot; // @[Core.scala 27:30]
  wire  InstBuffer_io_delay_sel_rst; // @[Core.scala 27:30]
  wire  InstBuffer_io_D_delay_rst; // @[Core.scala 27:30]
  wire  InstBuffer_io_E_delay_rst; // @[Core.scala 27:30]
  wire  InstBuffer_io_i_stall; // @[Core.scala 27:30]
  wire  InstBuffer_io_master_is_branch; // @[Core.scala 27:30]
  wire  InstBuffer_io_master_is_in_delayslot_o; // @[Core.scala 27:30]
  wire  InstBuffer_io_read_en_0; // @[Core.scala 27:30]
  wire  InstBuffer_io_read_en_1; // @[Core.scala 27:30]
  wire  InstBuffer_io_read_0_tlb_invalid; // @[Core.scala 27:30]
  wire [31:0] InstBuffer_io_read_0_data; // @[Core.scala 27:30]
  wire [31:0] InstBuffer_io_read_0_addr; // @[Core.scala 27:30]
  wire  InstBuffer_io_read_1_tlb_invalid; // @[Core.scala 27:30]
  wire [31:0] InstBuffer_io_read_1_data; // @[Core.scala 27:30]
  wire [31:0] InstBuffer_io_read_1_addr; // @[Core.scala 27:30]
  wire  InstBuffer_io_write_en_0; // @[Core.scala 27:30]
  wire  InstBuffer_io_write_en_1; // @[Core.scala 27:30]
  wire  InstBuffer_io_write_0_tlb_invalid; // @[Core.scala 27:30]
  wire [31:0] InstBuffer_io_write_0_data; // @[Core.scala 27:30]
  wire [31:0] InstBuffer_io_write_0_addr; // @[Core.scala 27:30]
  wire  InstBuffer_io_write_1_tlb_invalid; // @[Core.scala 27:30]
  wire [31:0] InstBuffer_io_write_1_data; // @[Core.scala 27:30]
  wire [31:0] InstBuffer_io_write_1_addr; // @[Core.scala 27:30]
  wire  InstBuffer_io_empty; // @[Core.scala 27:30]
  wire  InstBuffer_io_almost_empty; // @[Core.scala 27:30]
  wire  InstBuffer_io_full; // @[Core.scala 27:30]
  wire  DecoderUnit_io_instBuffer_inst_0_ready; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_instBuffer_inst_0_bits_pc; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_instBuffer_inst_0_bits_inst; // @[Core.scala 28:30]
  wire  DecoderUnit_io_instBuffer_inst_0_bits_tlb_invalid; // @[Core.scala 28:30]
  wire  DecoderUnit_io_instBuffer_inst_1_ready; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_instBuffer_inst_1_bits_pc; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_instBuffer_inst_1_bits_inst; // @[Core.scala 28:30]
  wire  DecoderUnit_io_instBuffer_inst_1_bits_tlb_invalid; // @[Core.scala 28:30]
  wire  DecoderUnit_io_instBuffer_info_inst0_is_in_delayslot; // @[Core.scala 28:30]
  wire  DecoderUnit_io_instBuffer_info_empty; // @[Core.scala 28:30]
  wire  DecoderUnit_io_instBuffer_info_almost_empty; // @[Core.scala 28:30]
  wire  DecoderUnit_io_instBuffer_inst0_is_jb; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_regfile_0_src1_raddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_regfile_0_src1_rdata; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_regfile_0_src2_raddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_regfile_0_src2_rdata; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_regfile_1_src1_raddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_regfile_1_src1_rdata; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_regfile_1_src2_raddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_regfile_1_src2_rdata; // @[Core.scala 28:30]
  wire  DecoderUnit_io_forward_0_exe_wen; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_forward_0_exe_waddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_forward_0_exe_wdata; // @[Core.scala 28:30]
  wire  DecoderUnit_io_forward_0_exe_mem_ren; // @[Core.scala 28:30]
  wire  DecoderUnit_io_forward_0_mem_wen; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_forward_0_mem_waddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_forward_0_mem_wdata; // @[Core.scala 28:30]
  wire  DecoderUnit_io_forward_1_exe_wen; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_forward_1_exe_waddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_forward_1_exe_wdata; // @[Core.scala 28:30]
  wire  DecoderUnit_io_forward_1_exe_mem_ren; // @[Core.scala 28:30]
  wire  DecoderUnit_io_forward_1_mem_wen; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_forward_1_mem_waddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_forward_1_mem_wdata; // @[Core.scala 28:30]
  wire  DecoderUnit_io_cp0_access_allowed; // @[Core.scala 28:30]
  wire  DecoderUnit_io_cp0_kernel_mode; // @[Core.scala 28:30]
  wire  DecoderUnit_io_cp0_intterupt_allowed; // @[Core.scala 28:30]
  wire [7:0] DecoderUnit_io_cp0_cause_ip; // @[Core.scala 28:30]
  wire [7:0] DecoderUnit_io_cp0_status_im; // @[Core.scala 28:30]
  wire  DecoderUnit_io_fetchUnit_branch; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_fetchUnit_target; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_bpu_pc; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_bpu_decoded_inst0_inst; // @[Core.scala 28:30]
  wire  DecoderUnit_io_bpu_inst_is_branch; // @[Core.scala 28:30]
  wire  DecoderUnit_io_bpu_pred_branch_flag; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_bpu_branch_target; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst0_pc; // @[Core.scala 28:30]
  wire [3:0] DecoderUnit_io_executeStage_inst0_inst_info_fusel; // @[Core.scala 28:30]
  wire [6:0] DecoderUnit_io_executeStage_inst0_inst_info_op; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst0_inst_info_reg_wen; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_executeStage_inst0_inst_info_reg_waddr; // @[Core.scala 28:30]
  wire [7:0] DecoderUnit_io_executeStage_inst0_inst_info_cp0_addr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst0_inst_info_inst; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst0_src_info_src1_data; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst0_src_info_src2_data; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst0_ex_flush_req; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst0_ex_tlb_refill; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst0_ex_eret; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst0_ex_badvaddr; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst0_ex_bd; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_executeStage_inst0_ex_excode; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst0_jb_info_jump_regiser_conflict; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst0_jb_info_is_branch; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst0_jb_info_pred_branch_flag; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst0_jb_info_branch_target; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst1_allow_to_go; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst1_pc; // @[Core.scala 28:30]
  wire [3:0] DecoderUnit_io_executeStage_inst1_inst_info_fusel; // @[Core.scala 28:30]
  wire [6:0] DecoderUnit_io_executeStage_inst1_inst_info_op; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst1_inst_info_reg_wen; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_executeStage_inst1_inst_info_reg_waddr; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst1_inst_info_inst; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst1_src_info_src1_data; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst1_src_info_src2_data; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst1_ex_flush_req; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst1_ex_tlb_refill; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst1_ex_eret; // @[Core.scala 28:30]
  wire [31:0] DecoderUnit_io_executeStage_inst1_ex_badvaddr; // @[Core.scala 28:30]
  wire  DecoderUnit_io_executeStage_inst1_ex_bd; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_executeStage_inst1_ex_excode; // @[Core.scala 28:30]
  wire  DecoderUnit_io_ctrl_inst0_src1_ren; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_ctrl_inst0_src1_raddr; // @[Core.scala 28:30]
  wire  DecoderUnit_io_ctrl_inst0_src2_ren; // @[Core.scala 28:30]
  wire [4:0] DecoderUnit_io_ctrl_inst0_src2_raddr; // @[Core.scala 28:30]
  wire  DecoderUnit_io_ctrl_branch_flag; // @[Core.scala 28:30]
  wire  DecoderUnit_io_ctrl_allow_to_go; // @[Core.scala 28:30]
  wire  ARegFile_clock; // @[Core.scala 29:30]
  wire  ARegFile_reset; // @[Core.scala 29:30]
  wire [4:0] ARegFile_io_read_0_src1_raddr; // @[Core.scala 29:30]
  wire [31:0] ARegFile_io_read_0_src1_rdata; // @[Core.scala 29:30]
  wire [4:0] ARegFile_io_read_0_src2_raddr; // @[Core.scala 29:30]
  wire [31:0] ARegFile_io_read_0_src2_rdata; // @[Core.scala 29:30]
  wire [4:0] ARegFile_io_read_1_src1_raddr; // @[Core.scala 29:30]
  wire [31:0] ARegFile_io_read_1_src1_rdata; // @[Core.scala 29:30]
  wire [4:0] ARegFile_io_read_1_src2_raddr; // @[Core.scala 29:30]
  wire [31:0] ARegFile_io_read_1_src2_rdata; // @[Core.scala 29:30]
  wire  ARegFile_io_write_0_wen; // @[Core.scala 29:30]
  wire [4:0] ARegFile_io_write_0_waddr; // @[Core.scala 29:30]
  wire [31:0] ARegFile_io_write_0_wdata; // @[Core.scala 29:30]
  wire  ARegFile_io_write_1_wen; // @[Core.scala 29:30]
  wire [4:0] ARegFile_io_write_1_waddr; // @[Core.scala 29:30]
  wire [31:0] ARegFile_io_write_1_wdata; // @[Core.scala 29:30]
  wire  ExecuteStage_clock; // @[Core.scala 30:30]
  wire  ExecuteStage_reset; // @[Core.scala 30:30]
  wire  ExecuteStage_io_ctrl_inst0_allow_to_go; // @[Core.scala 30:30]
  wire  ExecuteStage_io_ctrl_clear_0; // @[Core.scala 30:30]
  wire  ExecuteStage_io_ctrl_clear_1; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst0_pc; // @[Core.scala 30:30]
  wire [3:0] ExecuteStage_io_decoderUnit_inst0_inst_info_fusel; // @[Core.scala 30:30]
  wire [6:0] ExecuteStage_io_decoderUnit_inst0_inst_info_op; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst0_inst_info_reg_wen; // @[Core.scala 30:30]
  wire [4:0] ExecuteStage_io_decoderUnit_inst0_inst_info_reg_waddr; // @[Core.scala 30:30]
  wire [7:0] ExecuteStage_io_decoderUnit_inst0_inst_info_cp0_addr; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst0_inst_info_inst; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst0_src_info_src1_data; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst0_src_info_src2_data; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst0_ex_flush_req; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst0_ex_eret; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst0_ex_badvaddr; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst0_ex_bd; // @[Core.scala 30:30]
  wire [4:0] ExecuteStage_io_decoderUnit_inst0_ex_excode; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst0_jb_info_jump_regiser_conflict; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst0_jb_info_is_branch; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst0_jb_info_pred_branch_flag; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst0_jb_info_branch_target; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst1_allow_to_go; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst1_pc; // @[Core.scala 30:30]
  wire [3:0] ExecuteStage_io_decoderUnit_inst1_inst_info_fusel; // @[Core.scala 30:30]
  wire [6:0] ExecuteStage_io_decoderUnit_inst1_inst_info_op; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst1_inst_info_reg_wen; // @[Core.scala 30:30]
  wire [4:0] ExecuteStage_io_decoderUnit_inst1_inst_info_reg_waddr; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst1_inst_info_inst; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst1_src_info_src1_data; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst1_src_info_src2_data; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst1_ex_flush_req; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst1_ex_eret; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_decoderUnit_inst1_ex_badvaddr; // @[Core.scala 30:30]
  wire  ExecuteStage_io_decoderUnit_inst1_ex_bd; // @[Core.scala 30:30]
  wire [4:0] ExecuteStage_io_decoderUnit_inst1_ex_excode; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst0_pc; // @[Core.scala 30:30]
  wire [3:0] ExecuteStage_io_executeUnit_inst0_inst_info_fusel; // @[Core.scala 30:30]
  wire [6:0] ExecuteStage_io_executeUnit_inst0_inst_info_op; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst0_inst_info_reg_wen; // @[Core.scala 30:30]
  wire [4:0] ExecuteStage_io_executeUnit_inst0_inst_info_reg_waddr; // @[Core.scala 30:30]
  wire [7:0] ExecuteStage_io_executeUnit_inst0_inst_info_cp0_addr; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst0_inst_info_inst; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst0_src_info_src1_data; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst0_src_info_src2_data; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst0_ex_flush_req; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst0_ex_eret; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst0_ex_badvaddr; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst0_ex_bd; // @[Core.scala 30:30]
  wire [4:0] ExecuteStage_io_executeUnit_inst0_ex_excode; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst0_jb_info_jump_regiser_conflict; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst0_jb_info_is_branch; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst0_jb_info_pred_branch_flag; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst0_jb_info_branch_target; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst1_pc; // @[Core.scala 30:30]
  wire [3:0] ExecuteStage_io_executeUnit_inst1_inst_info_fusel; // @[Core.scala 30:30]
  wire [6:0] ExecuteStage_io_executeUnit_inst1_inst_info_op; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst1_inst_info_reg_wen; // @[Core.scala 30:30]
  wire [4:0] ExecuteStage_io_executeUnit_inst1_inst_info_reg_waddr; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst1_inst_info_inst; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst1_src_info_src1_data; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst1_src_info_src2_data; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst1_ex_flush_req; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst1_ex_eret; // @[Core.scala 30:30]
  wire [31:0] ExecuteStage_io_executeUnit_inst1_ex_badvaddr; // @[Core.scala 30:30]
  wire  ExecuteStage_io_executeUnit_inst1_ex_bd; // @[Core.scala 30:30]
  wire [4:0] ExecuteStage_io_executeUnit_inst1_ex_excode; // @[Core.scala 30:30]
  wire  ExecuteUnit_clock; // @[Core.scala 31:30]
  wire  ExecuteUnit_reset; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_ctrl_inst_0_mem_ren; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_ctrl_inst_0_reg_waddr; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_ctrl_inst_1_mem_ren; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_ctrl_inst_1_reg_waddr; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_ctrl_fu_stall; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_ctrl_branch_flag; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_ctrl_allow_to_go; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_ctrl_fu_allow_to_go; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_ctrl_fu_do_flush; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst0_pc; // @[Core.scala 31:30]
  wire [3:0] ExecuteUnit_io_executeStage_inst0_inst_info_fusel; // @[Core.scala 31:30]
  wire [6:0] ExecuteUnit_io_executeStage_inst0_inst_info_op; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst0_inst_info_reg_wen; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_executeStage_inst0_inst_info_reg_waddr; // @[Core.scala 31:30]
  wire [7:0] ExecuteUnit_io_executeStage_inst0_inst_info_cp0_addr; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst0_inst_info_inst; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst0_src_info_src1_data; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst0_src_info_src2_data; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst0_ex_flush_req; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst0_ex_eret; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst0_ex_badvaddr; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst0_ex_bd; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_executeStage_inst0_ex_excode; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst0_jb_info_jump_regiser_conflict; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst0_jb_info_is_branch; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst0_jb_info_pred_branch_flag; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst0_jb_info_branch_target; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst1_pc; // @[Core.scala 31:30]
  wire [3:0] ExecuteUnit_io_executeStage_inst1_inst_info_fusel; // @[Core.scala 31:30]
  wire [6:0] ExecuteUnit_io_executeStage_inst1_inst_info_op; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst1_inst_info_reg_wen; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_executeStage_inst1_inst_info_reg_waddr; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst1_inst_info_inst; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst1_src_info_src1_data; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst1_src_info_src2_data; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst1_ex_flush_req; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst1_ex_eret; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_executeStage_inst1_ex_badvaddr; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_executeStage_inst1_ex_bd; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_executeStage_inst1_ex_excode; // @[Core.scala 31:30]
  wire [6:0] ExecuteUnit_io_cp0_in_inst_info_op; // @[Core.scala 31:30]
  wire [7:0] ExecuteUnit_io_cp0_in_inst_info_cp0_addr; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_cp0_in_mtc0_wdata; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_cp0_out_cp0_rdata; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_cp0_out_debug_cp0_count; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_cp0_out_debug_cp0_random; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_cp0_out_debug_cp0_cause; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_bpu_pc; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_bpu_branch_flag; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_bpu_inst0_is_branch; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_fetchStage_branch; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_fetchStage_target; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_decoderUnit_forward_0_exe_wen; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_decoderUnit_forward_0_exe_waddr; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_decoderUnit_forward_0_exe_wdata; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_decoderUnit_forward_0_exe_mem_ren; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_decoderUnit_forward_1_exe_wen; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_decoderUnit_forward_1_exe_waddr; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_decoderUnit_forward_1_exe_wdata; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_decoderUnit_forward_1_exe_mem_ren; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_decoderUnit_inst0_bd; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_pc; // @[Core.scala 31:30]
  wire [3:0] ExecuteUnit_io_memoryStage_inst0_inst_info_fusel; // @[Core.scala 31:30]
  wire [6:0] ExecuteUnit_io_memoryStage_inst0_inst_info_op; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst0_inst_info_reg_wen; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_memoryStage_inst0_inst_info_reg_waddr; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_inst_info_inst; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_rd_info_wdata; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst0_ex_flush_req; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst0_ex_eret; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_ex_badvaddr; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst0_ex_bd; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_memoryStage_inst0_ex_excode; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_cp0_cp0_count; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_cp0_cp0_random; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_cp0_cp0_cause; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst0_mem_en; // @[Core.scala 31:30]
  wire [6:0] ExecuteUnit_io_memoryStage_inst0_mem_inst_info_op; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_mem_addr; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst0_mem_wdata; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst0_mem_sel_0; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst0_mem_sel_1; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst1_pc; // @[Core.scala 31:30]
  wire [3:0] ExecuteUnit_io_memoryStage_inst1_inst_info_fusel; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst1_inst_info_reg_wen; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_memoryStage_inst1_inst_info_reg_waddr; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst1_rd_info_wdata; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst1_ex_flush_req; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst1_ex_eret; // @[Core.scala 31:30]
  wire [31:0] ExecuteUnit_io_memoryStage_inst1_ex_badvaddr; // @[Core.scala 31:30]
  wire  ExecuteUnit_io_memoryStage_inst1_ex_bd; // @[Core.scala 31:30]
  wire [4:0] ExecuteUnit_io_memoryStage_inst1_ex_excode; // @[Core.scala 31:30]
  wire  Cp0_clock; // @[Core.scala 32:30]
  wire  Cp0_reset; // @[Core.scala 32:30]
  wire [5:0] Cp0_io_ext_int; // @[Core.scala 32:30]
  wire  Cp0_io_ctrl_exe_stall; // @[Core.scala 32:30]
  wire  Cp0_io_ctrl_mem_stall; // @[Core.scala 32:30]
  wire  Cp0_io_decoderUnit_access_allowed; // @[Core.scala 32:30]
  wire  Cp0_io_decoderUnit_kernel_mode; // @[Core.scala 32:30]
  wire  Cp0_io_decoderUnit_intterupt_allowed; // @[Core.scala 32:30]
  wire [7:0] Cp0_io_decoderUnit_cause_ip; // @[Core.scala 32:30]
  wire [7:0] Cp0_io_decoderUnit_status_im; // @[Core.scala 32:30]
  wire [6:0] Cp0_io_executeUnit_in_inst_info_op; // @[Core.scala 32:30]
  wire [7:0] Cp0_io_executeUnit_in_inst_info_cp0_addr; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_executeUnit_in_mtc0_wdata; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_executeUnit_out_cp0_rdata; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_executeUnit_out_debug_cp0_count; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_executeUnit_out_debug_cp0_random; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_executeUnit_out_debug_cp0_cause; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_memoryUnit_in_inst_0_pc; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_in_inst_0_ex_flush_req; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_in_inst_0_ex_tlb_refill; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_in_inst_0_ex_eret; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_memoryUnit_in_inst_0_ex_badvaddr; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_in_inst_0_ex_bd; // @[Core.scala 32:30]
  wire [4:0] Cp0_io_memoryUnit_in_inst_0_ex_excode; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_memoryUnit_in_inst_1_pc; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_in_inst_1_ex_flush_req; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_in_inst_1_ex_tlb_refill; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_in_inst_1_ex_eret; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_memoryUnit_in_inst_1_ex_badvaddr; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_in_inst_1_ex_bd; // @[Core.scala 32:30]
  wire [4:0] Cp0_io_memoryUnit_in_inst_1_ex_excode; // @[Core.scala 32:30]
  wire  Cp0_io_memoryUnit_out_flush; // @[Core.scala 32:30]
  wire [31:0] Cp0_io_memoryUnit_out_flush_pc; // @[Core.scala 32:30]
  wire [18:0] Cp0_io_tlb_0_vpn2; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_0_found; // @[Core.scala 32:30]
  wire [19:0] Cp0_io_tlb_0_info_pfn_0; // @[Core.scala 32:30]
  wire [19:0] Cp0_io_tlb_0_info_pfn_1; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_0_info_c_0; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_0_info_c_1; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_0_info_v_0; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_0_info_v_1; // @[Core.scala 32:30]
  wire [18:0] Cp0_io_tlb_1_vpn2; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_1_found; // @[Core.scala 32:30]
  wire [19:0] Cp0_io_tlb_1_info_pfn_0; // @[Core.scala 32:30]
  wire [19:0] Cp0_io_tlb_1_info_pfn_1; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_1_info_c_0; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_1_info_c_1; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_1_info_d_0; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_1_info_d_1; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_1_info_v_0; // @[Core.scala 32:30]
  wire  Cp0_io_tlb_1_info_v_1; // @[Core.scala 32:30]
  wire  MemoryStage_clock; // @[Core.scala 33:30]
  wire  MemoryStage_reset; // @[Core.scala 33:30]
  wire  MemoryStage_io_ctrl_allow_to_go; // @[Core.scala 33:30]
  wire  MemoryStage_io_ctrl_clear_0; // @[Core.scala 33:30]
  wire  MemoryStage_io_ctrl_clear_1; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_pc; // @[Core.scala 33:30]
  wire [3:0] MemoryStage_io_executeUnit_inst0_inst_info_fusel; // @[Core.scala 33:30]
  wire [6:0] MemoryStage_io_executeUnit_inst0_inst_info_op; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst0_inst_info_reg_wen; // @[Core.scala 33:30]
  wire [4:0] MemoryStage_io_executeUnit_inst0_inst_info_reg_waddr; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_inst_info_inst; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_rd_info_wdata; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst0_ex_flush_req; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst0_ex_eret; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_ex_badvaddr; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst0_ex_bd; // @[Core.scala 33:30]
  wire [4:0] MemoryStage_io_executeUnit_inst0_ex_excode; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_cp0_cp0_count; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_cp0_cp0_random; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_cp0_cp0_cause; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst0_mem_en; // @[Core.scala 33:30]
  wire [6:0] MemoryStage_io_executeUnit_inst0_mem_inst_info_op; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_mem_addr; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst0_mem_wdata; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst0_mem_sel_0; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst0_mem_sel_1; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst1_pc; // @[Core.scala 33:30]
  wire [3:0] MemoryStage_io_executeUnit_inst1_inst_info_fusel; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst1_inst_info_reg_wen; // @[Core.scala 33:30]
  wire [4:0] MemoryStage_io_executeUnit_inst1_inst_info_reg_waddr; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst1_rd_info_wdata; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst1_ex_flush_req; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst1_ex_eret; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_executeUnit_inst1_ex_badvaddr; // @[Core.scala 33:30]
  wire  MemoryStage_io_executeUnit_inst1_ex_bd; // @[Core.scala 33:30]
  wire [4:0] MemoryStage_io_executeUnit_inst1_ex_excode; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_pc; // @[Core.scala 33:30]
  wire [3:0] MemoryStage_io_memoryUnit_inst0_inst_info_fusel; // @[Core.scala 33:30]
  wire [6:0] MemoryStage_io_memoryUnit_inst0_inst_info_op; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst0_inst_info_reg_wen; // @[Core.scala 33:30]
  wire [4:0] MemoryStage_io_memoryUnit_inst0_inst_info_reg_waddr; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_inst_info_inst; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_rd_info_wdata; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst0_ex_flush_req; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst0_ex_eret; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_ex_badvaddr; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst0_ex_bd; // @[Core.scala 33:30]
  wire [4:0] MemoryStage_io_memoryUnit_inst0_ex_excode; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_cp0_cp0_count; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_cp0_cp0_random; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_cp0_cp0_cause; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst0_mem_en; // @[Core.scala 33:30]
  wire [6:0] MemoryStage_io_memoryUnit_inst0_mem_inst_info_op; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_mem_addr; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst0_mem_wdata; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst0_mem_sel_0; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst0_mem_sel_1; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst1_pc; // @[Core.scala 33:30]
  wire [3:0] MemoryStage_io_memoryUnit_inst1_inst_info_fusel; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst1_inst_info_reg_wen; // @[Core.scala 33:30]
  wire [4:0] MemoryStage_io_memoryUnit_inst1_inst_info_reg_waddr; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst1_rd_info_wdata; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst1_ex_flush_req; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst1_ex_eret; // @[Core.scala 33:30]
  wire [31:0] MemoryStage_io_memoryUnit_inst1_ex_badvaddr; // @[Core.scala 33:30]
  wire  MemoryStage_io_memoryUnit_inst1_ex_bd; // @[Core.scala 33:30]
  wire [4:0] MemoryStage_io_memoryUnit_inst1_ex_excode; // @[Core.scala 33:30]
  wire  MemoryUnit_io_ctrl_flush_req; // @[Core.scala 34:30]
  wire  MemoryUnit_io_ctrl_allow_to_go; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_pc; // @[Core.scala 34:30]
  wire [3:0] MemoryUnit_io_memoryStage_inst0_inst_info_fusel; // @[Core.scala 34:30]
  wire [6:0] MemoryUnit_io_memoryStage_inst0_inst_info_op; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst0_inst_info_reg_wen; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_memoryStage_inst0_inst_info_reg_waddr; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_inst_info_inst; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_rd_info_wdata; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst0_ex_flush_req; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst0_ex_eret; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_ex_badvaddr; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst0_ex_bd; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_memoryStage_inst0_ex_excode; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_cp0_cp0_count; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_cp0_cp0_random; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_cp0_cp0_cause; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst0_mem_en; // @[Core.scala 34:30]
  wire [6:0] MemoryUnit_io_memoryStage_inst0_mem_inst_info_op; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_mem_addr; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst0_mem_wdata; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst0_mem_sel_0; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst0_mem_sel_1; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst1_pc; // @[Core.scala 34:30]
  wire [3:0] MemoryUnit_io_memoryStage_inst1_inst_info_fusel; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst1_inst_info_reg_wen; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_memoryStage_inst1_inst_info_reg_waddr; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst1_rd_info_wdata; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst1_ex_flush_req; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst1_ex_eret; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_memoryStage_inst1_ex_badvaddr; // @[Core.scala 34:30]
  wire  MemoryUnit_io_memoryStage_inst1_ex_bd; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_memoryStage_inst1_ex_excode; // @[Core.scala 34:30]
  wire  MemoryUnit_io_fetchUnit_flush; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_fetchUnit_flush_pc; // @[Core.scala 34:30]
  wire  MemoryUnit_io_fetchUnit_ex_flush; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_fetchUnit_ex_flush_pc; // @[Core.scala 34:30]
  wire  MemoryUnit_io_decoderUnit_0_wen; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_decoderUnit_0_waddr; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_decoderUnit_0_wdata; // @[Core.scala 34:30]
  wire  MemoryUnit_io_decoderUnit_1_wen; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_decoderUnit_1_waddr; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_decoderUnit_1_wdata; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_cp0_in_inst_0_pc; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_in_inst_0_ex_flush_req; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_in_inst_0_ex_tlb_refill; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_in_inst_0_ex_eret; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_cp0_in_inst_0_ex_badvaddr; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_in_inst_0_ex_bd; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_cp0_in_inst_0_ex_excode; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_cp0_in_inst_1_pc; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_in_inst_1_ex_flush_req; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_in_inst_1_ex_tlb_refill; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_in_inst_1_ex_eret; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_cp0_in_inst_1_ex_badvaddr; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_in_inst_1_ex_bd; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_cp0_in_inst_1_ex_excode; // @[Core.scala 34:30]
  wire  MemoryUnit_io_cp0_out_flush; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_cp0_out_flush_pc; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst0_pc; // @[Core.scala 34:30]
  wire [3:0] MemoryUnit_io_writeBackStage_inst0_inst_info_fusel; // @[Core.scala 34:30]
  wire [6:0] MemoryUnit_io_writeBackStage_inst0_inst_info_op; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst0_inst_info_reg_wen; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_writeBackStage_inst0_inst_info_reg_waddr; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst0_inst_info_inst; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst0_rd_info_wdata; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst0_ex_flush_req; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst0_ex_tlb_refill; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst0_ex_eret; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst0_ex_badvaddr; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst0_ex_bd; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_writeBackStage_inst0_ex_excode; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst0_cp0_cp0_count; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst0_cp0_cp0_random; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst0_cp0_cp0_cause; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst1_pc; // @[Core.scala 34:30]
  wire [3:0] MemoryUnit_io_writeBackStage_inst1_inst_info_fusel; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst1_inst_info_reg_wen; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_writeBackStage_inst1_inst_info_reg_waddr; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst1_rd_info_wdata; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst1_ex_flush_req; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst1_ex_tlb_refill; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst1_ex_eret; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_writeBackStage_inst1_ex_badvaddr; // @[Core.scala 34:30]
  wire  MemoryUnit_io_writeBackStage_inst1_ex_bd; // @[Core.scala 34:30]
  wire [4:0] MemoryUnit_io_writeBackStage_inst1_ex_excode; // @[Core.scala 34:30]
  wire  MemoryUnit_io_dataMemory_in_tlb_invalid; // @[Core.scala 34:30]
  wire  MemoryUnit_io_dataMemory_in_tlb_refill; // @[Core.scala 34:30]
  wire  MemoryUnit_io_dataMemory_in_tlb_modify; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_dataMemory_in_rdata; // @[Core.scala 34:30]
  wire  MemoryUnit_io_dataMemory_out_en; // @[Core.scala 34:30]
  wire [1:0] MemoryUnit_io_dataMemory_out_rlen; // @[Core.scala 34:30]
  wire [3:0] MemoryUnit_io_dataMemory_out_wen; // @[Core.scala 34:30]
  wire [31:0] MemoryUnit_io_dataMemory_out_wdata; // @[Core.scala 34:30]
  wire  WriteBackStage_clock; // @[Core.scala 35:30]
  wire  WriteBackStage_reset; // @[Core.scala 35:30]
  wire  WriteBackStage_io_ctrl_allow_to_go; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_memoryUnit_inst0_pc; // @[Core.scala 35:30]
  wire  WriteBackStage_io_memoryUnit_inst0_inst_info_reg_wen; // @[Core.scala 35:30]
  wire [4:0] WriteBackStage_io_memoryUnit_inst0_inst_info_reg_waddr; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_memoryUnit_inst0_rd_info_wdata; // @[Core.scala 35:30]
  wire  WriteBackStage_io_memoryUnit_inst0_ex_flush_req; // @[Core.scala 35:30]
  wire [4:0] WriteBackStage_io_memoryUnit_inst0_ex_excode; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_memoryUnit_inst0_cp0_cp0_count; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_memoryUnit_inst0_cp0_cp0_random; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_memoryUnit_inst0_cp0_cp0_cause; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_memoryUnit_inst1_pc; // @[Core.scala 35:30]
  wire  WriteBackStage_io_memoryUnit_inst1_inst_info_reg_wen; // @[Core.scala 35:30]
  wire [4:0] WriteBackStage_io_memoryUnit_inst1_inst_info_reg_waddr; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_memoryUnit_inst1_rd_info_wdata; // @[Core.scala 35:30]
  wire  WriteBackStage_io_memoryUnit_inst1_ex_flush_req; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_writeBackUnit_inst0_pc; // @[Core.scala 35:30]
  wire  WriteBackStage_io_writeBackUnit_inst0_inst_info_reg_wen; // @[Core.scala 35:30]
  wire [4:0] WriteBackStage_io_writeBackUnit_inst0_inst_info_reg_waddr; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_writeBackUnit_inst0_rd_info_wdata; // @[Core.scala 35:30]
  wire  WriteBackStage_io_writeBackUnit_inst0_ex_flush_req; // @[Core.scala 35:30]
  wire [4:0] WriteBackStage_io_writeBackUnit_inst0_ex_excode; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_count; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_random; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_cause; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_writeBackUnit_inst1_pc; // @[Core.scala 35:30]
  wire  WriteBackStage_io_writeBackUnit_inst1_inst_info_reg_wen; // @[Core.scala 35:30]
  wire [4:0] WriteBackStage_io_writeBackUnit_inst1_inst_info_reg_waddr; // @[Core.scala 35:30]
  wire [31:0] WriteBackStage_io_writeBackUnit_inst1_rd_info_wdata; // @[Core.scala 35:30]
  wire  WriteBackStage_io_writeBackUnit_inst1_ex_flush_req; // @[Core.scala 35:30]
  wire  WriteBackUnit_clock; // @[Core.scala 36:30]
  wire  WriteBackUnit_reset; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_ctrl_allow_to_go; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_writeBackStage_inst0_pc; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_writeBackStage_inst0_inst_info_reg_wen; // @[Core.scala 36:30]
  wire [4:0] WriteBackUnit_io_writeBackStage_inst0_inst_info_reg_waddr; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_writeBackStage_inst0_rd_info_wdata; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_writeBackStage_inst0_ex_flush_req; // @[Core.scala 36:30]
  wire [4:0] WriteBackUnit_io_writeBackStage_inst0_ex_excode; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_count; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_random; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_cause; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_writeBackStage_inst1_pc; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_writeBackStage_inst1_inst_info_reg_wen; // @[Core.scala 36:30]
  wire [4:0] WriteBackUnit_io_writeBackStage_inst1_inst_info_reg_waddr; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_writeBackStage_inst1_rd_info_wdata; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_writeBackStage_inst1_ex_flush_req; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_regfile_0_wen; // @[Core.scala 36:30]
  wire [4:0] WriteBackUnit_io_regfile_0_waddr; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_regfile_0_wdata; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_regfile_1_wen; // @[Core.scala 36:30]
  wire [4:0] WriteBackUnit_io_regfile_1_waddr; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_regfile_1_wdata; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_debug_wb_pc; // @[Core.scala 36:30]
  wire [3:0] WriteBackUnit_io_debug_wb_rf_wen; // @[Core.scala 36:30]
  wire [4:0] WriteBackUnit_io_debug_wb_rf_wnum; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_debug_wb_rf_wdata; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_debug_cp0_count; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_debug_cp0_random; // @[Core.scala 36:30]
  wire [31:0] WriteBackUnit_io_debug_cp0_cause; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_debug_int; // @[Core.scala 36:30]
  wire  WriteBackUnit_io_debug_commit; // @[Core.scala 36:30]
  wire  _T_5 = ~(ExecuteUnit_io_memoryStage_inst1_ex_bd | DecoderUnit_io_executeStage_inst0_ex_bd); // @[Core.scala 74:5]
  wire  _T_6 = ~DecoderUnit_io_instBuffer_inst_1_ready; // @[Core.scala 77:7]
  wire  _T_7 = Ctrl_io_decoderUnit_branch_flag & _T_6; // @[Core.scala 75:8]
  wire  _T_13 = ~DecoderUnit_io_executeStage_inst0_ex_bd & Ctrl_io_executeUnit_do_flush &
    Ctrl_io_executeUnit_allow_to_go; // @[Core.scala 114:72]
  wire  _T_14 = Ctrl_io_memoryUnit_flush_req | _T_13; // @[Core.scala 113:59]
  wire  _T_16 = ~Ctrl_io_decoderUnit_allow_to_go & Ctrl_io_executeUnit_allow_to_go; // @[Core.scala 115:35]
  wire  _T_18 = Ctrl_io_executeUnit_do_flush & DecoderUnit_io_executeStage_inst1_allow_to_go; // @[Core.scala 117:32]
  wire  _T_19 = Ctrl_io_memoryUnit_flush_req | _T_18; // @[Core.scala 116:59]
  wire  _T_21 = Ctrl_io_executeUnit_allow_to_go & ~DecoderUnit_io_executeStage_inst1_allow_to_go; // @[Core.scala 118:35]
  Ctrl Ctrl ( // @[Core.scala 24:30]
    .io_cacheCtrl_iCache_stall(Ctrl_io_cacheCtrl_iCache_stall),
    .io_cacheCtrl_dCache_stall(Ctrl_io_cacheCtrl_dCache_stall),
    .io_fetchUnit_allow_to_go(Ctrl_io_fetchUnit_allow_to_go),
    .io_instBuffer_delay_slot_do_flush(Ctrl_io_instBuffer_delay_slot_do_flush),
    .io_decoderUnit_inst0_src1_ren(Ctrl_io_decoderUnit_inst0_src1_ren),
    .io_decoderUnit_inst0_src1_raddr(Ctrl_io_decoderUnit_inst0_src1_raddr),
    .io_decoderUnit_inst0_src2_ren(Ctrl_io_decoderUnit_inst0_src2_ren),
    .io_decoderUnit_inst0_src2_raddr(Ctrl_io_decoderUnit_inst0_src2_raddr),
    .io_decoderUnit_branch_flag(Ctrl_io_decoderUnit_branch_flag),
    .io_decoderUnit_allow_to_go(Ctrl_io_decoderUnit_allow_to_go),
    .io_decoderUnit_do_flush(Ctrl_io_decoderUnit_do_flush),
    .io_executeUnit_inst_0_mem_ren(Ctrl_io_executeUnit_inst_0_mem_ren),
    .io_executeUnit_inst_0_reg_waddr(Ctrl_io_executeUnit_inst_0_reg_waddr),
    .io_executeUnit_inst_1_mem_ren(Ctrl_io_executeUnit_inst_1_mem_ren),
    .io_executeUnit_inst_1_reg_waddr(Ctrl_io_executeUnit_inst_1_reg_waddr),
    .io_executeUnit_fu_stall(Ctrl_io_executeUnit_fu_stall),
    .io_executeUnit_branch_flag(Ctrl_io_executeUnit_branch_flag),
    .io_executeUnit_allow_to_go(Ctrl_io_executeUnit_allow_to_go),
    .io_executeUnit_do_flush(Ctrl_io_executeUnit_do_flush),
    .io_executeUnit_fu_allow_to_go(Ctrl_io_executeUnit_fu_allow_to_go),
    .io_executeUnit_fu_do_flush(Ctrl_io_executeUnit_fu_do_flush),
    .io_memoryUnit_flush_req(Ctrl_io_memoryUnit_flush_req),
    .io_memoryUnit_allow_to_go(Ctrl_io_memoryUnit_allow_to_go),
    .io_memoryUnit_do_flush(Ctrl_io_memoryUnit_do_flush),
    .io_writeBackUnit_allow_to_go(Ctrl_io_writeBackUnit_allow_to_go)
  );
  FetchStage FetchStage ( // @[Core.scala 25:30]
    .clock(FetchStage_clock),
    .reset(FetchStage_reset),
    .io_memory_ex(FetchStage_io_memory_ex),
    .io_memory_ex_pc(FetchStage_io_memory_ex_pc),
    .io_memory_flush(FetchStage_io_memory_flush),
    .io_memory_flush_pc(FetchStage_io_memory_flush_pc),
    .io_decoder_branch(FetchStage_io_decoder_branch),
    .io_decoder_target(FetchStage_io_decoder_target),
    .io_execute_branch(FetchStage_io_execute_branch),
    .io_execute_target(FetchStage_io_execute_target),
    .io_instBuffer_full(FetchStage_io_instBuffer_full),
    .io_iCache_inst_valid_0(FetchStage_io_iCache_inst_valid_0),
    .io_iCache_inst_valid_1(FetchStage_io_iCache_inst_valid_1),
    .io_iCache_pc(FetchStage_io_iCache_pc),
    .io_iCache_pc_next(FetchStage_io_iCache_pc_next)
  );
  BPU BPU ( // @[Core.scala 26:30]
    .clock(BPU_clock),
    .reset(BPU_reset),
    .io_instrD(BPU_io_instrD),
    .io_enaD(BPU_io_enaD),
    .io_pcD(BPU_io_pcD),
    .io_pc_plus4D(BPU_io_pc_plus4D),
    .io_pcE(BPU_io_pcE),
    .io_branchE(BPU_io_branchE),
    .io_actual_takeE(BPU_io_actual_takeE),
    .io_branchD(BPU_io_branchD),
    .io_pred_takeD(BPU_io_pred_takeD),
    .io_branch_targetD(BPU_io_branch_targetD)
  );
  InstBuffer InstBuffer ( // @[Core.scala 27:30]
    .clock(InstBuffer_clock),
    .reset(InstBuffer_reset),
    .io_fifo_rst(InstBuffer_io_fifo_rst),
    .io_flush_delay_slot(InstBuffer_io_flush_delay_slot),
    .io_delay_sel_rst(InstBuffer_io_delay_sel_rst),
    .io_D_delay_rst(InstBuffer_io_D_delay_rst),
    .io_E_delay_rst(InstBuffer_io_E_delay_rst),
    .io_i_stall(InstBuffer_io_i_stall),
    .io_master_is_branch(InstBuffer_io_master_is_branch),
    .io_master_is_in_delayslot_o(InstBuffer_io_master_is_in_delayslot_o),
    .io_read_en_0(InstBuffer_io_read_en_0),
    .io_read_en_1(InstBuffer_io_read_en_1),
    .io_read_0_tlb_invalid(InstBuffer_io_read_0_tlb_invalid),
    .io_read_0_data(InstBuffer_io_read_0_data),
    .io_read_0_addr(InstBuffer_io_read_0_addr),
    .io_read_1_tlb_invalid(InstBuffer_io_read_1_tlb_invalid),
    .io_read_1_data(InstBuffer_io_read_1_data),
    .io_read_1_addr(InstBuffer_io_read_1_addr),
    .io_write_en_0(InstBuffer_io_write_en_0),
    .io_write_en_1(InstBuffer_io_write_en_1),
    .io_write_0_tlb_invalid(InstBuffer_io_write_0_tlb_invalid),
    .io_write_0_data(InstBuffer_io_write_0_data),
    .io_write_0_addr(InstBuffer_io_write_0_addr),
    .io_write_1_tlb_invalid(InstBuffer_io_write_1_tlb_invalid),
    .io_write_1_data(InstBuffer_io_write_1_data),
    .io_write_1_addr(InstBuffer_io_write_1_addr),
    .io_empty(InstBuffer_io_empty),
    .io_almost_empty(InstBuffer_io_almost_empty),
    .io_full(InstBuffer_io_full)
  );
  DecoderUnit DecoderUnit ( // @[Core.scala 28:30]
    .io_instBuffer_inst_0_ready(DecoderUnit_io_instBuffer_inst_0_ready),
    .io_instBuffer_inst_0_bits_pc(DecoderUnit_io_instBuffer_inst_0_bits_pc),
    .io_instBuffer_inst_0_bits_inst(DecoderUnit_io_instBuffer_inst_0_bits_inst),
    .io_instBuffer_inst_0_bits_tlb_invalid(DecoderUnit_io_instBuffer_inst_0_bits_tlb_invalid),
    .io_instBuffer_inst_1_ready(DecoderUnit_io_instBuffer_inst_1_ready),
    .io_instBuffer_inst_1_bits_pc(DecoderUnit_io_instBuffer_inst_1_bits_pc),
    .io_instBuffer_inst_1_bits_inst(DecoderUnit_io_instBuffer_inst_1_bits_inst),
    .io_instBuffer_inst_1_bits_tlb_invalid(DecoderUnit_io_instBuffer_inst_1_bits_tlb_invalid),
    .io_instBuffer_info_inst0_is_in_delayslot(DecoderUnit_io_instBuffer_info_inst0_is_in_delayslot),
    .io_instBuffer_info_empty(DecoderUnit_io_instBuffer_info_empty),
    .io_instBuffer_info_almost_empty(DecoderUnit_io_instBuffer_info_almost_empty),
    .io_instBuffer_inst0_is_jb(DecoderUnit_io_instBuffer_inst0_is_jb),
    .io_regfile_0_src1_raddr(DecoderUnit_io_regfile_0_src1_raddr),
    .io_regfile_0_src1_rdata(DecoderUnit_io_regfile_0_src1_rdata),
    .io_regfile_0_src2_raddr(DecoderUnit_io_regfile_0_src2_raddr),
    .io_regfile_0_src2_rdata(DecoderUnit_io_regfile_0_src2_rdata),
    .io_regfile_1_src1_raddr(DecoderUnit_io_regfile_1_src1_raddr),
    .io_regfile_1_src1_rdata(DecoderUnit_io_regfile_1_src1_rdata),
    .io_regfile_1_src2_raddr(DecoderUnit_io_regfile_1_src2_raddr),
    .io_regfile_1_src2_rdata(DecoderUnit_io_regfile_1_src2_rdata),
    .io_forward_0_exe_wen(DecoderUnit_io_forward_0_exe_wen),
    .io_forward_0_exe_waddr(DecoderUnit_io_forward_0_exe_waddr),
    .io_forward_0_exe_wdata(DecoderUnit_io_forward_0_exe_wdata),
    .io_forward_0_exe_mem_ren(DecoderUnit_io_forward_0_exe_mem_ren),
    .io_forward_0_mem_wen(DecoderUnit_io_forward_0_mem_wen),
    .io_forward_0_mem_waddr(DecoderUnit_io_forward_0_mem_waddr),
    .io_forward_0_mem_wdata(DecoderUnit_io_forward_0_mem_wdata),
    .io_forward_1_exe_wen(DecoderUnit_io_forward_1_exe_wen),
    .io_forward_1_exe_waddr(DecoderUnit_io_forward_1_exe_waddr),
    .io_forward_1_exe_wdata(DecoderUnit_io_forward_1_exe_wdata),
    .io_forward_1_exe_mem_ren(DecoderUnit_io_forward_1_exe_mem_ren),
    .io_forward_1_mem_wen(DecoderUnit_io_forward_1_mem_wen),
    .io_forward_1_mem_waddr(DecoderUnit_io_forward_1_mem_waddr),
    .io_forward_1_mem_wdata(DecoderUnit_io_forward_1_mem_wdata),
    .io_cp0_access_allowed(DecoderUnit_io_cp0_access_allowed),
    .io_cp0_kernel_mode(DecoderUnit_io_cp0_kernel_mode),
    .io_cp0_intterupt_allowed(DecoderUnit_io_cp0_intterupt_allowed),
    .io_cp0_cause_ip(DecoderUnit_io_cp0_cause_ip),
    .io_cp0_status_im(DecoderUnit_io_cp0_status_im),
    .io_fetchUnit_branch(DecoderUnit_io_fetchUnit_branch),
    .io_fetchUnit_target(DecoderUnit_io_fetchUnit_target),
    .io_bpu_pc(DecoderUnit_io_bpu_pc),
    .io_bpu_decoded_inst0_inst(DecoderUnit_io_bpu_decoded_inst0_inst),
    .io_bpu_inst_is_branch(DecoderUnit_io_bpu_inst_is_branch),
    .io_bpu_pred_branch_flag(DecoderUnit_io_bpu_pred_branch_flag),
    .io_bpu_branch_target(DecoderUnit_io_bpu_branch_target),
    .io_executeStage_inst0_pc(DecoderUnit_io_executeStage_inst0_pc),
    .io_executeStage_inst0_inst_info_fusel(DecoderUnit_io_executeStage_inst0_inst_info_fusel),
    .io_executeStage_inst0_inst_info_op(DecoderUnit_io_executeStage_inst0_inst_info_op),
    .io_executeStage_inst0_inst_info_reg_wen(DecoderUnit_io_executeStage_inst0_inst_info_reg_wen),
    .io_executeStage_inst0_inst_info_reg_waddr(DecoderUnit_io_executeStage_inst0_inst_info_reg_waddr),
    .io_executeStage_inst0_inst_info_cp0_addr(DecoderUnit_io_executeStage_inst0_inst_info_cp0_addr),
    .io_executeStage_inst0_inst_info_inst(DecoderUnit_io_executeStage_inst0_inst_info_inst),
    .io_executeStage_inst0_src_info_src1_data(DecoderUnit_io_executeStage_inst0_src_info_src1_data),
    .io_executeStage_inst0_src_info_src2_data(DecoderUnit_io_executeStage_inst0_src_info_src2_data),
    .io_executeStage_inst0_ex_flush_req(DecoderUnit_io_executeStage_inst0_ex_flush_req),
    .io_executeStage_inst0_ex_tlb_refill(DecoderUnit_io_executeStage_inst0_ex_tlb_refill),
    .io_executeStage_inst0_ex_eret(DecoderUnit_io_executeStage_inst0_ex_eret),
    .io_executeStage_inst0_ex_badvaddr(DecoderUnit_io_executeStage_inst0_ex_badvaddr),
    .io_executeStage_inst0_ex_bd(DecoderUnit_io_executeStage_inst0_ex_bd),
    .io_executeStage_inst0_ex_excode(DecoderUnit_io_executeStage_inst0_ex_excode),
    .io_executeStage_inst0_jb_info_jump_regiser_conflict(DecoderUnit_io_executeStage_inst0_jb_info_jump_regiser_conflict
      ),
    .io_executeStage_inst0_jb_info_is_branch(DecoderUnit_io_executeStage_inst0_jb_info_is_branch),
    .io_executeStage_inst0_jb_info_pred_branch_flag(DecoderUnit_io_executeStage_inst0_jb_info_pred_branch_flag),
    .io_executeStage_inst0_jb_info_branch_target(DecoderUnit_io_executeStage_inst0_jb_info_branch_target),
    .io_executeStage_inst1_allow_to_go(DecoderUnit_io_executeStage_inst1_allow_to_go),
    .io_executeStage_inst1_pc(DecoderUnit_io_executeStage_inst1_pc),
    .io_executeStage_inst1_inst_info_fusel(DecoderUnit_io_executeStage_inst1_inst_info_fusel),
    .io_executeStage_inst1_inst_info_op(DecoderUnit_io_executeStage_inst1_inst_info_op),
    .io_executeStage_inst1_inst_info_reg_wen(DecoderUnit_io_executeStage_inst1_inst_info_reg_wen),
    .io_executeStage_inst1_inst_info_reg_waddr(DecoderUnit_io_executeStage_inst1_inst_info_reg_waddr),
    .io_executeStage_inst1_inst_info_inst(DecoderUnit_io_executeStage_inst1_inst_info_inst),
    .io_executeStage_inst1_src_info_src1_data(DecoderUnit_io_executeStage_inst1_src_info_src1_data),
    .io_executeStage_inst1_src_info_src2_data(DecoderUnit_io_executeStage_inst1_src_info_src2_data),
    .io_executeStage_inst1_ex_flush_req(DecoderUnit_io_executeStage_inst1_ex_flush_req),
    .io_executeStage_inst1_ex_tlb_refill(DecoderUnit_io_executeStage_inst1_ex_tlb_refill),
    .io_executeStage_inst1_ex_eret(DecoderUnit_io_executeStage_inst1_ex_eret),
    .io_executeStage_inst1_ex_badvaddr(DecoderUnit_io_executeStage_inst1_ex_badvaddr),
    .io_executeStage_inst1_ex_bd(DecoderUnit_io_executeStage_inst1_ex_bd),
    .io_executeStage_inst1_ex_excode(DecoderUnit_io_executeStage_inst1_ex_excode),
    .io_ctrl_inst0_src1_ren(DecoderUnit_io_ctrl_inst0_src1_ren),
    .io_ctrl_inst0_src1_raddr(DecoderUnit_io_ctrl_inst0_src1_raddr),
    .io_ctrl_inst0_src2_ren(DecoderUnit_io_ctrl_inst0_src2_ren),
    .io_ctrl_inst0_src2_raddr(DecoderUnit_io_ctrl_inst0_src2_raddr),
    .io_ctrl_branch_flag(DecoderUnit_io_ctrl_branch_flag),
    .io_ctrl_allow_to_go(DecoderUnit_io_ctrl_allow_to_go)
  );
  ARegFile ARegFile ( // @[Core.scala 29:30]
    .clock(ARegFile_clock),
    .reset(ARegFile_reset),
    .io_read_0_src1_raddr(ARegFile_io_read_0_src1_raddr),
    .io_read_0_src1_rdata(ARegFile_io_read_0_src1_rdata),
    .io_read_0_src2_raddr(ARegFile_io_read_0_src2_raddr),
    .io_read_0_src2_rdata(ARegFile_io_read_0_src2_rdata),
    .io_read_1_src1_raddr(ARegFile_io_read_1_src1_raddr),
    .io_read_1_src1_rdata(ARegFile_io_read_1_src1_rdata),
    .io_read_1_src2_raddr(ARegFile_io_read_1_src2_raddr),
    .io_read_1_src2_rdata(ARegFile_io_read_1_src2_rdata),
    .io_write_0_wen(ARegFile_io_write_0_wen),
    .io_write_0_waddr(ARegFile_io_write_0_waddr),
    .io_write_0_wdata(ARegFile_io_write_0_wdata),
    .io_write_1_wen(ARegFile_io_write_1_wen),
    .io_write_1_waddr(ARegFile_io_write_1_waddr),
    .io_write_1_wdata(ARegFile_io_write_1_wdata)
  );
  ExecuteStage ExecuteStage ( // @[Core.scala 30:30]
    .clock(ExecuteStage_clock),
    .reset(ExecuteStage_reset),
    .io_ctrl_inst0_allow_to_go(ExecuteStage_io_ctrl_inst0_allow_to_go),
    .io_ctrl_clear_0(ExecuteStage_io_ctrl_clear_0),
    .io_ctrl_clear_1(ExecuteStage_io_ctrl_clear_1),
    .io_decoderUnit_inst0_pc(ExecuteStage_io_decoderUnit_inst0_pc),
    .io_decoderUnit_inst0_inst_info_fusel(ExecuteStage_io_decoderUnit_inst0_inst_info_fusel),
    .io_decoderUnit_inst0_inst_info_op(ExecuteStage_io_decoderUnit_inst0_inst_info_op),
    .io_decoderUnit_inst0_inst_info_reg_wen(ExecuteStage_io_decoderUnit_inst0_inst_info_reg_wen),
    .io_decoderUnit_inst0_inst_info_reg_waddr(ExecuteStage_io_decoderUnit_inst0_inst_info_reg_waddr),
    .io_decoderUnit_inst0_inst_info_cp0_addr(ExecuteStage_io_decoderUnit_inst0_inst_info_cp0_addr),
    .io_decoderUnit_inst0_inst_info_inst(ExecuteStage_io_decoderUnit_inst0_inst_info_inst),
    .io_decoderUnit_inst0_src_info_src1_data(ExecuteStage_io_decoderUnit_inst0_src_info_src1_data),
    .io_decoderUnit_inst0_src_info_src2_data(ExecuteStage_io_decoderUnit_inst0_src_info_src2_data),
    .io_decoderUnit_inst0_ex_flush_req(ExecuteStage_io_decoderUnit_inst0_ex_flush_req),
    .io_decoderUnit_inst0_ex_eret(ExecuteStage_io_decoderUnit_inst0_ex_eret),
    .io_decoderUnit_inst0_ex_badvaddr(ExecuteStage_io_decoderUnit_inst0_ex_badvaddr),
    .io_decoderUnit_inst0_ex_bd(ExecuteStage_io_decoderUnit_inst0_ex_bd),
    .io_decoderUnit_inst0_ex_excode(ExecuteStage_io_decoderUnit_inst0_ex_excode),
    .io_decoderUnit_inst0_jb_info_jump_regiser_conflict(ExecuteStage_io_decoderUnit_inst0_jb_info_jump_regiser_conflict)
      ,
    .io_decoderUnit_inst0_jb_info_is_branch(ExecuteStage_io_decoderUnit_inst0_jb_info_is_branch),
    .io_decoderUnit_inst0_jb_info_pred_branch_flag(ExecuteStage_io_decoderUnit_inst0_jb_info_pred_branch_flag),
    .io_decoderUnit_inst0_jb_info_branch_target(ExecuteStage_io_decoderUnit_inst0_jb_info_branch_target),
    .io_decoderUnit_inst1_allow_to_go(ExecuteStage_io_decoderUnit_inst1_allow_to_go),
    .io_decoderUnit_inst1_pc(ExecuteStage_io_decoderUnit_inst1_pc),
    .io_decoderUnit_inst1_inst_info_fusel(ExecuteStage_io_decoderUnit_inst1_inst_info_fusel),
    .io_decoderUnit_inst1_inst_info_op(ExecuteStage_io_decoderUnit_inst1_inst_info_op),
    .io_decoderUnit_inst1_inst_info_reg_wen(ExecuteStage_io_decoderUnit_inst1_inst_info_reg_wen),
    .io_decoderUnit_inst1_inst_info_reg_waddr(ExecuteStage_io_decoderUnit_inst1_inst_info_reg_waddr),
    .io_decoderUnit_inst1_inst_info_inst(ExecuteStage_io_decoderUnit_inst1_inst_info_inst),
    .io_decoderUnit_inst1_src_info_src1_data(ExecuteStage_io_decoderUnit_inst1_src_info_src1_data),
    .io_decoderUnit_inst1_src_info_src2_data(ExecuteStage_io_decoderUnit_inst1_src_info_src2_data),
    .io_decoderUnit_inst1_ex_flush_req(ExecuteStage_io_decoderUnit_inst1_ex_flush_req),
    .io_decoderUnit_inst1_ex_eret(ExecuteStage_io_decoderUnit_inst1_ex_eret),
    .io_decoderUnit_inst1_ex_badvaddr(ExecuteStage_io_decoderUnit_inst1_ex_badvaddr),
    .io_decoderUnit_inst1_ex_bd(ExecuteStage_io_decoderUnit_inst1_ex_bd),
    .io_decoderUnit_inst1_ex_excode(ExecuteStage_io_decoderUnit_inst1_ex_excode),
    .io_executeUnit_inst0_pc(ExecuteStage_io_executeUnit_inst0_pc),
    .io_executeUnit_inst0_inst_info_fusel(ExecuteStage_io_executeUnit_inst0_inst_info_fusel),
    .io_executeUnit_inst0_inst_info_op(ExecuteStage_io_executeUnit_inst0_inst_info_op),
    .io_executeUnit_inst0_inst_info_reg_wen(ExecuteStage_io_executeUnit_inst0_inst_info_reg_wen),
    .io_executeUnit_inst0_inst_info_reg_waddr(ExecuteStage_io_executeUnit_inst0_inst_info_reg_waddr),
    .io_executeUnit_inst0_inst_info_cp0_addr(ExecuteStage_io_executeUnit_inst0_inst_info_cp0_addr),
    .io_executeUnit_inst0_inst_info_inst(ExecuteStage_io_executeUnit_inst0_inst_info_inst),
    .io_executeUnit_inst0_src_info_src1_data(ExecuteStage_io_executeUnit_inst0_src_info_src1_data),
    .io_executeUnit_inst0_src_info_src2_data(ExecuteStage_io_executeUnit_inst0_src_info_src2_data),
    .io_executeUnit_inst0_ex_flush_req(ExecuteStage_io_executeUnit_inst0_ex_flush_req),
    .io_executeUnit_inst0_ex_eret(ExecuteStage_io_executeUnit_inst0_ex_eret),
    .io_executeUnit_inst0_ex_badvaddr(ExecuteStage_io_executeUnit_inst0_ex_badvaddr),
    .io_executeUnit_inst0_ex_bd(ExecuteStage_io_executeUnit_inst0_ex_bd),
    .io_executeUnit_inst0_ex_excode(ExecuteStage_io_executeUnit_inst0_ex_excode),
    .io_executeUnit_inst0_jb_info_jump_regiser_conflict(ExecuteStage_io_executeUnit_inst0_jb_info_jump_regiser_conflict)
      ,
    .io_executeUnit_inst0_jb_info_is_branch(ExecuteStage_io_executeUnit_inst0_jb_info_is_branch),
    .io_executeUnit_inst0_jb_info_pred_branch_flag(ExecuteStage_io_executeUnit_inst0_jb_info_pred_branch_flag),
    .io_executeUnit_inst0_jb_info_branch_target(ExecuteStage_io_executeUnit_inst0_jb_info_branch_target),
    .io_executeUnit_inst1_pc(ExecuteStage_io_executeUnit_inst1_pc),
    .io_executeUnit_inst1_inst_info_fusel(ExecuteStage_io_executeUnit_inst1_inst_info_fusel),
    .io_executeUnit_inst1_inst_info_op(ExecuteStage_io_executeUnit_inst1_inst_info_op),
    .io_executeUnit_inst1_inst_info_reg_wen(ExecuteStage_io_executeUnit_inst1_inst_info_reg_wen),
    .io_executeUnit_inst1_inst_info_reg_waddr(ExecuteStage_io_executeUnit_inst1_inst_info_reg_waddr),
    .io_executeUnit_inst1_inst_info_inst(ExecuteStage_io_executeUnit_inst1_inst_info_inst),
    .io_executeUnit_inst1_src_info_src1_data(ExecuteStage_io_executeUnit_inst1_src_info_src1_data),
    .io_executeUnit_inst1_src_info_src2_data(ExecuteStage_io_executeUnit_inst1_src_info_src2_data),
    .io_executeUnit_inst1_ex_flush_req(ExecuteStage_io_executeUnit_inst1_ex_flush_req),
    .io_executeUnit_inst1_ex_eret(ExecuteStage_io_executeUnit_inst1_ex_eret),
    .io_executeUnit_inst1_ex_badvaddr(ExecuteStage_io_executeUnit_inst1_ex_badvaddr),
    .io_executeUnit_inst1_ex_bd(ExecuteStage_io_executeUnit_inst1_ex_bd),
    .io_executeUnit_inst1_ex_excode(ExecuteStage_io_executeUnit_inst1_ex_excode)
  );
  ExecuteUnit ExecuteUnit ( // @[Core.scala 31:30]
    .clock(ExecuteUnit_clock),
    .reset(ExecuteUnit_reset),
    .io_ctrl_inst_0_mem_ren(ExecuteUnit_io_ctrl_inst_0_mem_ren),
    .io_ctrl_inst_0_reg_waddr(ExecuteUnit_io_ctrl_inst_0_reg_waddr),
    .io_ctrl_inst_1_mem_ren(ExecuteUnit_io_ctrl_inst_1_mem_ren),
    .io_ctrl_inst_1_reg_waddr(ExecuteUnit_io_ctrl_inst_1_reg_waddr),
    .io_ctrl_fu_stall(ExecuteUnit_io_ctrl_fu_stall),
    .io_ctrl_branch_flag(ExecuteUnit_io_ctrl_branch_flag),
    .io_ctrl_allow_to_go(ExecuteUnit_io_ctrl_allow_to_go),
    .io_ctrl_fu_allow_to_go(ExecuteUnit_io_ctrl_fu_allow_to_go),
    .io_ctrl_fu_do_flush(ExecuteUnit_io_ctrl_fu_do_flush),
    .io_executeStage_inst0_pc(ExecuteUnit_io_executeStage_inst0_pc),
    .io_executeStage_inst0_inst_info_fusel(ExecuteUnit_io_executeStage_inst0_inst_info_fusel),
    .io_executeStage_inst0_inst_info_op(ExecuteUnit_io_executeStage_inst0_inst_info_op),
    .io_executeStage_inst0_inst_info_reg_wen(ExecuteUnit_io_executeStage_inst0_inst_info_reg_wen),
    .io_executeStage_inst0_inst_info_reg_waddr(ExecuteUnit_io_executeStage_inst0_inst_info_reg_waddr),
    .io_executeStage_inst0_inst_info_cp0_addr(ExecuteUnit_io_executeStage_inst0_inst_info_cp0_addr),
    .io_executeStage_inst0_inst_info_inst(ExecuteUnit_io_executeStage_inst0_inst_info_inst),
    .io_executeStage_inst0_src_info_src1_data(ExecuteUnit_io_executeStage_inst0_src_info_src1_data),
    .io_executeStage_inst0_src_info_src2_data(ExecuteUnit_io_executeStage_inst0_src_info_src2_data),
    .io_executeStage_inst0_ex_flush_req(ExecuteUnit_io_executeStage_inst0_ex_flush_req),
    .io_executeStage_inst0_ex_eret(ExecuteUnit_io_executeStage_inst0_ex_eret),
    .io_executeStage_inst0_ex_badvaddr(ExecuteUnit_io_executeStage_inst0_ex_badvaddr),
    .io_executeStage_inst0_ex_bd(ExecuteUnit_io_executeStage_inst0_ex_bd),
    .io_executeStage_inst0_ex_excode(ExecuteUnit_io_executeStage_inst0_ex_excode),
    .io_executeStage_inst0_jb_info_jump_regiser_conflict(ExecuteUnit_io_executeStage_inst0_jb_info_jump_regiser_conflict
      ),
    .io_executeStage_inst0_jb_info_is_branch(ExecuteUnit_io_executeStage_inst0_jb_info_is_branch),
    .io_executeStage_inst0_jb_info_pred_branch_flag(ExecuteUnit_io_executeStage_inst0_jb_info_pred_branch_flag),
    .io_executeStage_inst0_jb_info_branch_target(ExecuteUnit_io_executeStage_inst0_jb_info_branch_target),
    .io_executeStage_inst1_pc(ExecuteUnit_io_executeStage_inst1_pc),
    .io_executeStage_inst1_inst_info_fusel(ExecuteUnit_io_executeStage_inst1_inst_info_fusel),
    .io_executeStage_inst1_inst_info_op(ExecuteUnit_io_executeStage_inst1_inst_info_op),
    .io_executeStage_inst1_inst_info_reg_wen(ExecuteUnit_io_executeStage_inst1_inst_info_reg_wen),
    .io_executeStage_inst1_inst_info_reg_waddr(ExecuteUnit_io_executeStage_inst1_inst_info_reg_waddr),
    .io_executeStage_inst1_inst_info_inst(ExecuteUnit_io_executeStage_inst1_inst_info_inst),
    .io_executeStage_inst1_src_info_src1_data(ExecuteUnit_io_executeStage_inst1_src_info_src1_data),
    .io_executeStage_inst1_src_info_src2_data(ExecuteUnit_io_executeStage_inst1_src_info_src2_data),
    .io_executeStage_inst1_ex_flush_req(ExecuteUnit_io_executeStage_inst1_ex_flush_req),
    .io_executeStage_inst1_ex_eret(ExecuteUnit_io_executeStage_inst1_ex_eret),
    .io_executeStage_inst1_ex_badvaddr(ExecuteUnit_io_executeStage_inst1_ex_badvaddr),
    .io_executeStage_inst1_ex_bd(ExecuteUnit_io_executeStage_inst1_ex_bd),
    .io_executeStage_inst1_ex_excode(ExecuteUnit_io_executeStage_inst1_ex_excode),
    .io_cp0_in_inst_info_op(ExecuteUnit_io_cp0_in_inst_info_op),
    .io_cp0_in_inst_info_cp0_addr(ExecuteUnit_io_cp0_in_inst_info_cp0_addr),
    .io_cp0_in_mtc0_wdata(ExecuteUnit_io_cp0_in_mtc0_wdata),
    .io_cp0_out_cp0_rdata(ExecuteUnit_io_cp0_out_cp0_rdata),
    .io_cp0_out_debug_cp0_count(ExecuteUnit_io_cp0_out_debug_cp0_count),
    .io_cp0_out_debug_cp0_random(ExecuteUnit_io_cp0_out_debug_cp0_random),
    .io_cp0_out_debug_cp0_cause(ExecuteUnit_io_cp0_out_debug_cp0_cause),
    .io_bpu_pc(ExecuteUnit_io_bpu_pc),
    .io_bpu_branch_flag(ExecuteUnit_io_bpu_branch_flag),
    .io_bpu_inst0_is_branch(ExecuteUnit_io_bpu_inst0_is_branch),
    .io_fetchStage_branch(ExecuteUnit_io_fetchStage_branch),
    .io_fetchStage_target(ExecuteUnit_io_fetchStage_target),
    .io_decoderUnit_forward_0_exe_wen(ExecuteUnit_io_decoderUnit_forward_0_exe_wen),
    .io_decoderUnit_forward_0_exe_waddr(ExecuteUnit_io_decoderUnit_forward_0_exe_waddr),
    .io_decoderUnit_forward_0_exe_wdata(ExecuteUnit_io_decoderUnit_forward_0_exe_wdata),
    .io_decoderUnit_forward_0_exe_mem_ren(ExecuteUnit_io_decoderUnit_forward_0_exe_mem_ren),
    .io_decoderUnit_forward_1_exe_wen(ExecuteUnit_io_decoderUnit_forward_1_exe_wen),
    .io_decoderUnit_forward_1_exe_waddr(ExecuteUnit_io_decoderUnit_forward_1_exe_waddr),
    .io_decoderUnit_forward_1_exe_wdata(ExecuteUnit_io_decoderUnit_forward_1_exe_wdata),
    .io_decoderUnit_forward_1_exe_mem_ren(ExecuteUnit_io_decoderUnit_forward_1_exe_mem_ren),
    .io_decoderUnit_inst0_bd(ExecuteUnit_io_decoderUnit_inst0_bd),
    .io_memoryStage_inst0_pc(ExecuteUnit_io_memoryStage_inst0_pc),
    .io_memoryStage_inst0_inst_info_fusel(ExecuteUnit_io_memoryStage_inst0_inst_info_fusel),
    .io_memoryStage_inst0_inst_info_op(ExecuteUnit_io_memoryStage_inst0_inst_info_op),
    .io_memoryStage_inst0_inst_info_reg_wen(ExecuteUnit_io_memoryStage_inst0_inst_info_reg_wen),
    .io_memoryStage_inst0_inst_info_reg_waddr(ExecuteUnit_io_memoryStage_inst0_inst_info_reg_waddr),
    .io_memoryStage_inst0_inst_info_inst(ExecuteUnit_io_memoryStage_inst0_inst_info_inst),
    .io_memoryStage_inst0_rd_info_wdata(ExecuteUnit_io_memoryStage_inst0_rd_info_wdata),
    .io_memoryStage_inst0_ex_flush_req(ExecuteUnit_io_memoryStage_inst0_ex_flush_req),
    .io_memoryStage_inst0_ex_eret(ExecuteUnit_io_memoryStage_inst0_ex_eret),
    .io_memoryStage_inst0_ex_badvaddr(ExecuteUnit_io_memoryStage_inst0_ex_badvaddr),
    .io_memoryStage_inst0_ex_bd(ExecuteUnit_io_memoryStage_inst0_ex_bd),
    .io_memoryStage_inst0_ex_excode(ExecuteUnit_io_memoryStage_inst0_ex_excode),
    .io_memoryStage_inst0_cp0_cp0_count(ExecuteUnit_io_memoryStage_inst0_cp0_cp0_count),
    .io_memoryStage_inst0_cp0_cp0_random(ExecuteUnit_io_memoryStage_inst0_cp0_cp0_random),
    .io_memoryStage_inst0_cp0_cp0_cause(ExecuteUnit_io_memoryStage_inst0_cp0_cp0_cause),
    .io_memoryStage_inst0_mem_en(ExecuteUnit_io_memoryStage_inst0_mem_en),
    .io_memoryStage_inst0_mem_inst_info_op(ExecuteUnit_io_memoryStage_inst0_mem_inst_info_op),
    .io_memoryStage_inst0_mem_addr(ExecuteUnit_io_memoryStage_inst0_mem_addr),
    .io_memoryStage_inst0_mem_wdata(ExecuteUnit_io_memoryStage_inst0_mem_wdata),
    .io_memoryStage_inst0_mem_sel_0(ExecuteUnit_io_memoryStage_inst0_mem_sel_0),
    .io_memoryStage_inst0_mem_sel_1(ExecuteUnit_io_memoryStage_inst0_mem_sel_1),
    .io_memoryStage_inst1_pc(ExecuteUnit_io_memoryStage_inst1_pc),
    .io_memoryStage_inst1_inst_info_fusel(ExecuteUnit_io_memoryStage_inst1_inst_info_fusel),
    .io_memoryStage_inst1_inst_info_reg_wen(ExecuteUnit_io_memoryStage_inst1_inst_info_reg_wen),
    .io_memoryStage_inst1_inst_info_reg_waddr(ExecuteUnit_io_memoryStage_inst1_inst_info_reg_waddr),
    .io_memoryStage_inst1_rd_info_wdata(ExecuteUnit_io_memoryStage_inst1_rd_info_wdata),
    .io_memoryStage_inst1_ex_flush_req(ExecuteUnit_io_memoryStage_inst1_ex_flush_req),
    .io_memoryStage_inst1_ex_eret(ExecuteUnit_io_memoryStage_inst1_ex_eret),
    .io_memoryStage_inst1_ex_badvaddr(ExecuteUnit_io_memoryStage_inst1_ex_badvaddr),
    .io_memoryStage_inst1_ex_bd(ExecuteUnit_io_memoryStage_inst1_ex_bd),
    .io_memoryStage_inst1_ex_excode(ExecuteUnit_io_memoryStage_inst1_ex_excode)
  );
  Cp0 Cp0 ( // @[Core.scala 32:30]
    .clock(Cp0_clock),
    .reset(Cp0_reset),
    .io_ext_int(Cp0_io_ext_int),
    .io_ctrl_exe_stall(Cp0_io_ctrl_exe_stall),
    .io_ctrl_mem_stall(Cp0_io_ctrl_mem_stall),
    .io_decoderUnit_access_allowed(Cp0_io_decoderUnit_access_allowed),
    .io_decoderUnit_kernel_mode(Cp0_io_decoderUnit_kernel_mode),
    .io_decoderUnit_intterupt_allowed(Cp0_io_decoderUnit_intterupt_allowed),
    .io_decoderUnit_cause_ip(Cp0_io_decoderUnit_cause_ip),
    .io_decoderUnit_status_im(Cp0_io_decoderUnit_status_im),
    .io_executeUnit_in_inst_info_op(Cp0_io_executeUnit_in_inst_info_op),
    .io_executeUnit_in_inst_info_cp0_addr(Cp0_io_executeUnit_in_inst_info_cp0_addr),
    .io_executeUnit_in_mtc0_wdata(Cp0_io_executeUnit_in_mtc0_wdata),
    .io_executeUnit_out_cp0_rdata(Cp0_io_executeUnit_out_cp0_rdata),
    .io_executeUnit_out_debug_cp0_count(Cp0_io_executeUnit_out_debug_cp0_count),
    .io_executeUnit_out_debug_cp0_random(Cp0_io_executeUnit_out_debug_cp0_random),
    .io_executeUnit_out_debug_cp0_cause(Cp0_io_executeUnit_out_debug_cp0_cause),
    .io_memoryUnit_in_inst_0_pc(Cp0_io_memoryUnit_in_inst_0_pc),
    .io_memoryUnit_in_inst_0_ex_flush_req(Cp0_io_memoryUnit_in_inst_0_ex_flush_req),
    .io_memoryUnit_in_inst_0_ex_tlb_refill(Cp0_io_memoryUnit_in_inst_0_ex_tlb_refill),
    .io_memoryUnit_in_inst_0_ex_eret(Cp0_io_memoryUnit_in_inst_0_ex_eret),
    .io_memoryUnit_in_inst_0_ex_badvaddr(Cp0_io_memoryUnit_in_inst_0_ex_badvaddr),
    .io_memoryUnit_in_inst_0_ex_bd(Cp0_io_memoryUnit_in_inst_0_ex_bd),
    .io_memoryUnit_in_inst_0_ex_excode(Cp0_io_memoryUnit_in_inst_0_ex_excode),
    .io_memoryUnit_in_inst_1_pc(Cp0_io_memoryUnit_in_inst_1_pc),
    .io_memoryUnit_in_inst_1_ex_flush_req(Cp0_io_memoryUnit_in_inst_1_ex_flush_req),
    .io_memoryUnit_in_inst_1_ex_tlb_refill(Cp0_io_memoryUnit_in_inst_1_ex_tlb_refill),
    .io_memoryUnit_in_inst_1_ex_eret(Cp0_io_memoryUnit_in_inst_1_ex_eret),
    .io_memoryUnit_in_inst_1_ex_badvaddr(Cp0_io_memoryUnit_in_inst_1_ex_badvaddr),
    .io_memoryUnit_in_inst_1_ex_bd(Cp0_io_memoryUnit_in_inst_1_ex_bd),
    .io_memoryUnit_in_inst_1_ex_excode(Cp0_io_memoryUnit_in_inst_1_ex_excode),
    .io_memoryUnit_out_flush(Cp0_io_memoryUnit_out_flush),
    .io_memoryUnit_out_flush_pc(Cp0_io_memoryUnit_out_flush_pc),
    .io_tlb_0_vpn2(Cp0_io_tlb_0_vpn2),
    .io_tlb_0_found(Cp0_io_tlb_0_found),
    .io_tlb_0_info_pfn_0(Cp0_io_tlb_0_info_pfn_0),
    .io_tlb_0_info_pfn_1(Cp0_io_tlb_0_info_pfn_1),
    .io_tlb_0_info_c_0(Cp0_io_tlb_0_info_c_0),
    .io_tlb_0_info_c_1(Cp0_io_tlb_0_info_c_1),
    .io_tlb_0_info_v_0(Cp0_io_tlb_0_info_v_0),
    .io_tlb_0_info_v_1(Cp0_io_tlb_0_info_v_1),
    .io_tlb_1_vpn2(Cp0_io_tlb_1_vpn2),
    .io_tlb_1_found(Cp0_io_tlb_1_found),
    .io_tlb_1_info_pfn_0(Cp0_io_tlb_1_info_pfn_0),
    .io_tlb_1_info_pfn_1(Cp0_io_tlb_1_info_pfn_1),
    .io_tlb_1_info_c_0(Cp0_io_tlb_1_info_c_0),
    .io_tlb_1_info_c_1(Cp0_io_tlb_1_info_c_1),
    .io_tlb_1_info_d_0(Cp0_io_tlb_1_info_d_0),
    .io_tlb_1_info_d_1(Cp0_io_tlb_1_info_d_1),
    .io_tlb_1_info_v_0(Cp0_io_tlb_1_info_v_0),
    .io_tlb_1_info_v_1(Cp0_io_tlb_1_info_v_1)
  );
  MemoryStage MemoryStage ( // @[Core.scala 33:30]
    .clock(MemoryStage_clock),
    .reset(MemoryStage_reset),
    .io_ctrl_allow_to_go(MemoryStage_io_ctrl_allow_to_go),
    .io_ctrl_clear_0(MemoryStage_io_ctrl_clear_0),
    .io_ctrl_clear_1(MemoryStage_io_ctrl_clear_1),
    .io_executeUnit_inst0_pc(MemoryStage_io_executeUnit_inst0_pc),
    .io_executeUnit_inst0_inst_info_fusel(MemoryStage_io_executeUnit_inst0_inst_info_fusel),
    .io_executeUnit_inst0_inst_info_op(MemoryStage_io_executeUnit_inst0_inst_info_op),
    .io_executeUnit_inst0_inst_info_reg_wen(MemoryStage_io_executeUnit_inst0_inst_info_reg_wen),
    .io_executeUnit_inst0_inst_info_reg_waddr(MemoryStage_io_executeUnit_inst0_inst_info_reg_waddr),
    .io_executeUnit_inst0_inst_info_inst(MemoryStage_io_executeUnit_inst0_inst_info_inst),
    .io_executeUnit_inst0_rd_info_wdata(MemoryStage_io_executeUnit_inst0_rd_info_wdata),
    .io_executeUnit_inst0_ex_flush_req(MemoryStage_io_executeUnit_inst0_ex_flush_req),
    .io_executeUnit_inst0_ex_eret(MemoryStage_io_executeUnit_inst0_ex_eret),
    .io_executeUnit_inst0_ex_badvaddr(MemoryStage_io_executeUnit_inst0_ex_badvaddr),
    .io_executeUnit_inst0_ex_bd(MemoryStage_io_executeUnit_inst0_ex_bd),
    .io_executeUnit_inst0_ex_excode(MemoryStage_io_executeUnit_inst0_ex_excode),
    .io_executeUnit_inst0_cp0_cp0_count(MemoryStage_io_executeUnit_inst0_cp0_cp0_count),
    .io_executeUnit_inst0_cp0_cp0_random(MemoryStage_io_executeUnit_inst0_cp0_cp0_random),
    .io_executeUnit_inst0_cp0_cp0_cause(MemoryStage_io_executeUnit_inst0_cp0_cp0_cause),
    .io_executeUnit_inst0_mem_en(MemoryStage_io_executeUnit_inst0_mem_en),
    .io_executeUnit_inst0_mem_inst_info_op(MemoryStage_io_executeUnit_inst0_mem_inst_info_op),
    .io_executeUnit_inst0_mem_addr(MemoryStage_io_executeUnit_inst0_mem_addr),
    .io_executeUnit_inst0_mem_wdata(MemoryStage_io_executeUnit_inst0_mem_wdata),
    .io_executeUnit_inst0_mem_sel_0(MemoryStage_io_executeUnit_inst0_mem_sel_0),
    .io_executeUnit_inst0_mem_sel_1(MemoryStage_io_executeUnit_inst0_mem_sel_1),
    .io_executeUnit_inst1_pc(MemoryStage_io_executeUnit_inst1_pc),
    .io_executeUnit_inst1_inst_info_fusel(MemoryStage_io_executeUnit_inst1_inst_info_fusel),
    .io_executeUnit_inst1_inst_info_reg_wen(MemoryStage_io_executeUnit_inst1_inst_info_reg_wen),
    .io_executeUnit_inst1_inst_info_reg_waddr(MemoryStage_io_executeUnit_inst1_inst_info_reg_waddr),
    .io_executeUnit_inst1_rd_info_wdata(MemoryStage_io_executeUnit_inst1_rd_info_wdata),
    .io_executeUnit_inst1_ex_flush_req(MemoryStage_io_executeUnit_inst1_ex_flush_req),
    .io_executeUnit_inst1_ex_eret(MemoryStage_io_executeUnit_inst1_ex_eret),
    .io_executeUnit_inst1_ex_badvaddr(MemoryStage_io_executeUnit_inst1_ex_badvaddr),
    .io_executeUnit_inst1_ex_bd(MemoryStage_io_executeUnit_inst1_ex_bd),
    .io_executeUnit_inst1_ex_excode(MemoryStage_io_executeUnit_inst1_ex_excode),
    .io_memoryUnit_inst0_pc(MemoryStage_io_memoryUnit_inst0_pc),
    .io_memoryUnit_inst0_inst_info_fusel(MemoryStage_io_memoryUnit_inst0_inst_info_fusel),
    .io_memoryUnit_inst0_inst_info_op(MemoryStage_io_memoryUnit_inst0_inst_info_op),
    .io_memoryUnit_inst0_inst_info_reg_wen(MemoryStage_io_memoryUnit_inst0_inst_info_reg_wen),
    .io_memoryUnit_inst0_inst_info_reg_waddr(MemoryStage_io_memoryUnit_inst0_inst_info_reg_waddr),
    .io_memoryUnit_inst0_inst_info_inst(MemoryStage_io_memoryUnit_inst0_inst_info_inst),
    .io_memoryUnit_inst0_rd_info_wdata(MemoryStage_io_memoryUnit_inst0_rd_info_wdata),
    .io_memoryUnit_inst0_ex_flush_req(MemoryStage_io_memoryUnit_inst0_ex_flush_req),
    .io_memoryUnit_inst0_ex_eret(MemoryStage_io_memoryUnit_inst0_ex_eret),
    .io_memoryUnit_inst0_ex_badvaddr(MemoryStage_io_memoryUnit_inst0_ex_badvaddr),
    .io_memoryUnit_inst0_ex_bd(MemoryStage_io_memoryUnit_inst0_ex_bd),
    .io_memoryUnit_inst0_ex_excode(MemoryStage_io_memoryUnit_inst0_ex_excode),
    .io_memoryUnit_inst0_cp0_cp0_count(MemoryStage_io_memoryUnit_inst0_cp0_cp0_count),
    .io_memoryUnit_inst0_cp0_cp0_random(MemoryStage_io_memoryUnit_inst0_cp0_cp0_random),
    .io_memoryUnit_inst0_cp0_cp0_cause(MemoryStage_io_memoryUnit_inst0_cp0_cp0_cause),
    .io_memoryUnit_inst0_mem_en(MemoryStage_io_memoryUnit_inst0_mem_en),
    .io_memoryUnit_inst0_mem_inst_info_op(MemoryStage_io_memoryUnit_inst0_mem_inst_info_op),
    .io_memoryUnit_inst0_mem_addr(MemoryStage_io_memoryUnit_inst0_mem_addr),
    .io_memoryUnit_inst0_mem_wdata(MemoryStage_io_memoryUnit_inst0_mem_wdata),
    .io_memoryUnit_inst0_mem_sel_0(MemoryStage_io_memoryUnit_inst0_mem_sel_0),
    .io_memoryUnit_inst0_mem_sel_1(MemoryStage_io_memoryUnit_inst0_mem_sel_1),
    .io_memoryUnit_inst1_pc(MemoryStage_io_memoryUnit_inst1_pc),
    .io_memoryUnit_inst1_inst_info_fusel(MemoryStage_io_memoryUnit_inst1_inst_info_fusel),
    .io_memoryUnit_inst1_inst_info_reg_wen(MemoryStage_io_memoryUnit_inst1_inst_info_reg_wen),
    .io_memoryUnit_inst1_inst_info_reg_waddr(MemoryStage_io_memoryUnit_inst1_inst_info_reg_waddr),
    .io_memoryUnit_inst1_rd_info_wdata(MemoryStage_io_memoryUnit_inst1_rd_info_wdata),
    .io_memoryUnit_inst1_ex_flush_req(MemoryStage_io_memoryUnit_inst1_ex_flush_req),
    .io_memoryUnit_inst1_ex_eret(MemoryStage_io_memoryUnit_inst1_ex_eret),
    .io_memoryUnit_inst1_ex_badvaddr(MemoryStage_io_memoryUnit_inst1_ex_badvaddr),
    .io_memoryUnit_inst1_ex_bd(MemoryStage_io_memoryUnit_inst1_ex_bd),
    .io_memoryUnit_inst1_ex_excode(MemoryStage_io_memoryUnit_inst1_ex_excode)
  );
  MemoryUnit MemoryUnit ( // @[Core.scala 34:30]
    .io_ctrl_flush_req(MemoryUnit_io_ctrl_flush_req),
    .io_ctrl_allow_to_go(MemoryUnit_io_ctrl_allow_to_go),
    .io_memoryStage_inst0_pc(MemoryUnit_io_memoryStage_inst0_pc),
    .io_memoryStage_inst0_inst_info_fusel(MemoryUnit_io_memoryStage_inst0_inst_info_fusel),
    .io_memoryStage_inst0_inst_info_op(MemoryUnit_io_memoryStage_inst0_inst_info_op),
    .io_memoryStage_inst0_inst_info_reg_wen(MemoryUnit_io_memoryStage_inst0_inst_info_reg_wen),
    .io_memoryStage_inst0_inst_info_reg_waddr(MemoryUnit_io_memoryStage_inst0_inst_info_reg_waddr),
    .io_memoryStage_inst0_inst_info_inst(MemoryUnit_io_memoryStage_inst0_inst_info_inst),
    .io_memoryStage_inst0_rd_info_wdata(MemoryUnit_io_memoryStage_inst0_rd_info_wdata),
    .io_memoryStage_inst0_ex_flush_req(MemoryUnit_io_memoryStage_inst0_ex_flush_req),
    .io_memoryStage_inst0_ex_eret(MemoryUnit_io_memoryStage_inst0_ex_eret),
    .io_memoryStage_inst0_ex_badvaddr(MemoryUnit_io_memoryStage_inst0_ex_badvaddr),
    .io_memoryStage_inst0_ex_bd(MemoryUnit_io_memoryStage_inst0_ex_bd),
    .io_memoryStage_inst0_ex_excode(MemoryUnit_io_memoryStage_inst0_ex_excode),
    .io_memoryStage_inst0_cp0_cp0_count(MemoryUnit_io_memoryStage_inst0_cp0_cp0_count),
    .io_memoryStage_inst0_cp0_cp0_random(MemoryUnit_io_memoryStage_inst0_cp0_cp0_random),
    .io_memoryStage_inst0_cp0_cp0_cause(MemoryUnit_io_memoryStage_inst0_cp0_cp0_cause),
    .io_memoryStage_inst0_mem_en(MemoryUnit_io_memoryStage_inst0_mem_en),
    .io_memoryStage_inst0_mem_inst_info_op(MemoryUnit_io_memoryStage_inst0_mem_inst_info_op),
    .io_memoryStage_inst0_mem_addr(MemoryUnit_io_memoryStage_inst0_mem_addr),
    .io_memoryStage_inst0_mem_wdata(MemoryUnit_io_memoryStage_inst0_mem_wdata),
    .io_memoryStage_inst0_mem_sel_0(MemoryUnit_io_memoryStage_inst0_mem_sel_0),
    .io_memoryStage_inst0_mem_sel_1(MemoryUnit_io_memoryStage_inst0_mem_sel_1),
    .io_memoryStage_inst1_pc(MemoryUnit_io_memoryStage_inst1_pc),
    .io_memoryStage_inst1_inst_info_fusel(MemoryUnit_io_memoryStage_inst1_inst_info_fusel),
    .io_memoryStage_inst1_inst_info_reg_wen(MemoryUnit_io_memoryStage_inst1_inst_info_reg_wen),
    .io_memoryStage_inst1_inst_info_reg_waddr(MemoryUnit_io_memoryStage_inst1_inst_info_reg_waddr),
    .io_memoryStage_inst1_rd_info_wdata(MemoryUnit_io_memoryStage_inst1_rd_info_wdata),
    .io_memoryStage_inst1_ex_flush_req(MemoryUnit_io_memoryStage_inst1_ex_flush_req),
    .io_memoryStage_inst1_ex_eret(MemoryUnit_io_memoryStage_inst1_ex_eret),
    .io_memoryStage_inst1_ex_badvaddr(MemoryUnit_io_memoryStage_inst1_ex_badvaddr),
    .io_memoryStage_inst1_ex_bd(MemoryUnit_io_memoryStage_inst1_ex_bd),
    .io_memoryStage_inst1_ex_excode(MemoryUnit_io_memoryStage_inst1_ex_excode),
    .io_fetchUnit_flush(MemoryUnit_io_fetchUnit_flush),
    .io_fetchUnit_flush_pc(MemoryUnit_io_fetchUnit_flush_pc),
    .io_fetchUnit_ex_flush(MemoryUnit_io_fetchUnit_ex_flush),
    .io_fetchUnit_ex_flush_pc(MemoryUnit_io_fetchUnit_ex_flush_pc),
    .io_decoderUnit_0_wen(MemoryUnit_io_decoderUnit_0_wen),
    .io_decoderUnit_0_waddr(MemoryUnit_io_decoderUnit_0_waddr),
    .io_decoderUnit_0_wdata(MemoryUnit_io_decoderUnit_0_wdata),
    .io_decoderUnit_1_wen(MemoryUnit_io_decoderUnit_1_wen),
    .io_decoderUnit_1_waddr(MemoryUnit_io_decoderUnit_1_waddr),
    .io_decoderUnit_1_wdata(MemoryUnit_io_decoderUnit_1_wdata),
    .io_cp0_in_inst_0_pc(MemoryUnit_io_cp0_in_inst_0_pc),
    .io_cp0_in_inst_0_ex_flush_req(MemoryUnit_io_cp0_in_inst_0_ex_flush_req),
    .io_cp0_in_inst_0_ex_tlb_refill(MemoryUnit_io_cp0_in_inst_0_ex_tlb_refill),
    .io_cp0_in_inst_0_ex_eret(MemoryUnit_io_cp0_in_inst_0_ex_eret),
    .io_cp0_in_inst_0_ex_badvaddr(MemoryUnit_io_cp0_in_inst_0_ex_badvaddr),
    .io_cp0_in_inst_0_ex_bd(MemoryUnit_io_cp0_in_inst_0_ex_bd),
    .io_cp0_in_inst_0_ex_excode(MemoryUnit_io_cp0_in_inst_0_ex_excode),
    .io_cp0_in_inst_1_pc(MemoryUnit_io_cp0_in_inst_1_pc),
    .io_cp0_in_inst_1_ex_flush_req(MemoryUnit_io_cp0_in_inst_1_ex_flush_req),
    .io_cp0_in_inst_1_ex_tlb_refill(MemoryUnit_io_cp0_in_inst_1_ex_tlb_refill),
    .io_cp0_in_inst_1_ex_eret(MemoryUnit_io_cp0_in_inst_1_ex_eret),
    .io_cp0_in_inst_1_ex_badvaddr(MemoryUnit_io_cp0_in_inst_1_ex_badvaddr),
    .io_cp0_in_inst_1_ex_bd(MemoryUnit_io_cp0_in_inst_1_ex_bd),
    .io_cp0_in_inst_1_ex_excode(MemoryUnit_io_cp0_in_inst_1_ex_excode),
    .io_cp0_out_flush(MemoryUnit_io_cp0_out_flush),
    .io_cp0_out_flush_pc(MemoryUnit_io_cp0_out_flush_pc),
    .io_writeBackStage_inst0_pc(MemoryUnit_io_writeBackStage_inst0_pc),
    .io_writeBackStage_inst0_inst_info_fusel(MemoryUnit_io_writeBackStage_inst0_inst_info_fusel),
    .io_writeBackStage_inst0_inst_info_op(MemoryUnit_io_writeBackStage_inst0_inst_info_op),
    .io_writeBackStage_inst0_inst_info_reg_wen(MemoryUnit_io_writeBackStage_inst0_inst_info_reg_wen),
    .io_writeBackStage_inst0_inst_info_reg_waddr(MemoryUnit_io_writeBackStage_inst0_inst_info_reg_waddr),
    .io_writeBackStage_inst0_inst_info_inst(MemoryUnit_io_writeBackStage_inst0_inst_info_inst),
    .io_writeBackStage_inst0_rd_info_wdata(MemoryUnit_io_writeBackStage_inst0_rd_info_wdata),
    .io_writeBackStage_inst0_ex_flush_req(MemoryUnit_io_writeBackStage_inst0_ex_flush_req),
    .io_writeBackStage_inst0_ex_tlb_refill(MemoryUnit_io_writeBackStage_inst0_ex_tlb_refill),
    .io_writeBackStage_inst0_ex_eret(MemoryUnit_io_writeBackStage_inst0_ex_eret),
    .io_writeBackStage_inst0_ex_badvaddr(MemoryUnit_io_writeBackStage_inst0_ex_badvaddr),
    .io_writeBackStage_inst0_ex_bd(MemoryUnit_io_writeBackStage_inst0_ex_bd),
    .io_writeBackStage_inst0_ex_excode(MemoryUnit_io_writeBackStage_inst0_ex_excode),
    .io_writeBackStage_inst0_cp0_cp0_count(MemoryUnit_io_writeBackStage_inst0_cp0_cp0_count),
    .io_writeBackStage_inst0_cp0_cp0_random(MemoryUnit_io_writeBackStage_inst0_cp0_cp0_random),
    .io_writeBackStage_inst0_cp0_cp0_cause(MemoryUnit_io_writeBackStage_inst0_cp0_cp0_cause),
    .io_writeBackStage_inst1_pc(MemoryUnit_io_writeBackStage_inst1_pc),
    .io_writeBackStage_inst1_inst_info_fusel(MemoryUnit_io_writeBackStage_inst1_inst_info_fusel),
    .io_writeBackStage_inst1_inst_info_reg_wen(MemoryUnit_io_writeBackStage_inst1_inst_info_reg_wen),
    .io_writeBackStage_inst1_inst_info_reg_waddr(MemoryUnit_io_writeBackStage_inst1_inst_info_reg_waddr),
    .io_writeBackStage_inst1_rd_info_wdata(MemoryUnit_io_writeBackStage_inst1_rd_info_wdata),
    .io_writeBackStage_inst1_ex_flush_req(MemoryUnit_io_writeBackStage_inst1_ex_flush_req),
    .io_writeBackStage_inst1_ex_tlb_refill(MemoryUnit_io_writeBackStage_inst1_ex_tlb_refill),
    .io_writeBackStage_inst1_ex_eret(MemoryUnit_io_writeBackStage_inst1_ex_eret),
    .io_writeBackStage_inst1_ex_badvaddr(MemoryUnit_io_writeBackStage_inst1_ex_badvaddr),
    .io_writeBackStage_inst1_ex_bd(MemoryUnit_io_writeBackStage_inst1_ex_bd),
    .io_writeBackStage_inst1_ex_excode(MemoryUnit_io_writeBackStage_inst1_ex_excode),
    .io_dataMemory_in_tlb_invalid(MemoryUnit_io_dataMemory_in_tlb_invalid),
    .io_dataMemory_in_tlb_refill(MemoryUnit_io_dataMemory_in_tlb_refill),
    .io_dataMemory_in_tlb_modify(MemoryUnit_io_dataMemory_in_tlb_modify),
    .io_dataMemory_in_rdata(MemoryUnit_io_dataMemory_in_rdata),
    .io_dataMemory_out_en(MemoryUnit_io_dataMemory_out_en),
    .io_dataMemory_out_rlen(MemoryUnit_io_dataMemory_out_rlen),
    .io_dataMemory_out_wen(MemoryUnit_io_dataMemory_out_wen),
    .io_dataMemory_out_wdata(MemoryUnit_io_dataMemory_out_wdata)
  );
  WriteBackStage WriteBackStage ( // @[Core.scala 35:30]
    .clock(WriteBackStage_clock),
    .reset(WriteBackStage_reset),
    .io_ctrl_allow_to_go(WriteBackStage_io_ctrl_allow_to_go),
    .io_memoryUnit_inst0_pc(WriteBackStage_io_memoryUnit_inst0_pc),
    .io_memoryUnit_inst0_inst_info_reg_wen(WriteBackStage_io_memoryUnit_inst0_inst_info_reg_wen),
    .io_memoryUnit_inst0_inst_info_reg_waddr(WriteBackStage_io_memoryUnit_inst0_inst_info_reg_waddr),
    .io_memoryUnit_inst0_rd_info_wdata(WriteBackStage_io_memoryUnit_inst0_rd_info_wdata),
    .io_memoryUnit_inst0_ex_flush_req(WriteBackStage_io_memoryUnit_inst0_ex_flush_req),
    .io_memoryUnit_inst0_ex_excode(WriteBackStage_io_memoryUnit_inst0_ex_excode),
    .io_memoryUnit_inst0_cp0_cp0_count(WriteBackStage_io_memoryUnit_inst0_cp0_cp0_count),
    .io_memoryUnit_inst0_cp0_cp0_random(WriteBackStage_io_memoryUnit_inst0_cp0_cp0_random),
    .io_memoryUnit_inst0_cp0_cp0_cause(WriteBackStage_io_memoryUnit_inst0_cp0_cp0_cause),
    .io_memoryUnit_inst1_pc(WriteBackStage_io_memoryUnit_inst1_pc),
    .io_memoryUnit_inst1_inst_info_reg_wen(WriteBackStage_io_memoryUnit_inst1_inst_info_reg_wen),
    .io_memoryUnit_inst1_inst_info_reg_waddr(WriteBackStage_io_memoryUnit_inst1_inst_info_reg_waddr),
    .io_memoryUnit_inst1_rd_info_wdata(WriteBackStage_io_memoryUnit_inst1_rd_info_wdata),
    .io_memoryUnit_inst1_ex_flush_req(WriteBackStage_io_memoryUnit_inst1_ex_flush_req),
    .io_writeBackUnit_inst0_pc(WriteBackStage_io_writeBackUnit_inst0_pc),
    .io_writeBackUnit_inst0_inst_info_reg_wen(WriteBackStage_io_writeBackUnit_inst0_inst_info_reg_wen),
    .io_writeBackUnit_inst0_inst_info_reg_waddr(WriteBackStage_io_writeBackUnit_inst0_inst_info_reg_waddr),
    .io_writeBackUnit_inst0_rd_info_wdata(WriteBackStage_io_writeBackUnit_inst0_rd_info_wdata),
    .io_writeBackUnit_inst0_ex_flush_req(WriteBackStage_io_writeBackUnit_inst0_ex_flush_req),
    .io_writeBackUnit_inst0_ex_excode(WriteBackStage_io_writeBackUnit_inst0_ex_excode),
    .io_writeBackUnit_inst0_cp0_cp0_count(WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_count),
    .io_writeBackUnit_inst0_cp0_cp0_random(WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_random),
    .io_writeBackUnit_inst0_cp0_cp0_cause(WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_cause),
    .io_writeBackUnit_inst1_pc(WriteBackStage_io_writeBackUnit_inst1_pc),
    .io_writeBackUnit_inst1_inst_info_reg_wen(WriteBackStage_io_writeBackUnit_inst1_inst_info_reg_wen),
    .io_writeBackUnit_inst1_inst_info_reg_waddr(WriteBackStage_io_writeBackUnit_inst1_inst_info_reg_waddr),
    .io_writeBackUnit_inst1_rd_info_wdata(WriteBackStage_io_writeBackUnit_inst1_rd_info_wdata),
    .io_writeBackUnit_inst1_ex_flush_req(WriteBackStage_io_writeBackUnit_inst1_ex_flush_req)
  );
  WriteBackUnit WriteBackUnit ( // @[Core.scala 36:30]
    .clock(WriteBackUnit_clock),
    .reset(WriteBackUnit_reset),
    .io_ctrl_allow_to_go(WriteBackUnit_io_ctrl_allow_to_go),
    .io_writeBackStage_inst0_pc(WriteBackUnit_io_writeBackStage_inst0_pc),
    .io_writeBackStage_inst0_inst_info_reg_wen(WriteBackUnit_io_writeBackStage_inst0_inst_info_reg_wen),
    .io_writeBackStage_inst0_inst_info_reg_waddr(WriteBackUnit_io_writeBackStage_inst0_inst_info_reg_waddr),
    .io_writeBackStage_inst0_rd_info_wdata(WriteBackUnit_io_writeBackStage_inst0_rd_info_wdata),
    .io_writeBackStage_inst0_ex_flush_req(WriteBackUnit_io_writeBackStage_inst0_ex_flush_req),
    .io_writeBackStage_inst0_ex_excode(WriteBackUnit_io_writeBackStage_inst0_ex_excode),
    .io_writeBackStage_inst0_cp0_cp0_count(WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_count),
    .io_writeBackStage_inst0_cp0_cp0_random(WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_random),
    .io_writeBackStage_inst0_cp0_cp0_cause(WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_cause),
    .io_writeBackStage_inst1_pc(WriteBackUnit_io_writeBackStage_inst1_pc),
    .io_writeBackStage_inst1_inst_info_reg_wen(WriteBackUnit_io_writeBackStage_inst1_inst_info_reg_wen),
    .io_writeBackStage_inst1_inst_info_reg_waddr(WriteBackUnit_io_writeBackStage_inst1_inst_info_reg_waddr),
    .io_writeBackStage_inst1_rd_info_wdata(WriteBackUnit_io_writeBackStage_inst1_rd_info_wdata),
    .io_writeBackStage_inst1_ex_flush_req(WriteBackUnit_io_writeBackStage_inst1_ex_flush_req),
    .io_regfile_0_wen(WriteBackUnit_io_regfile_0_wen),
    .io_regfile_0_waddr(WriteBackUnit_io_regfile_0_waddr),
    .io_regfile_0_wdata(WriteBackUnit_io_regfile_0_wdata),
    .io_regfile_1_wen(WriteBackUnit_io_regfile_1_wen),
    .io_regfile_1_waddr(WriteBackUnit_io_regfile_1_waddr),
    .io_regfile_1_wdata(WriteBackUnit_io_regfile_1_wdata),
    .io_debug_wb_pc(WriteBackUnit_io_debug_wb_pc),
    .io_debug_wb_rf_wen(WriteBackUnit_io_debug_wb_rf_wen),
    .io_debug_wb_rf_wnum(WriteBackUnit_io_debug_wb_rf_wnum),
    .io_debug_wb_rf_wdata(WriteBackUnit_io_debug_wb_rf_wdata),
    .io_debug_cp0_count(WriteBackUnit_io_debug_cp0_count),
    .io_debug_cp0_random(WriteBackUnit_io_debug_cp0_random),
    .io_debug_cp0_cause(WriteBackUnit_io_debug_cp0_cause),
    .io_debug_int(WriteBackUnit_io_debug_int),
    .io_debug_commit(WriteBackUnit_io_debug_commit)
  );
  assign io_inst_req = ~(reset | InstBuffer_io_full); // @[Core.scala 181:29]
  assign io_inst_addr_0 = FetchStage_io_iCache_pc; // @[Core.scala 53:31]
  assign io_inst_addr_1 = FetchStage_io_iCache_pc_next; // @[Core.scala 54:31]
  assign io_inst_cpu_stall = ~Ctrl_io_fetchUnit_allow_to_go; // @[Core.scala 182:29]
  assign io_inst_tlb2_found = Cp0_io_tlb_0_found; // @[Core.scala 131:22]
  assign io_inst_tlb2_entry_pfn_0 = Cp0_io_tlb_0_info_pfn_0; // @[Core.scala 133:22]
  assign io_inst_tlb2_entry_pfn_1 = Cp0_io_tlb_0_info_pfn_1; // @[Core.scala 133:22]
  assign io_inst_tlb2_entry_c_0 = Cp0_io_tlb_0_info_c_0; // @[Core.scala 133:22]
  assign io_inst_tlb2_entry_c_1 = Cp0_io_tlb_0_info_c_1; // @[Core.scala 133:22]
  assign io_inst_tlb2_entry_v_0 = Cp0_io_tlb_0_info_v_0; // @[Core.scala 133:22]
  assign io_inst_tlb2_entry_v_1 = Cp0_io_tlb_0_info_v_1; // @[Core.scala 133:22]
  assign io_inst_fence_value = ~ExecuteUnit_io_memoryStage_inst0_inst_info_inst[16] &
    ExecuteUnit_io_memoryStage_inst0_inst_info_op == 7'h4c; // @[Core.scala 173:86]
  assign io_inst_fence_addr = ExecuteUnit_io_memoryStage_inst0_rd_info_wdata; // @[Core.scala 174:26]
  assign io_inst_fence_tlb = 7'h12 == ExecuteUnit_io_executeStage_inst0_inst_info_op | 7'h4a ==
    ExecuteUnit_io_executeStage_inst0_inst_info_op | 7'h4b == ExecuteUnit_io_executeStage_inst0_inst_info_op; // @[Core.scala 177:77]
  assign io_data_stallM = ~Ctrl_io_memoryUnit_allow_to_go; // @[Core.scala 183:29]
  assign io_data_E_mem_va = ExecuteUnit_io_memoryStage_inst0_mem_addr; // @[Core.scala 179:26]
  assign io_data_M_mem_va = MemoryUnit_io_memoryStage_inst0_mem_addr; // @[Core.scala 180:26]
  assign io_data_M_fence_addr = MemoryUnit_io_writeBackStage_inst0_rd_info_wdata; // @[Core.scala 176:26]
  assign io_data_M_fence_d = MemoryUnit_io_writeBackStage_inst0_inst_info_inst[16] &
    MemoryUnit_io_writeBackStage_inst0_inst_info_op == 7'h4c; // @[Core.scala 175:88]
  assign io_data_M_mem_en = MemoryUnit_io_dataMemory_out_en; // @[Core.scala 148:40]
  assign io_data_M_mem_write = |MemoryUnit_io_dataMemory_out_wen; // @[Core.scala 149:73]
  assign io_data_M_wmask = MemoryUnit_io_dataMemory_out_wen; // @[Core.scala 151:40]
  assign io_data_M_mem_size = MemoryUnit_io_dataMemory_out_rlen; // @[Core.scala 150:40]
  assign io_data_M_wdata = MemoryUnit_io_dataMemory_out_wdata; // @[Core.scala 152:40]
  assign io_data_tlb_found = Cp0_io_tlb_1_found; // @[Core.scala 132:22]
  assign io_data_tlb_entry_pfn_0 = Cp0_io_tlb_1_info_pfn_0; // @[Core.scala 134:22]
  assign io_data_tlb_entry_pfn_1 = Cp0_io_tlb_1_info_pfn_1; // @[Core.scala 134:22]
  assign io_data_tlb_entry_c_0 = Cp0_io_tlb_1_info_c_0; // @[Core.scala 134:22]
  assign io_data_tlb_entry_c_1 = Cp0_io_tlb_1_info_c_1; // @[Core.scala 134:22]
  assign io_data_tlb_entry_d_0 = Cp0_io_tlb_1_info_d_0; // @[Core.scala 134:22]
  assign io_data_tlb_entry_d_1 = Cp0_io_tlb_1_info_d_1; // @[Core.scala 134:22]
  assign io_data_tlb_entry_v_0 = Cp0_io_tlb_1_info_v_0; // @[Core.scala 134:22]
  assign io_data_tlb_entry_v_1 = Cp0_io_tlb_1_info_v_1; // @[Core.scala 134:22]
  assign io_data_fence_tlb = 7'h12 == MemoryUnit_io_memoryStage_inst0_inst_info_op | 7'h4a ==
    MemoryUnit_io_memoryStage_inst0_inst_info_op | 7'h4b == MemoryUnit_io_memoryStage_inst0_inst_info_op; // @[Core.scala 178:77]
  assign io_debug_wb_pc = WriteBackUnit_io_debug_wb_pc; // @[Core.scala 165:24]
  assign io_debug_wb_rf_wen = WriteBackUnit_io_debug_wb_rf_wen; // @[Core.scala 166:24]
  assign io_debug_wb_rf_wnum = WriteBackUnit_io_debug_wb_rf_wnum; // @[Core.scala 167:24]
  assign io_debug_wb_rf_wdata = WriteBackUnit_io_debug_wb_rf_wdata; // @[Core.scala 168:24]
  assign io_debug_cp0_count = WriteBackUnit_io_debug_cp0_count; // @[Core.scala 169:24]
  assign io_debug_cp0_random = WriteBackUnit_io_debug_cp0_random; // @[Core.scala 170:24]
  assign io_debug_cp0_cause = WriteBackUnit_io_debug_cp0_cause; // @[Core.scala 171:24]
  assign io_debug_int = WriteBackUnit_io_debug_int; // @[Core.scala 164:24]
  assign io_debug_commit = WriteBackUnit_io_debug_commit; // @[Core.scala 163:24]
  assign Ctrl_io_cacheCtrl_iCache_stall = io_inst_icache_stall; // @[Core.scala 42:31]
  assign Ctrl_io_cacheCtrl_dCache_stall = io_data_dstall; // @[Core.scala 43:31]
  assign Ctrl_io_decoderUnit_inst0_src1_ren = DecoderUnit_io_ctrl_inst0_src1_ren; // @[Core.scala 38:20]
  assign Ctrl_io_decoderUnit_inst0_src1_raddr = DecoderUnit_io_ctrl_inst0_src1_raddr; // @[Core.scala 38:20]
  assign Ctrl_io_decoderUnit_inst0_src2_ren = DecoderUnit_io_ctrl_inst0_src2_ren; // @[Core.scala 38:20]
  assign Ctrl_io_decoderUnit_inst0_src2_raddr = DecoderUnit_io_ctrl_inst0_src2_raddr; // @[Core.scala 38:20]
  assign Ctrl_io_decoderUnit_branch_flag = DecoderUnit_io_ctrl_branch_flag; // @[Core.scala 38:20]
  assign Ctrl_io_executeUnit_inst_0_mem_ren = ExecuteUnit_io_ctrl_inst_0_mem_ren; // @[Core.scala 39:20]
  assign Ctrl_io_executeUnit_inst_0_reg_waddr = ExecuteUnit_io_ctrl_inst_0_reg_waddr; // @[Core.scala 39:20]
  assign Ctrl_io_executeUnit_inst_1_mem_ren = ExecuteUnit_io_ctrl_inst_1_mem_ren; // @[Core.scala 39:20]
  assign Ctrl_io_executeUnit_inst_1_reg_waddr = ExecuteUnit_io_ctrl_inst_1_reg_waddr; // @[Core.scala 39:20]
  assign Ctrl_io_executeUnit_fu_stall = ExecuteUnit_io_ctrl_fu_stall; // @[Core.scala 39:20]
  assign Ctrl_io_executeUnit_branch_flag = ExecuteUnit_io_ctrl_branch_flag; // @[Core.scala 39:20]
  assign Ctrl_io_memoryUnit_flush_req = MemoryUnit_io_ctrl_flush_req; // @[Core.scala 40:19]
  assign FetchStage_clock = clock;
  assign FetchStage_reset = reset;
  assign FetchStage_io_memory_ex = MemoryUnit_io_fetchUnit_ex_flush; // @[Core.scala 45:29]
  assign FetchStage_io_memory_ex_pc = MemoryUnit_io_fetchUnit_ex_flush_pc; // @[Core.scala 46:29]
  assign FetchStage_io_memory_flush = MemoryUnit_io_fetchUnit_flush; // @[Core.scala 47:29]
  assign FetchStage_io_memory_flush_pc = MemoryUnit_io_fetchUnit_flush_pc; // @[Core.scala 48:29]
  assign FetchStage_io_decoder_branch = DecoderUnit_io_fetchUnit_branch; // @[Core.scala 50:21]
  assign FetchStage_io_decoder_target = DecoderUnit_io_fetchUnit_target; // @[Core.scala 50:21]
  assign FetchStage_io_execute_branch = ExecuteUnit_io_fetchStage_branch; // @[Core.scala 49:21]
  assign FetchStage_io_execute_target = ExecuteUnit_io_fetchStage_target; // @[Core.scala 49:21]
  assign FetchStage_io_instBuffer_full = InstBuffer_io_full; // @[Core.scala 51:31]
  assign FetchStage_io_iCache_inst_valid_0 = io_inst_inst_valid_0; // @[Core.scala 52:31]
  assign FetchStage_io_iCache_inst_valid_1 = io_inst_inst_valid_1; // @[Core.scala 52:31]
  assign BPU_clock = clock;
  assign BPU_reset = reset;
  assign BPU_io_instrD = DecoderUnit_io_bpu_decoded_inst0_inst; // @[Core.scala 57:36]
  assign BPU_io_enaD = Ctrl_io_decoderUnit_allow_to_go; // @[Core.scala 56:36]
  assign BPU_io_pcD = DecoderUnit_io_bpu_pc; // @[Core.scala 58:36]
  assign BPU_io_pc_plus4D = DecoderUnit_io_bpu_pc + 32'h4; // @[Core.scala 59:58]
  assign BPU_io_pcE = ExecuteUnit_io_bpu_pc; // @[Core.scala 60:36]
  assign BPU_io_branchE = ExecuteUnit_io_bpu_inst0_is_branch; // @[Core.scala 61:36]
  assign BPU_io_actual_takeE = ExecuteUnit_io_bpu_branch_flag; // @[Core.scala 62:36]
  assign InstBuffer_clock = clock;
  assign InstBuffer_reset = reset;
  assign InstBuffer_io_fifo_rst = reset | Ctrl_io_decoderUnit_do_flush; // @[Core.scala 67:47]
  assign InstBuffer_io_flush_delay_slot = Ctrl_io_instBuffer_delay_slot_do_flush; // @[Core.scala 68:31]
  assign InstBuffer_io_delay_sel_rst = Ctrl_io_executeUnit_branch_flag ? _T_5 : _T_7; // @[Core.scala 72:34]
  assign InstBuffer_io_D_delay_rst = Ctrl_io_decoderUnit_branch_flag; // @[Core.scala 81:26]
  assign InstBuffer_io_E_delay_rst = Ctrl_io_executeUnit_branch_flag; // @[Core.scala 82:26]
  assign InstBuffer_io_i_stall = io_inst_icache_stall; // @[Core.scala 70:31]
  assign InstBuffer_io_master_is_branch = DecoderUnit_io_instBuffer_inst0_is_jb; // @[Core.scala 71:31]
  assign InstBuffer_io_read_en_0 = DecoderUnit_io_instBuffer_inst_0_ready; // @[Core.scala 84:53]
  assign InstBuffer_io_read_en_1 = DecoderUnit_io_instBuffer_inst_1_ready; // @[Core.scala 84:53]
  assign InstBuffer_io_write_en_0 = io_inst_inst_valid_0; // @[Core.scala 91:32]
  assign InstBuffer_io_write_en_1 = io_inst_inst_valid_1; // @[Core.scala 91:32]
  assign InstBuffer_io_write_0_tlb_invalid = io_inst_tlb1_invalid; // @[Core.scala 94:35]
  assign InstBuffer_io_write_0_data = io_inst_inst_0; // @[Core.scala 98:35]
  assign InstBuffer_io_write_0_addr = io_inst_addr_0; // @[Core.scala 96:35]
  assign InstBuffer_io_write_1_tlb_invalid = io_inst_tlb1_invalid; // @[Core.scala 95:35]
  assign InstBuffer_io_write_1_data = io_inst_inst_1; // @[Core.scala 99:35]
  assign InstBuffer_io_write_1_addr = io_inst_addr_0 + 32'h4; // @[Core.scala 97:54]
  assign DecoderUnit_io_instBuffer_inst_0_bits_pc = InstBuffer_io_read_0_addr; // @[Core.scala 88:53]
  assign DecoderUnit_io_instBuffer_inst_0_bits_inst = InstBuffer_io_read_0_data; // @[Core.scala 89:53]
  assign DecoderUnit_io_instBuffer_inst_0_bits_tlb_invalid = InstBuffer_io_read_0_tlb_invalid; // @[Core.scala 87:53]
  assign DecoderUnit_io_instBuffer_inst_1_bits_pc = InstBuffer_io_read_1_addr; // @[Core.scala 88:53]
  assign DecoderUnit_io_instBuffer_inst_1_bits_inst = InstBuffer_io_read_1_data; // @[Core.scala 89:53]
  assign DecoderUnit_io_instBuffer_inst_1_bits_tlb_invalid = InstBuffer_io_read_1_tlb_invalid; // @[Core.scala 87:53]
  assign DecoderUnit_io_instBuffer_info_inst0_is_in_delayslot = InstBuffer_io_master_is_in_delayslot_o; // @[Core.scala 103:53]
  assign DecoderUnit_io_instBuffer_info_empty = InstBuffer_io_empty; // @[Core.scala 101:53]
  assign DecoderUnit_io_instBuffer_info_almost_empty = InstBuffer_io_almost_empty; // @[Core.scala 102:53]
  assign DecoderUnit_io_regfile_0_src1_rdata = ARegFile_io_read_0_src1_rdata; // @[Core.scala 104:23]
  assign DecoderUnit_io_regfile_0_src2_rdata = ARegFile_io_read_0_src2_rdata; // @[Core.scala 104:23]
  assign DecoderUnit_io_regfile_1_src1_rdata = ARegFile_io_read_1_src1_rdata; // @[Core.scala 104:23]
  assign DecoderUnit_io_regfile_1_src2_rdata = ARegFile_io_read_1_src2_rdata; // @[Core.scala 104:23]
  assign DecoderUnit_io_forward_0_exe_wen = ExecuteUnit_io_decoderUnit_forward_0_exe_wen; // @[Core.scala 106:40]
  assign DecoderUnit_io_forward_0_exe_waddr = ExecuteUnit_io_decoderUnit_forward_0_exe_waddr; // @[Core.scala 106:40]
  assign DecoderUnit_io_forward_0_exe_wdata = ExecuteUnit_io_decoderUnit_forward_0_exe_wdata; // @[Core.scala 106:40]
  assign DecoderUnit_io_forward_0_exe_mem_ren = ExecuteUnit_io_decoderUnit_forward_0_exe_mem_ren; // @[Core.scala 107:40]
  assign DecoderUnit_io_forward_0_mem_wen = MemoryUnit_io_decoderUnit_0_wen; // @[Core.scala 108:40]
  assign DecoderUnit_io_forward_0_mem_waddr = MemoryUnit_io_decoderUnit_0_waddr; // @[Core.scala 108:40]
  assign DecoderUnit_io_forward_0_mem_wdata = MemoryUnit_io_decoderUnit_0_wdata; // @[Core.scala 108:40]
  assign DecoderUnit_io_forward_1_exe_wen = ExecuteUnit_io_decoderUnit_forward_1_exe_wen; // @[Core.scala 106:40]
  assign DecoderUnit_io_forward_1_exe_waddr = ExecuteUnit_io_decoderUnit_forward_1_exe_waddr; // @[Core.scala 106:40]
  assign DecoderUnit_io_forward_1_exe_wdata = ExecuteUnit_io_decoderUnit_forward_1_exe_wdata; // @[Core.scala 106:40]
  assign DecoderUnit_io_forward_1_exe_mem_ren = ExecuteUnit_io_decoderUnit_forward_1_exe_mem_ren; // @[Core.scala 107:40]
  assign DecoderUnit_io_forward_1_mem_wen = MemoryUnit_io_decoderUnit_1_wen; // @[Core.scala 108:40]
  assign DecoderUnit_io_forward_1_mem_waddr = MemoryUnit_io_decoderUnit_1_waddr; // @[Core.scala 108:40]
  assign DecoderUnit_io_forward_1_mem_wdata = MemoryUnit_io_decoderUnit_1_wdata; // @[Core.scala 108:40]
  assign DecoderUnit_io_cp0_access_allowed = Cp0_io_decoderUnit_access_allowed; // @[Core.scala 110:19]
  assign DecoderUnit_io_cp0_kernel_mode = Cp0_io_decoderUnit_kernel_mode; // @[Core.scala 110:19]
  assign DecoderUnit_io_cp0_intterupt_allowed = Cp0_io_decoderUnit_intterupt_allowed; // @[Core.scala 110:19]
  assign DecoderUnit_io_cp0_cause_ip = Cp0_io_decoderUnit_cause_ip; // @[Core.scala 110:19]
  assign DecoderUnit_io_cp0_status_im = Cp0_io_decoderUnit_status_im; // @[Core.scala 110:19]
  assign DecoderUnit_io_bpu_inst_is_branch = BPU_io_branchD; // @[Core.scala 63:36]
  assign DecoderUnit_io_bpu_pred_branch_flag = BPU_io_pred_takeD; // @[Core.scala 64:36]
  assign DecoderUnit_io_bpu_branch_target = BPU_io_branch_targetD; // @[Core.scala 65:36]
  assign DecoderUnit_io_ctrl_allow_to_go = Ctrl_io_decoderUnit_allow_to_go; // @[Core.scala 38:20]
  assign ARegFile_clock = clock;
  assign ARegFile_reset = reset;
  assign ARegFile_io_read_0_src1_raddr = DecoderUnit_io_regfile_0_src1_raddr; // @[Core.scala 104:23]
  assign ARegFile_io_read_0_src2_raddr = DecoderUnit_io_regfile_0_src2_raddr; // @[Core.scala 104:23]
  assign ARegFile_io_read_1_src1_raddr = DecoderUnit_io_regfile_1_src1_raddr; // @[Core.scala 104:23]
  assign ARegFile_io_read_1_src2_raddr = DecoderUnit_io_regfile_1_src2_raddr; // @[Core.scala 104:23]
  assign ARegFile_io_write_0_wen = WriteBackUnit_io_regfile_0_wen; // @[Core.scala 161:17]
  assign ARegFile_io_write_0_waddr = WriteBackUnit_io_regfile_0_waddr; // @[Core.scala 161:17]
  assign ARegFile_io_write_0_wdata = WriteBackUnit_io_regfile_0_wdata; // @[Core.scala 161:17]
  assign ARegFile_io_write_1_wen = WriteBackUnit_io_regfile_1_wen; // @[Core.scala 161:17]
  assign ARegFile_io_write_1_waddr = WriteBackUnit_io_regfile_1_waddr; // @[Core.scala 161:17]
  assign ARegFile_io_write_1_wdata = WriteBackUnit_io_regfile_1_wdata; // @[Core.scala 161:17]
  assign ExecuteStage_clock = clock;
  assign ExecuteStage_reset = reset;
  assign ExecuteStage_io_ctrl_inst0_allow_to_go = Ctrl_io_executeUnit_allow_to_go; // @[Core.scala 119:39]
  assign ExecuteStage_io_ctrl_clear_0 = _T_14 | _T_16; // @[Core.scala 114:104]
  assign ExecuteStage_io_ctrl_clear_1 = _T_19 | _T_21; // @[Core.scala 117:79]
  assign ExecuteStage_io_decoderUnit_inst0_pc = DecoderUnit_io_executeStage_inst0_pc; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_inst_info_fusel = DecoderUnit_io_executeStage_inst0_inst_info_fusel; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_inst_info_op = DecoderUnit_io_executeStage_inst0_inst_info_op; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_inst_info_reg_wen = DecoderUnit_io_executeStage_inst0_inst_info_reg_wen; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_inst_info_reg_waddr = DecoderUnit_io_executeStage_inst0_inst_info_reg_waddr; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_inst_info_cp0_addr = DecoderUnit_io_executeStage_inst0_inst_info_cp0_addr; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_inst_info_inst = DecoderUnit_io_executeStage_inst0_inst_info_inst; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_src_info_src1_data = DecoderUnit_io_executeStage_inst0_src_info_src1_data; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_src_info_src2_data = DecoderUnit_io_executeStage_inst0_src_info_src2_data; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_ex_flush_req = DecoderUnit_io_executeStage_inst0_ex_flush_req; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_ex_eret = DecoderUnit_io_executeStage_inst0_ex_eret; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_ex_badvaddr = DecoderUnit_io_executeStage_inst0_ex_badvaddr; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_ex_bd = DecoderUnit_io_executeStage_inst0_ex_bd; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_ex_excode = DecoderUnit_io_executeStage_inst0_ex_excode; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_jb_info_jump_regiser_conflict =
    DecoderUnit_io_executeStage_inst0_jb_info_jump_regiser_conflict; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_jb_info_is_branch = DecoderUnit_io_executeStage_inst0_jb_info_is_branch; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_jb_info_pred_branch_flag =
    DecoderUnit_io_executeStage_inst0_jb_info_pred_branch_flag; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst0_jb_info_branch_target =
    DecoderUnit_io_executeStage_inst0_jb_info_branch_target; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_allow_to_go = DecoderUnit_io_executeStage_inst1_allow_to_go; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_pc = DecoderUnit_io_executeStage_inst1_pc; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_inst_info_fusel = DecoderUnit_io_executeStage_inst1_inst_info_fusel; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_inst_info_op = DecoderUnit_io_executeStage_inst1_inst_info_op; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_inst_info_reg_wen = DecoderUnit_io_executeStage_inst1_inst_info_reg_wen; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_inst_info_reg_waddr = DecoderUnit_io_executeStage_inst1_inst_info_reg_waddr; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_inst_info_inst = DecoderUnit_io_executeStage_inst1_inst_info_inst; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_src_info_src1_data = DecoderUnit_io_executeStage_inst1_src_info_src1_data; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_src_info_src2_data = DecoderUnit_io_executeStage_inst1_src_info_src2_data; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_ex_flush_req = DecoderUnit_io_executeStage_inst1_ex_flush_req; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_ex_eret = DecoderUnit_io_executeStage_inst1_ex_eret; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_ex_badvaddr = DecoderUnit_io_executeStage_inst1_ex_badvaddr; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_ex_bd = DecoderUnit_io_executeStage_inst1_ex_bd; // @[Core.scala 111:28]
  assign ExecuteStage_io_decoderUnit_inst1_ex_excode = DecoderUnit_io_executeStage_inst1_ex_excode; // @[Core.scala 111:28]
  assign ExecuteUnit_clock = clock;
  assign ExecuteUnit_reset = reset;
  assign ExecuteUnit_io_ctrl_allow_to_go = Ctrl_io_executeUnit_allow_to_go; // @[Core.scala 39:20]
  assign ExecuteUnit_io_ctrl_fu_allow_to_go = Ctrl_io_executeUnit_fu_allow_to_go; // @[Core.scala 39:20]
  assign ExecuteUnit_io_ctrl_fu_do_flush = Ctrl_io_executeUnit_fu_do_flush; // @[Core.scala 39:20]
  assign ExecuteUnit_io_executeStage_inst0_pc = ExecuteStage_io_executeUnit_inst0_pc; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_inst_info_fusel = ExecuteStage_io_executeUnit_inst0_inst_info_fusel; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_inst_info_op = ExecuteStage_io_executeUnit_inst0_inst_info_op; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_inst_info_reg_wen = ExecuteStage_io_executeUnit_inst0_inst_info_reg_wen; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_inst_info_reg_waddr = ExecuteStage_io_executeUnit_inst0_inst_info_reg_waddr; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_inst_info_cp0_addr = ExecuteStage_io_executeUnit_inst0_inst_info_cp0_addr; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_inst_info_inst = ExecuteStage_io_executeUnit_inst0_inst_info_inst; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_src_info_src1_data = ExecuteStage_io_executeUnit_inst0_src_info_src1_data; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_src_info_src2_data = ExecuteStage_io_executeUnit_inst0_src_info_src2_data; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_ex_flush_req = ExecuteStage_io_executeUnit_inst0_ex_flush_req; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_ex_eret = ExecuteStage_io_executeUnit_inst0_ex_eret; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_ex_badvaddr = ExecuteStage_io_executeUnit_inst0_ex_badvaddr; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_ex_bd = ExecuteStage_io_executeUnit_inst0_ex_bd; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_ex_excode = ExecuteStage_io_executeUnit_inst0_ex_excode; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_jb_info_jump_regiser_conflict =
    ExecuteStage_io_executeUnit_inst0_jb_info_jump_regiser_conflict; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_jb_info_is_branch = ExecuteStage_io_executeUnit_inst0_jb_info_is_branch; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_jb_info_pred_branch_flag =
    ExecuteStage_io_executeUnit_inst0_jb_info_pred_branch_flag; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst0_jb_info_branch_target =
    ExecuteStage_io_executeUnit_inst0_jb_info_branch_target; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_pc = ExecuteStage_io_executeUnit_inst1_pc; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_inst_info_fusel = ExecuteStage_io_executeUnit_inst1_inst_info_fusel; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_inst_info_op = ExecuteStage_io_executeUnit_inst1_inst_info_op; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_inst_info_reg_wen = ExecuteStage_io_executeUnit_inst1_inst_info_reg_wen; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_inst_info_reg_waddr = ExecuteStage_io_executeUnit_inst1_inst_info_reg_waddr; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_inst_info_inst = ExecuteStage_io_executeUnit_inst1_inst_info_inst; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_src_info_src1_data = ExecuteStage_io_executeUnit_inst1_src_info_src1_data; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_src_info_src2_data = ExecuteStage_io_executeUnit_inst1_src_info_src2_data; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_ex_flush_req = ExecuteStage_io_executeUnit_inst1_ex_flush_req; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_ex_eret = ExecuteStage_io_executeUnit_inst1_ex_eret; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_ex_badvaddr = ExecuteStage_io_executeUnit_inst1_ex_badvaddr; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_ex_bd = ExecuteStage_io_executeUnit_inst1_ex_bd; // @[Core.scala 122:28]
  assign ExecuteUnit_io_executeStage_inst1_ex_excode = ExecuteStage_io_executeUnit_inst1_ex_excode; // @[Core.scala 122:28]
  assign ExecuteUnit_io_cp0_out_cp0_rdata = Cp0_io_executeUnit_out_cp0_rdata; // @[Core.scala 123:19]
  assign ExecuteUnit_io_cp0_out_debug_cp0_count = Cp0_io_executeUnit_out_debug_cp0_count; // @[Core.scala 123:19]
  assign ExecuteUnit_io_cp0_out_debug_cp0_random = Cp0_io_executeUnit_out_debug_cp0_random; // @[Core.scala 123:19]
  assign ExecuteUnit_io_cp0_out_debug_cp0_cause = Cp0_io_executeUnit_out_debug_cp0_cause; // @[Core.scala 123:19]
  assign ExecuteUnit_io_decoderUnit_inst0_bd = DecoderUnit_io_executeStage_inst0_ex_bd; // @[Core.scala 121:36]
  assign Cp0_clock = clock;
  assign Cp0_reset = reset;
  assign Cp0_io_ext_int = io_ext_int; // @[Core.scala 130:22]
  assign Cp0_io_ctrl_exe_stall = ~Ctrl_io_executeUnit_allow_to_go; // @[Core.scala 126:25]
  assign Cp0_io_ctrl_mem_stall = ~Ctrl_io_memoryUnit_allow_to_go; // @[Core.scala 127:25]
  assign Cp0_io_executeUnit_in_inst_info_op = ExecuteUnit_io_cp0_in_inst_info_op; // @[Core.scala 123:19]
  assign Cp0_io_executeUnit_in_inst_info_cp0_addr = ExecuteUnit_io_cp0_in_inst_info_cp0_addr; // @[Core.scala 123:19]
  assign Cp0_io_executeUnit_in_mtc0_wdata = ExecuteUnit_io_cp0_in_mtc0_wdata; // @[Core.scala 123:19]
  assign Cp0_io_memoryUnit_in_inst_0_pc = MemoryUnit_io_cp0_in_inst_0_pc; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_0_ex_flush_req = MemoryUnit_io_cp0_in_inst_0_ex_flush_req; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_0_ex_tlb_refill = MemoryUnit_io_cp0_in_inst_0_ex_tlb_refill; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_0_ex_eret = MemoryUnit_io_cp0_in_inst_0_ex_eret; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_0_ex_badvaddr = MemoryUnit_io_cp0_in_inst_0_ex_badvaddr; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_0_ex_bd = MemoryUnit_io_cp0_in_inst_0_ex_bd; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_0_ex_excode = MemoryUnit_io_cp0_in_inst_0_ex_excode; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_1_pc = MemoryUnit_io_cp0_in_inst_1_pc; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_1_ex_flush_req = MemoryUnit_io_cp0_in_inst_1_ex_flush_req; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_1_ex_tlb_refill = MemoryUnit_io_cp0_in_inst_1_ex_tlb_refill; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_1_ex_eret = MemoryUnit_io_cp0_in_inst_1_ex_eret; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_1_ex_badvaddr = MemoryUnit_io_cp0_in_inst_1_ex_badvaddr; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_1_ex_bd = MemoryUnit_io_cp0_in_inst_1_ex_bd; // @[Core.scala 141:18]
  assign Cp0_io_memoryUnit_in_inst_1_ex_excode = MemoryUnit_io_cp0_in_inst_1_ex_excode; // @[Core.scala 141:18]
  assign Cp0_io_tlb_0_vpn2 = io_inst_tlb2_vpn; // @[Core.scala 128:22]
  assign Cp0_io_tlb_1_vpn2 = io_data_tlb_vpn2; // @[Core.scala 129:22]
  assign MemoryStage_clock = clock;
  assign MemoryStage_reset = reset;
  assign MemoryStage_io_ctrl_allow_to_go = Ctrl_io_memoryUnit_allow_to_go; // @[Core.scala 136:32]
  assign MemoryStage_io_ctrl_clear_0 = Ctrl_io_memoryUnit_do_flush; // @[Core.scala 137:32]
  assign MemoryStage_io_ctrl_clear_1 = Ctrl_io_memoryUnit_do_flush; // @[Core.scala 138:32]
  assign MemoryStage_io_executeUnit_inst0_pc = ExecuteUnit_io_memoryStage_inst0_pc; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_inst_info_fusel = ExecuteUnit_io_memoryStage_inst0_inst_info_fusel; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_inst_info_op = ExecuteUnit_io_memoryStage_inst0_inst_info_op; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_inst_info_reg_wen = ExecuteUnit_io_memoryStage_inst0_inst_info_reg_wen; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_inst_info_reg_waddr = ExecuteUnit_io_memoryStage_inst0_inst_info_reg_waddr; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_inst_info_inst = ExecuteUnit_io_memoryStage_inst0_inst_info_inst; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_rd_info_wdata = ExecuteUnit_io_memoryStage_inst0_rd_info_wdata; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_ex_flush_req = ExecuteUnit_io_memoryStage_inst0_ex_flush_req; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_ex_eret = ExecuteUnit_io_memoryStage_inst0_ex_eret; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_ex_badvaddr = ExecuteUnit_io_memoryStage_inst0_ex_badvaddr; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_ex_bd = ExecuteUnit_io_memoryStage_inst0_ex_bd; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_ex_excode = ExecuteUnit_io_memoryStage_inst0_ex_excode; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_cp0_cp0_count = ExecuteUnit_io_memoryStage_inst0_cp0_cp0_count; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_cp0_cp0_random = ExecuteUnit_io_memoryStage_inst0_cp0_cp0_random; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_cp0_cp0_cause = ExecuteUnit_io_memoryStage_inst0_cp0_cp0_cause; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_mem_en = ExecuteUnit_io_memoryStage_inst0_mem_en; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_mem_inst_info_op = ExecuteUnit_io_memoryStage_inst0_mem_inst_info_op; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_mem_addr = ExecuteUnit_io_memoryStage_inst0_mem_addr; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_mem_wdata = ExecuteUnit_io_memoryStage_inst0_mem_wdata; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_mem_sel_0 = ExecuteUnit_io_memoryStage_inst0_mem_sel_0; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst0_mem_sel_1 = ExecuteUnit_io_memoryStage_inst0_mem_sel_1; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_pc = ExecuteUnit_io_memoryStage_inst1_pc; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_inst_info_fusel = ExecuteUnit_io_memoryStage_inst1_inst_info_fusel; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_inst_info_reg_wen = ExecuteUnit_io_memoryStage_inst1_inst_info_reg_wen; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_inst_info_reg_waddr = ExecuteUnit_io_memoryStage_inst1_inst_info_reg_waddr; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_rd_info_wdata = ExecuteUnit_io_memoryStage_inst1_rd_info_wdata; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_ex_flush_req = ExecuteUnit_io_memoryStage_inst1_ex_flush_req; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_ex_eret = ExecuteUnit_io_memoryStage_inst1_ex_eret; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_ex_badvaddr = ExecuteUnit_io_memoryStage_inst1_ex_badvaddr; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_ex_bd = ExecuteUnit_io_memoryStage_inst1_ex_bd; // @[Core.scala 124:27]
  assign MemoryStage_io_executeUnit_inst1_ex_excode = ExecuteUnit_io_memoryStage_inst1_ex_excode; // @[Core.scala 124:27]
  assign MemoryUnit_io_ctrl_allow_to_go = Ctrl_io_memoryUnit_allow_to_go; // @[Core.scala 40:19]
  assign MemoryUnit_io_memoryStage_inst0_pc = MemoryStage_io_memoryUnit_inst0_pc; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_inst_info_fusel = MemoryStage_io_memoryUnit_inst0_inst_info_fusel; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_inst_info_op = MemoryStage_io_memoryUnit_inst0_inst_info_op; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_inst_info_reg_wen = MemoryStage_io_memoryUnit_inst0_inst_info_reg_wen; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_inst_info_reg_waddr = MemoryStage_io_memoryUnit_inst0_inst_info_reg_waddr; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_inst_info_inst = MemoryStage_io_memoryUnit_inst0_inst_info_inst; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_rd_info_wdata = MemoryStage_io_memoryUnit_inst0_rd_info_wdata; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_ex_flush_req = MemoryStage_io_memoryUnit_inst0_ex_flush_req; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_ex_eret = MemoryStage_io_memoryUnit_inst0_ex_eret; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_ex_badvaddr = MemoryStage_io_memoryUnit_inst0_ex_badvaddr; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_ex_bd = MemoryStage_io_memoryUnit_inst0_ex_bd; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_ex_excode = MemoryStage_io_memoryUnit_inst0_ex_excode; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_cp0_cp0_count = MemoryStage_io_memoryUnit_inst0_cp0_cp0_count; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_cp0_cp0_random = MemoryStage_io_memoryUnit_inst0_cp0_cp0_random; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_cp0_cp0_cause = MemoryStage_io_memoryUnit_inst0_cp0_cp0_cause; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_mem_en = MemoryStage_io_memoryUnit_inst0_mem_en; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_mem_inst_info_op = MemoryStage_io_memoryUnit_inst0_mem_inst_info_op; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_mem_addr = MemoryStage_io_memoryUnit_inst0_mem_addr; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_mem_wdata = MemoryStage_io_memoryUnit_inst0_mem_wdata; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_mem_sel_0 = MemoryStage_io_memoryUnit_inst0_mem_sel_0; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst0_mem_sel_1 = MemoryStage_io_memoryUnit_inst0_mem_sel_1; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_pc = MemoryStage_io_memoryUnit_inst1_pc; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_inst_info_fusel = MemoryStage_io_memoryUnit_inst1_inst_info_fusel; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_inst_info_reg_wen = MemoryStage_io_memoryUnit_inst1_inst_info_reg_wen; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_inst_info_reg_waddr = MemoryStage_io_memoryUnit_inst1_inst_info_reg_waddr; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_rd_info_wdata = MemoryStage_io_memoryUnit_inst1_rd_info_wdata; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_ex_flush_req = MemoryStage_io_memoryUnit_inst1_ex_flush_req; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_ex_eret = MemoryStage_io_memoryUnit_inst1_ex_eret; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_ex_badvaddr = MemoryStage_io_memoryUnit_inst1_ex_badvaddr; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_ex_bd = MemoryStage_io_memoryUnit_inst1_ex_bd; // @[Core.scala 140:26]
  assign MemoryUnit_io_memoryStage_inst1_ex_excode = MemoryStage_io_memoryUnit_inst1_ex_excode; // @[Core.scala 140:26]
  assign MemoryUnit_io_cp0_out_flush = Cp0_io_memoryUnit_out_flush; // @[Core.scala 141:18]
  assign MemoryUnit_io_cp0_out_flush_pc = Cp0_io_memoryUnit_out_flush_pc; // @[Core.scala 141:18]
  assign MemoryUnit_io_dataMemory_in_tlb_invalid = io_data_data_tlb_invalid; // @[Core.scala 144:40]
  assign MemoryUnit_io_dataMemory_in_tlb_refill = io_data_data_tlb_refill; // @[Core.scala 145:40]
  assign MemoryUnit_io_dataMemory_in_tlb_modify = io_data_data_tlb_mod; // @[Core.scala 146:40]
  assign MemoryUnit_io_dataMemory_in_rdata = io_data_M_rdata; // @[Core.scala 147:40]
  assign WriteBackStage_clock = clock;
  assign WriteBackStage_reset = reset;
  assign WriteBackStage_io_ctrl_allow_to_go = Ctrl_io_writeBackUnit_allow_to_go; // @[Core.scala 155:35]
  assign WriteBackStage_io_memoryUnit_inst0_pc = MemoryUnit_io_writeBackStage_inst0_pc; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst0_inst_info_reg_wen = MemoryUnit_io_writeBackStage_inst0_inst_info_reg_wen; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst0_inst_info_reg_waddr = MemoryUnit_io_writeBackStage_inst0_inst_info_reg_waddr
    ; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst0_rd_info_wdata = MemoryUnit_io_writeBackStage_inst0_rd_info_wdata; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst0_ex_flush_req = MemoryUnit_io_writeBackStage_inst0_ex_flush_req; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst0_ex_excode = MemoryUnit_io_writeBackStage_inst0_ex_excode; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst0_cp0_cp0_count = MemoryUnit_io_writeBackStage_inst0_cp0_cp0_count; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst0_cp0_cp0_random = MemoryUnit_io_writeBackStage_inst0_cp0_cp0_random; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst0_cp0_cp0_cause = MemoryUnit_io_writeBackStage_inst0_cp0_cp0_cause; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst1_pc = MemoryUnit_io_writeBackStage_inst1_pc; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst1_inst_info_reg_wen = MemoryUnit_io_writeBackStage_inst1_inst_info_reg_wen; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst1_inst_info_reg_waddr = MemoryUnit_io_writeBackStage_inst1_inst_info_reg_waddr
    ; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst1_rd_info_wdata = MemoryUnit_io_writeBackStage_inst1_rd_info_wdata; // @[Core.scala 154:29]
  assign WriteBackStage_io_memoryUnit_inst1_ex_flush_req = MemoryUnit_io_writeBackStage_inst1_ex_flush_req; // @[Core.scala 154:29]
  assign WriteBackUnit_clock = clock;
  assign WriteBackUnit_reset = reset;
  assign WriteBackUnit_io_ctrl_allow_to_go = Ctrl_io_writeBackUnit_allow_to_go; // @[Core.scala 160:22]
  assign WriteBackUnit_io_writeBackStage_inst0_pc = WriteBackStage_io_writeBackUnit_inst0_pc; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst0_inst_info_reg_wen =
    WriteBackStage_io_writeBackUnit_inst0_inst_info_reg_wen; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst0_inst_info_reg_waddr =
    WriteBackStage_io_writeBackUnit_inst0_inst_info_reg_waddr; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst0_rd_info_wdata = WriteBackStage_io_writeBackUnit_inst0_rd_info_wdata; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst0_ex_flush_req = WriteBackStage_io_writeBackUnit_inst0_ex_flush_req; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst0_ex_excode = WriteBackStage_io_writeBackUnit_inst0_ex_excode; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_count = WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_count; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_random = WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_random; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst0_cp0_cp0_cause = WriteBackStage_io_writeBackUnit_inst0_cp0_cp0_cause; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst1_pc = WriteBackStage_io_writeBackUnit_inst1_pc; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst1_inst_info_reg_wen =
    WriteBackStage_io_writeBackUnit_inst1_inst_info_reg_wen; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst1_inst_info_reg_waddr =
    WriteBackStage_io_writeBackUnit_inst1_inst_info_reg_waddr; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst1_rd_info_wdata = WriteBackStage_io_writeBackUnit_inst1_rd_info_wdata; // @[Core.scala 159:32]
  assign WriteBackUnit_io_writeBackStage_inst1_ex_flush_req = WriteBackStage_io_writeBackUnit_inst1_ex_flush_req; // @[Core.scala 159:32]
endmodule
module SimpleDualPortRam(
  input         clock,
  input         reset,
  input  [8:0]  io_raddr,
  output [31:0] io_rdata,
  input  [8:0]  io_waddr,
  input         io_wen,
  input  [3:0]  io_wstrb,
  input  [31:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] bank_0 [0:511]; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_0_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  wire [8:0] bank_0_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_0_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_0_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [8:0] bank_0_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_0_MPORT_mask; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_0_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  reg  bank_0_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_0_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_1 [0:511]; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_1_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  wire [8:0] bank_1_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_1_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_1_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [8:0] bank_1_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_1_MPORT_mask; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_1_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  reg  bank_1_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_1_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_2 [0:511]; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_2_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  wire [8:0] bank_2_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_2_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_2_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [8:0] bank_2_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_2_MPORT_mask; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_2_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  reg  bank_2_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_2_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_3 [0:511]; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_3_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  wire [8:0] bank_3_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_3_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_3_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [8:0] bank_3_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_3_MPORT_mask; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_3_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  reg  bank_3_io_rdata_MPORT_en_pipe_0;
  reg [8:0] bank_3_io_rdata_MPORT_addr_pipe_0;
  wire  _T_2 = |io_wstrb | ~io_wen; // @[SimpleDualPortRam.scala 64:20]
  wire [15:0] io_rdata_lo = {bank_1_io_rdata_MPORT_data,bank_0_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 70:44]
  wire [15:0] io_rdata_hi = {bank_3_io_rdata_MPORT_data,bank_2_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 70:44]
  assign bank_0_io_rdata_MPORT_en = bank_0_io_rdata_MPORT_en_pipe_0;
  assign bank_0_io_rdata_MPORT_addr = bank_0_io_rdata_MPORT_addr_pipe_0;
  assign bank_0_io_rdata_MPORT_data = bank_0[bank_0_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 68:29]
  assign bank_0_MPORT_data = io_wdata[7:0];
  assign bank_0_MPORT_addr = io_waddr;
  assign bank_0_MPORT_mask = io_wstrb[0];
  assign bank_0_MPORT_en = io_wen;
  assign bank_1_io_rdata_MPORT_en = bank_1_io_rdata_MPORT_en_pipe_0;
  assign bank_1_io_rdata_MPORT_addr = bank_1_io_rdata_MPORT_addr_pipe_0;
  assign bank_1_io_rdata_MPORT_data = bank_1[bank_1_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 68:29]
  assign bank_1_MPORT_data = io_wdata[15:8];
  assign bank_1_MPORT_addr = io_waddr;
  assign bank_1_MPORT_mask = io_wstrb[1];
  assign bank_1_MPORT_en = io_wen;
  assign bank_2_io_rdata_MPORT_en = bank_2_io_rdata_MPORT_en_pipe_0;
  assign bank_2_io_rdata_MPORT_addr = bank_2_io_rdata_MPORT_addr_pipe_0;
  assign bank_2_io_rdata_MPORT_data = bank_2[bank_2_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 68:29]
  assign bank_2_MPORT_data = io_wdata[23:16];
  assign bank_2_MPORT_addr = io_waddr;
  assign bank_2_MPORT_mask = io_wstrb[2];
  assign bank_2_MPORT_en = io_wen;
  assign bank_3_io_rdata_MPORT_en = bank_3_io_rdata_MPORT_en_pipe_0;
  assign bank_3_io_rdata_MPORT_addr = bank_3_io_rdata_MPORT_addr_pipe_0;
  assign bank_3_io_rdata_MPORT_data = bank_3[bank_3_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 68:29]
  assign bank_3_MPORT_data = io_wdata[31:24];
  assign bank_3_MPORT_addr = io_waddr;
  assign bank_3_MPORT_mask = io_wstrb[3];
  assign bank_3_MPORT_en = io_wen;
  assign io_rdata = {io_rdata_hi,io_rdata_lo}; // @[SimpleDualPortRam.scala 70:44]
  always @(posedge clock) begin
    if (bank_0_MPORT_en & bank_0_MPORT_mask) begin
      bank_0[bank_0_MPORT_addr] <= bank_0_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
    end
    bank_0_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_0_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_1_MPORT_en & bank_1_MPORT_mask) begin
      bank_1[bank_1_MPORT_addr] <= bank_1_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
    end
    bank_1_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_1_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_2_MPORT_en & bank_2_MPORT_mask) begin
      bank_2[bank_2_MPORT_addr] <= bank_2_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
    end
    bank_2_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_2_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_3_MPORT_en & bank_3_MPORT_mask) begin
      bank_3[bank_3_MPORT_addr] <= bank_3_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
    end
    bank_3_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_3_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed: when write port enable is high, write vector cannot be all 0\n    at SimpleDualPortRam.scala:63 assert(\n"
            ); // @[SimpleDualPortRam.scala 63:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & ~reset) begin
          $fatal; // @[SimpleDualPortRam.scala 63:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_0[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_1[initvar] = _RAND_3[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_2[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    bank_3[initvar] = _RAND_9[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bank_0_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bank_0_io_rdata_MPORT_addr_pipe_0 = _RAND_2[8:0];
  _RAND_4 = {1{`RANDOM}};
  bank_1_io_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  bank_1_io_rdata_MPORT_addr_pipe_0 = _RAND_5[8:0];
  _RAND_7 = {1{`RANDOM}};
  bank_2_io_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  bank_2_io_rdata_MPORT_addr_pipe_0 = _RAND_8[8:0];
  _RAND_10 = {1{`RANDOM}};
  bank_3_io_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  bank_3_io_rdata_MPORT_addr_pipe_0 = _RAND_11[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleDualPortRam_1(
  input         clock,
  input         reset,
  input  [5:0]  io_raddr,
  output [19:0] io_rdata,
  input  [5:0]  io_waddr,
  input         io_wen,
  input         io_wstrb,
  input  [19:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] bank [0:63]; // @[SimpleDualPortRam.scala 78:29]
  wire  bank_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 78:29]
  wire [5:0] bank_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 78:29]
  wire [19:0] bank_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 78:29]
  wire [19:0] bank_MPORT_data; // @[SimpleDualPortRam.scala 78:29]
  wire [5:0] bank_MPORT_addr; // @[SimpleDualPortRam.scala 78:29]
  wire  bank_MPORT_mask; // @[SimpleDualPortRam.scala 78:29]
  wire  bank_MPORT_en; // @[SimpleDualPortRam.scala 78:29]
  reg  bank_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_io_rdata_MPORT_addr_pipe_0;
  wire  _T_2 = |io_wstrb | ~io_wen; // @[SimpleDualPortRam.scala 64:20]
  wire [31:0] _GEN_7 = {{12'd0}, bank_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 80:20 81:18 83:18]
  assign bank_io_rdata_MPORT_en = bank_io_rdata_MPORT_en_pipe_0;
  assign bank_io_rdata_MPORT_addr = bank_io_rdata_MPORT_addr_pipe_0;
  assign bank_io_rdata_MPORT_data = bank[bank_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 78:29]
  assign bank_MPORT_data = io_wdata;
  assign bank_MPORT_addr = io_waddr;
  assign bank_MPORT_mask = 1'h1;
  assign bank_MPORT_en = io_wen;
  assign io_rdata = _GEN_7[19:0];
  always @(posedge clock) begin
    if (bank_MPORT_en & bank_MPORT_mask) begin
      bank[bank_MPORT_addr] <= bank_MPORT_data; // @[SimpleDualPortRam.scala 78:29]
    end
    bank_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed: when write port enable is high, write vector cannot be all 0\n    at SimpleDualPortRam.scala:63 assert(\n"
            ); // @[SimpleDualPortRam.scala 63:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & ~reset) begin
          $fatal; // @[SimpleDualPortRam.scala 63:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bank_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bank_io_rdata_MPORT_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input         clock,
  input         reset,
  input         io_cpu_req,
  input  [31:0] io_cpu_addr_0,
  input  [31:0] io_cpu_addr_1,
  output [31:0] io_cpu_inst_0,
  output [31:0] io_cpu_inst_1,
  output        io_cpu_inst_valid_0,
  output        io_cpu_inst_valid_1,
  input         io_cpu_cpu_stall,
  output        io_cpu_icache_stall,
  output        io_cpu_tlb1_invalid,
  output [18:0] io_cpu_tlb2_vpn,
  input         io_cpu_tlb2_found,
  input  [19:0] io_cpu_tlb2_entry_pfn_0,
  input  [19:0] io_cpu_tlb2_entry_pfn_1,
  input         io_cpu_tlb2_entry_c_0,
  input         io_cpu_tlb2_entry_c_1,
  input         io_cpu_tlb2_entry_v_0,
  input         io_cpu_tlb2_entry_v_1,
  input         io_cpu_fence_value,
  input  [31:0] io_cpu_fence_addr,
  input         io_cpu_fence_tlb,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output [7:0]  io_axi_ar_bits_len,
  output [2:0]  io_axi_ar_bits_size,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [31:0] io_axi_r_bits_data,
  input         io_axi_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
`endif // RANDOMIZE_REG_INIT
  wire  bank_clock; // @[ICache.scala 122:22]
  wire  bank_reset; // @[ICache.scala 122:22]
  wire [8:0] bank_io_raddr; // @[ICache.scala 122:22]
  wire [31:0] bank_io_rdata; // @[ICache.scala 122:22]
  wire [8:0] bank_io_waddr; // @[ICache.scala 122:22]
  wire  bank_io_wen; // @[ICache.scala 122:22]
  wire [3:0] bank_io_wstrb; // @[ICache.scala 122:22]
  wire [31:0] bank_io_wdata; // @[ICache.scala 122:22]
  wire  tag_bram_clock; // @[ICache.scala 132:26]
  wire  tag_bram_reset; // @[ICache.scala 132:26]
  wire [5:0] tag_bram_io_raddr; // @[ICache.scala 132:26]
  wire [19:0] tag_bram_io_rdata; // @[ICache.scala 132:26]
  wire [5:0] tag_bram_io_waddr; // @[ICache.scala 132:26]
  wire  tag_bram_io_wen; // @[ICache.scala 132:26]
  wire  tag_bram_io_wstrb; // @[ICache.scala 132:26]
  wire [19:0] tag_bram_io_wdata; // @[ICache.scala 132:26]
  wire  bank_1_clock; // @[ICache.scala 122:22]
  wire  bank_1_reset; // @[ICache.scala 122:22]
  wire [8:0] bank_1_io_raddr; // @[ICache.scala 122:22]
  wire [31:0] bank_1_io_rdata; // @[ICache.scala 122:22]
  wire [8:0] bank_1_io_waddr; // @[ICache.scala 122:22]
  wire  bank_1_io_wen; // @[ICache.scala 122:22]
  wire [3:0] bank_1_io_wstrb; // @[ICache.scala 122:22]
  wire [31:0] bank_1_io_wdata; // @[ICache.scala 122:22]
  wire  tag_bram_1_clock; // @[ICache.scala 132:26]
  wire  tag_bram_1_reset; // @[ICache.scala 132:26]
  wire [5:0] tag_bram_1_io_raddr; // @[ICache.scala 132:26]
  wire [19:0] tag_bram_1_io_rdata; // @[ICache.scala 132:26]
  wire [5:0] tag_bram_1_io_waddr; // @[ICache.scala 132:26]
  wire  tag_bram_1_io_wen; // @[ICache.scala 132:26]
  wire  tag_bram_1_io_wstrb; // @[ICache.scala 132:26]
  wire [19:0] tag_bram_1_io_wdata; // @[ICache.scala 132:26]
  wire  bank_2_clock; // @[ICache.scala 122:22]
  wire  bank_2_reset; // @[ICache.scala 122:22]
  wire [8:0] bank_2_io_raddr; // @[ICache.scala 122:22]
  wire [31:0] bank_2_io_rdata; // @[ICache.scala 122:22]
  wire [8:0] bank_2_io_waddr; // @[ICache.scala 122:22]
  wire  bank_2_io_wen; // @[ICache.scala 122:22]
  wire [3:0] bank_2_io_wstrb; // @[ICache.scala 122:22]
  wire [31:0] bank_2_io_wdata; // @[ICache.scala 122:22]
  wire  tag_bram_2_clock; // @[ICache.scala 132:26]
  wire  tag_bram_2_reset; // @[ICache.scala 132:26]
  wire [5:0] tag_bram_2_io_raddr; // @[ICache.scala 132:26]
  wire [19:0] tag_bram_2_io_rdata; // @[ICache.scala 132:26]
  wire [5:0] tag_bram_2_io_waddr; // @[ICache.scala 132:26]
  wire  tag_bram_2_io_wen; // @[ICache.scala 132:26]
  wire  tag_bram_2_io_wstrb; // @[ICache.scala 132:26]
  wire [19:0] tag_bram_2_io_wdata; // @[ICache.scala 132:26]
  wire  bank_3_clock; // @[ICache.scala 122:22]
  wire  bank_3_reset; // @[ICache.scala 122:22]
  wire [8:0] bank_3_io_raddr; // @[ICache.scala 122:22]
  wire [31:0] bank_3_io_rdata; // @[ICache.scala 122:22]
  wire [8:0] bank_3_io_waddr; // @[ICache.scala 122:22]
  wire  bank_3_io_wen; // @[ICache.scala 122:22]
  wire [3:0] bank_3_io_wstrb; // @[ICache.scala 122:22]
  wire [31:0] bank_3_io_wdata; // @[ICache.scala 122:22]
  wire  tag_bram_3_clock; // @[ICache.scala 132:26]
  wire  tag_bram_3_reset; // @[ICache.scala 132:26]
  wire [5:0] tag_bram_3_io_raddr; // @[ICache.scala 132:26]
  wire [19:0] tag_bram_3_io_rdata; // @[ICache.scala 132:26]
  wire [5:0] tag_bram_3_io_waddr; // @[ICache.scala 132:26]
  wire  tag_bram_3_io_wen; // @[ICache.scala 132:26]
  wire  tag_bram_3_io_wstrb; // @[ICache.scala 132:26]
  wire [19:0] tag_bram_3_io_wdata; // @[ICache.scala 132:26]
  reg [2:0] state; // @[ICache.scala 39:81]
  reg  valid_0_0; // @[ICache.scala 52:22]
  reg  valid_0_1; // @[ICache.scala 52:22]
  reg  valid_1_0; // @[ICache.scala 52:22]
  reg  valid_1_1; // @[ICache.scala 52:22]
  reg  valid_2_0; // @[ICache.scala 52:22]
  reg  valid_2_1; // @[ICache.scala 52:22]
  reg  valid_3_0; // @[ICache.scala 52:22]
  reg  valid_3_1; // @[ICache.scala 52:22]
  reg  valid_4_0; // @[ICache.scala 52:22]
  reg  valid_4_1; // @[ICache.scala 52:22]
  reg  valid_5_0; // @[ICache.scala 52:22]
  reg  valid_5_1; // @[ICache.scala 52:22]
  reg  valid_6_0; // @[ICache.scala 52:22]
  reg  valid_6_1; // @[ICache.scala 52:22]
  reg  valid_7_0; // @[ICache.scala 52:22]
  reg  valid_7_1; // @[ICache.scala 52:22]
  reg  valid_8_0; // @[ICache.scala 52:22]
  reg  valid_8_1; // @[ICache.scala 52:22]
  reg  valid_9_0; // @[ICache.scala 52:22]
  reg  valid_9_1; // @[ICache.scala 52:22]
  reg  valid_10_0; // @[ICache.scala 52:22]
  reg  valid_10_1; // @[ICache.scala 52:22]
  reg  valid_11_0; // @[ICache.scala 52:22]
  reg  valid_11_1; // @[ICache.scala 52:22]
  reg  valid_12_0; // @[ICache.scala 52:22]
  reg  valid_12_1; // @[ICache.scala 52:22]
  reg  valid_13_0; // @[ICache.scala 52:22]
  reg  valid_13_1; // @[ICache.scala 52:22]
  reg  valid_14_0; // @[ICache.scala 52:22]
  reg  valid_14_1; // @[ICache.scala 52:22]
  reg  valid_15_0; // @[ICache.scala 52:22]
  reg  valid_15_1; // @[ICache.scala 52:22]
  reg  valid_16_0; // @[ICache.scala 52:22]
  reg  valid_16_1; // @[ICache.scala 52:22]
  reg  valid_17_0; // @[ICache.scala 52:22]
  reg  valid_17_1; // @[ICache.scala 52:22]
  reg  valid_18_0; // @[ICache.scala 52:22]
  reg  valid_18_1; // @[ICache.scala 52:22]
  reg  valid_19_0; // @[ICache.scala 52:22]
  reg  valid_19_1; // @[ICache.scala 52:22]
  reg  valid_20_0; // @[ICache.scala 52:22]
  reg  valid_20_1; // @[ICache.scala 52:22]
  reg  valid_21_0; // @[ICache.scala 52:22]
  reg  valid_21_1; // @[ICache.scala 52:22]
  reg  valid_22_0; // @[ICache.scala 52:22]
  reg  valid_22_1; // @[ICache.scala 52:22]
  reg  valid_23_0; // @[ICache.scala 52:22]
  reg  valid_23_1; // @[ICache.scala 52:22]
  reg  valid_24_0; // @[ICache.scala 52:22]
  reg  valid_24_1; // @[ICache.scala 52:22]
  reg  valid_25_0; // @[ICache.scala 52:22]
  reg  valid_25_1; // @[ICache.scala 52:22]
  reg  valid_26_0; // @[ICache.scala 52:22]
  reg  valid_26_1; // @[ICache.scala 52:22]
  reg  valid_27_0; // @[ICache.scala 52:22]
  reg  valid_27_1; // @[ICache.scala 52:22]
  reg  valid_28_0; // @[ICache.scala 52:22]
  reg  valid_28_1; // @[ICache.scala 52:22]
  reg  valid_29_0; // @[ICache.scala 52:22]
  reg  valid_29_1; // @[ICache.scala 52:22]
  reg  valid_30_0; // @[ICache.scala 52:22]
  reg  valid_30_1; // @[ICache.scala 52:22]
  reg  valid_31_0; // @[ICache.scala 52:22]
  reg  valid_31_1; // @[ICache.scala 52:22]
  reg  valid_32_0; // @[ICache.scala 52:22]
  reg  valid_32_1; // @[ICache.scala 52:22]
  reg  valid_33_0; // @[ICache.scala 52:22]
  reg  valid_33_1; // @[ICache.scala 52:22]
  reg  valid_34_0; // @[ICache.scala 52:22]
  reg  valid_34_1; // @[ICache.scala 52:22]
  reg  valid_35_0; // @[ICache.scala 52:22]
  reg  valid_35_1; // @[ICache.scala 52:22]
  reg  valid_36_0; // @[ICache.scala 52:22]
  reg  valid_36_1; // @[ICache.scala 52:22]
  reg  valid_37_0; // @[ICache.scala 52:22]
  reg  valid_37_1; // @[ICache.scala 52:22]
  reg  valid_38_0; // @[ICache.scala 52:22]
  reg  valid_38_1; // @[ICache.scala 52:22]
  reg  valid_39_0; // @[ICache.scala 52:22]
  reg  valid_39_1; // @[ICache.scala 52:22]
  reg  valid_40_0; // @[ICache.scala 52:22]
  reg  valid_40_1; // @[ICache.scala 52:22]
  reg  valid_41_0; // @[ICache.scala 52:22]
  reg  valid_41_1; // @[ICache.scala 52:22]
  reg  valid_42_0; // @[ICache.scala 52:22]
  reg  valid_42_1; // @[ICache.scala 52:22]
  reg  valid_43_0; // @[ICache.scala 52:22]
  reg  valid_43_1; // @[ICache.scala 52:22]
  reg  valid_44_0; // @[ICache.scala 52:22]
  reg  valid_44_1; // @[ICache.scala 52:22]
  reg  valid_45_0; // @[ICache.scala 52:22]
  reg  valid_45_1; // @[ICache.scala 52:22]
  reg  valid_46_0; // @[ICache.scala 52:22]
  reg  valid_46_1; // @[ICache.scala 52:22]
  reg  valid_47_0; // @[ICache.scala 52:22]
  reg  valid_47_1; // @[ICache.scala 52:22]
  reg  valid_48_0; // @[ICache.scala 52:22]
  reg  valid_48_1; // @[ICache.scala 52:22]
  reg  valid_49_0; // @[ICache.scala 52:22]
  reg  valid_49_1; // @[ICache.scala 52:22]
  reg  valid_50_0; // @[ICache.scala 52:22]
  reg  valid_50_1; // @[ICache.scala 52:22]
  reg  valid_51_0; // @[ICache.scala 52:22]
  reg  valid_51_1; // @[ICache.scala 52:22]
  reg  valid_52_0; // @[ICache.scala 52:22]
  reg  valid_52_1; // @[ICache.scala 52:22]
  reg  valid_53_0; // @[ICache.scala 52:22]
  reg  valid_53_1; // @[ICache.scala 52:22]
  reg  valid_54_0; // @[ICache.scala 52:22]
  reg  valid_54_1; // @[ICache.scala 52:22]
  reg  valid_55_0; // @[ICache.scala 52:22]
  reg  valid_55_1; // @[ICache.scala 52:22]
  reg  valid_56_0; // @[ICache.scala 52:22]
  reg  valid_56_1; // @[ICache.scala 52:22]
  reg  valid_57_0; // @[ICache.scala 52:22]
  reg  valid_57_1; // @[ICache.scala 52:22]
  reg  valid_58_0; // @[ICache.scala 52:22]
  reg  valid_58_1; // @[ICache.scala 52:22]
  reg  valid_59_0; // @[ICache.scala 52:22]
  reg  valid_59_1; // @[ICache.scala 52:22]
  reg  valid_60_0; // @[ICache.scala 52:22]
  reg  valid_60_1; // @[ICache.scala 52:22]
  reg  valid_61_0; // @[ICache.scala 52:22]
  reg  valid_61_1; // @[ICache.scala 52:22]
  reg  valid_62_0; // @[ICache.scala 52:22]
  reg  valid_62_1; // @[ICache.scala 52:22]
  reg  valid_63_0; // @[ICache.scala 52:22]
  reg  valid_63_1; // @[ICache.scala 52:22]
  reg  valid_64_0; // @[ICache.scala 52:22]
  reg  valid_64_1; // @[ICache.scala 52:22]
  reg  valid_65_0; // @[ICache.scala 52:22]
  reg  valid_65_1; // @[ICache.scala 52:22]
  reg  valid_66_0; // @[ICache.scala 52:22]
  reg  valid_66_1; // @[ICache.scala 52:22]
  reg  valid_67_0; // @[ICache.scala 52:22]
  reg  valid_67_1; // @[ICache.scala 52:22]
  reg  valid_68_0; // @[ICache.scala 52:22]
  reg  valid_68_1; // @[ICache.scala 52:22]
  reg  valid_69_0; // @[ICache.scala 52:22]
  reg  valid_69_1; // @[ICache.scala 52:22]
  reg  valid_70_0; // @[ICache.scala 52:22]
  reg  valid_70_1; // @[ICache.scala 52:22]
  reg  valid_71_0; // @[ICache.scala 52:22]
  reg  valid_71_1; // @[ICache.scala 52:22]
  reg  valid_72_0; // @[ICache.scala 52:22]
  reg  valid_72_1; // @[ICache.scala 52:22]
  reg  valid_73_0; // @[ICache.scala 52:22]
  reg  valid_73_1; // @[ICache.scala 52:22]
  reg  valid_74_0; // @[ICache.scala 52:22]
  reg  valid_74_1; // @[ICache.scala 52:22]
  reg  valid_75_0; // @[ICache.scala 52:22]
  reg  valid_75_1; // @[ICache.scala 52:22]
  reg  valid_76_0; // @[ICache.scala 52:22]
  reg  valid_76_1; // @[ICache.scala 52:22]
  reg  valid_77_0; // @[ICache.scala 52:22]
  reg  valid_77_1; // @[ICache.scala 52:22]
  reg  valid_78_0; // @[ICache.scala 52:22]
  reg  valid_78_1; // @[ICache.scala 52:22]
  reg  valid_79_0; // @[ICache.scala 52:22]
  reg  valid_79_1; // @[ICache.scala 52:22]
  reg  valid_80_0; // @[ICache.scala 52:22]
  reg  valid_80_1; // @[ICache.scala 52:22]
  reg  valid_81_0; // @[ICache.scala 52:22]
  reg  valid_81_1; // @[ICache.scala 52:22]
  reg  valid_82_0; // @[ICache.scala 52:22]
  reg  valid_82_1; // @[ICache.scala 52:22]
  reg  valid_83_0; // @[ICache.scala 52:22]
  reg  valid_83_1; // @[ICache.scala 52:22]
  reg  valid_84_0; // @[ICache.scala 52:22]
  reg  valid_84_1; // @[ICache.scala 52:22]
  reg  valid_85_0; // @[ICache.scala 52:22]
  reg  valid_85_1; // @[ICache.scala 52:22]
  reg  valid_86_0; // @[ICache.scala 52:22]
  reg  valid_86_1; // @[ICache.scala 52:22]
  reg  valid_87_0; // @[ICache.scala 52:22]
  reg  valid_87_1; // @[ICache.scala 52:22]
  reg  valid_88_0; // @[ICache.scala 52:22]
  reg  valid_88_1; // @[ICache.scala 52:22]
  reg  valid_89_0; // @[ICache.scala 52:22]
  reg  valid_89_1; // @[ICache.scala 52:22]
  reg  valid_90_0; // @[ICache.scala 52:22]
  reg  valid_90_1; // @[ICache.scala 52:22]
  reg  valid_91_0; // @[ICache.scala 52:22]
  reg  valid_91_1; // @[ICache.scala 52:22]
  reg  valid_92_0; // @[ICache.scala 52:22]
  reg  valid_92_1; // @[ICache.scala 52:22]
  reg  valid_93_0; // @[ICache.scala 52:22]
  reg  valid_93_1; // @[ICache.scala 52:22]
  reg  valid_94_0; // @[ICache.scala 52:22]
  reg  valid_94_1; // @[ICache.scala 52:22]
  reg  valid_95_0; // @[ICache.scala 52:22]
  reg  valid_95_1; // @[ICache.scala 52:22]
  reg  valid_96_0; // @[ICache.scala 52:22]
  reg  valid_96_1; // @[ICache.scala 52:22]
  reg  valid_97_0; // @[ICache.scala 52:22]
  reg  valid_97_1; // @[ICache.scala 52:22]
  reg  valid_98_0; // @[ICache.scala 52:22]
  reg  valid_98_1; // @[ICache.scala 52:22]
  reg  valid_99_0; // @[ICache.scala 52:22]
  reg  valid_99_1; // @[ICache.scala 52:22]
  reg  valid_100_0; // @[ICache.scala 52:22]
  reg  valid_100_1; // @[ICache.scala 52:22]
  reg  valid_101_0; // @[ICache.scala 52:22]
  reg  valid_101_1; // @[ICache.scala 52:22]
  reg  valid_102_0; // @[ICache.scala 52:22]
  reg  valid_102_1; // @[ICache.scala 52:22]
  reg  valid_103_0; // @[ICache.scala 52:22]
  reg  valid_103_1; // @[ICache.scala 52:22]
  reg  valid_104_0; // @[ICache.scala 52:22]
  reg  valid_104_1; // @[ICache.scala 52:22]
  reg  valid_105_0; // @[ICache.scala 52:22]
  reg  valid_105_1; // @[ICache.scala 52:22]
  reg  valid_106_0; // @[ICache.scala 52:22]
  reg  valid_106_1; // @[ICache.scala 52:22]
  reg  valid_107_0; // @[ICache.scala 52:22]
  reg  valid_107_1; // @[ICache.scala 52:22]
  reg  valid_108_0; // @[ICache.scala 52:22]
  reg  valid_108_1; // @[ICache.scala 52:22]
  reg  valid_109_0; // @[ICache.scala 52:22]
  reg  valid_109_1; // @[ICache.scala 52:22]
  reg  valid_110_0; // @[ICache.scala 52:22]
  reg  valid_110_1; // @[ICache.scala 52:22]
  reg  valid_111_0; // @[ICache.scala 52:22]
  reg  valid_111_1; // @[ICache.scala 52:22]
  reg  valid_112_0; // @[ICache.scala 52:22]
  reg  valid_112_1; // @[ICache.scala 52:22]
  reg  valid_113_0; // @[ICache.scala 52:22]
  reg  valid_113_1; // @[ICache.scala 52:22]
  reg  valid_114_0; // @[ICache.scala 52:22]
  reg  valid_114_1; // @[ICache.scala 52:22]
  reg  valid_115_0; // @[ICache.scala 52:22]
  reg  valid_115_1; // @[ICache.scala 52:22]
  reg  valid_116_0; // @[ICache.scala 52:22]
  reg  valid_116_1; // @[ICache.scala 52:22]
  reg  valid_117_0; // @[ICache.scala 52:22]
  reg  valid_117_1; // @[ICache.scala 52:22]
  reg  valid_118_0; // @[ICache.scala 52:22]
  reg  valid_118_1; // @[ICache.scala 52:22]
  reg  valid_119_0; // @[ICache.scala 52:22]
  reg  valid_119_1; // @[ICache.scala 52:22]
  reg  valid_120_0; // @[ICache.scala 52:22]
  reg  valid_120_1; // @[ICache.scala 52:22]
  reg  valid_121_0; // @[ICache.scala 52:22]
  reg  valid_121_1; // @[ICache.scala 52:22]
  reg  valid_122_0; // @[ICache.scala 52:22]
  reg  valid_122_1; // @[ICache.scala 52:22]
  reg  valid_123_0; // @[ICache.scala 52:22]
  reg  valid_123_1; // @[ICache.scala 52:22]
  reg  valid_124_0; // @[ICache.scala 52:22]
  reg  valid_124_1; // @[ICache.scala 52:22]
  reg  valid_125_0; // @[ICache.scala 52:22]
  reg  valid_125_1; // @[ICache.scala 52:22]
  reg  valid_126_0; // @[ICache.scala 52:22]
  reg  valid_126_1; // @[ICache.scala 52:22]
  reg  valid_127_0; // @[ICache.scala 52:22]
  reg  valid_127_1; // @[ICache.scala 52:22]
  reg  valid_128_0; // @[ICache.scala 52:22]
  reg  valid_128_1; // @[ICache.scala 52:22]
  reg  valid_129_0; // @[ICache.scala 52:22]
  reg  valid_129_1; // @[ICache.scala 52:22]
  reg  valid_130_0; // @[ICache.scala 52:22]
  reg  valid_130_1; // @[ICache.scala 52:22]
  reg  valid_131_0; // @[ICache.scala 52:22]
  reg  valid_131_1; // @[ICache.scala 52:22]
  reg  valid_132_0; // @[ICache.scala 52:22]
  reg  valid_132_1; // @[ICache.scala 52:22]
  reg  valid_133_0; // @[ICache.scala 52:22]
  reg  valid_133_1; // @[ICache.scala 52:22]
  reg  valid_134_0; // @[ICache.scala 52:22]
  reg  valid_134_1; // @[ICache.scala 52:22]
  reg  valid_135_0; // @[ICache.scala 52:22]
  reg  valid_135_1; // @[ICache.scala 52:22]
  reg  valid_136_0; // @[ICache.scala 52:22]
  reg  valid_136_1; // @[ICache.scala 52:22]
  reg  valid_137_0; // @[ICache.scala 52:22]
  reg  valid_137_1; // @[ICache.scala 52:22]
  reg  valid_138_0; // @[ICache.scala 52:22]
  reg  valid_138_1; // @[ICache.scala 52:22]
  reg  valid_139_0; // @[ICache.scala 52:22]
  reg  valid_139_1; // @[ICache.scala 52:22]
  reg  valid_140_0; // @[ICache.scala 52:22]
  reg  valid_140_1; // @[ICache.scala 52:22]
  reg  valid_141_0; // @[ICache.scala 52:22]
  reg  valid_141_1; // @[ICache.scala 52:22]
  reg  valid_142_0; // @[ICache.scala 52:22]
  reg  valid_142_1; // @[ICache.scala 52:22]
  reg  valid_143_0; // @[ICache.scala 52:22]
  reg  valid_143_1; // @[ICache.scala 52:22]
  reg  valid_144_0; // @[ICache.scala 52:22]
  reg  valid_144_1; // @[ICache.scala 52:22]
  reg  valid_145_0; // @[ICache.scala 52:22]
  reg  valid_145_1; // @[ICache.scala 52:22]
  reg  valid_146_0; // @[ICache.scala 52:22]
  reg  valid_146_1; // @[ICache.scala 52:22]
  reg  valid_147_0; // @[ICache.scala 52:22]
  reg  valid_147_1; // @[ICache.scala 52:22]
  reg  valid_148_0; // @[ICache.scala 52:22]
  reg  valid_148_1; // @[ICache.scala 52:22]
  reg  valid_149_0; // @[ICache.scala 52:22]
  reg  valid_149_1; // @[ICache.scala 52:22]
  reg  valid_150_0; // @[ICache.scala 52:22]
  reg  valid_150_1; // @[ICache.scala 52:22]
  reg  valid_151_0; // @[ICache.scala 52:22]
  reg  valid_151_1; // @[ICache.scala 52:22]
  reg  valid_152_0; // @[ICache.scala 52:22]
  reg  valid_152_1; // @[ICache.scala 52:22]
  reg  valid_153_0; // @[ICache.scala 52:22]
  reg  valid_153_1; // @[ICache.scala 52:22]
  reg  valid_154_0; // @[ICache.scala 52:22]
  reg  valid_154_1; // @[ICache.scala 52:22]
  reg  valid_155_0; // @[ICache.scala 52:22]
  reg  valid_155_1; // @[ICache.scala 52:22]
  reg  valid_156_0; // @[ICache.scala 52:22]
  reg  valid_156_1; // @[ICache.scala 52:22]
  reg  valid_157_0; // @[ICache.scala 52:22]
  reg  valid_157_1; // @[ICache.scala 52:22]
  reg  valid_158_0; // @[ICache.scala 52:22]
  reg  valid_158_1; // @[ICache.scala 52:22]
  reg  valid_159_0; // @[ICache.scala 52:22]
  reg  valid_159_1; // @[ICache.scala 52:22]
  reg  valid_160_0; // @[ICache.scala 52:22]
  reg  valid_160_1; // @[ICache.scala 52:22]
  reg  valid_161_0; // @[ICache.scala 52:22]
  reg  valid_161_1; // @[ICache.scala 52:22]
  reg  valid_162_0; // @[ICache.scala 52:22]
  reg  valid_162_1; // @[ICache.scala 52:22]
  reg  valid_163_0; // @[ICache.scala 52:22]
  reg  valid_163_1; // @[ICache.scala 52:22]
  reg  valid_164_0; // @[ICache.scala 52:22]
  reg  valid_164_1; // @[ICache.scala 52:22]
  reg  valid_165_0; // @[ICache.scala 52:22]
  reg  valid_165_1; // @[ICache.scala 52:22]
  reg  valid_166_0; // @[ICache.scala 52:22]
  reg  valid_166_1; // @[ICache.scala 52:22]
  reg  valid_167_0; // @[ICache.scala 52:22]
  reg  valid_167_1; // @[ICache.scala 52:22]
  reg  valid_168_0; // @[ICache.scala 52:22]
  reg  valid_168_1; // @[ICache.scala 52:22]
  reg  valid_169_0; // @[ICache.scala 52:22]
  reg  valid_169_1; // @[ICache.scala 52:22]
  reg  valid_170_0; // @[ICache.scala 52:22]
  reg  valid_170_1; // @[ICache.scala 52:22]
  reg  valid_171_0; // @[ICache.scala 52:22]
  reg  valid_171_1; // @[ICache.scala 52:22]
  reg  valid_172_0; // @[ICache.scala 52:22]
  reg  valid_172_1; // @[ICache.scala 52:22]
  reg  valid_173_0; // @[ICache.scala 52:22]
  reg  valid_173_1; // @[ICache.scala 52:22]
  reg  valid_174_0; // @[ICache.scala 52:22]
  reg  valid_174_1; // @[ICache.scala 52:22]
  reg  valid_175_0; // @[ICache.scala 52:22]
  reg  valid_175_1; // @[ICache.scala 52:22]
  reg  valid_176_0; // @[ICache.scala 52:22]
  reg  valid_176_1; // @[ICache.scala 52:22]
  reg  valid_177_0; // @[ICache.scala 52:22]
  reg  valid_177_1; // @[ICache.scala 52:22]
  reg  valid_178_0; // @[ICache.scala 52:22]
  reg  valid_178_1; // @[ICache.scala 52:22]
  reg  valid_179_0; // @[ICache.scala 52:22]
  reg  valid_179_1; // @[ICache.scala 52:22]
  reg  valid_180_0; // @[ICache.scala 52:22]
  reg  valid_180_1; // @[ICache.scala 52:22]
  reg  valid_181_0; // @[ICache.scala 52:22]
  reg  valid_181_1; // @[ICache.scala 52:22]
  reg  valid_182_0; // @[ICache.scala 52:22]
  reg  valid_182_1; // @[ICache.scala 52:22]
  reg  valid_183_0; // @[ICache.scala 52:22]
  reg  valid_183_1; // @[ICache.scala 52:22]
  reg  valid_184_0; // @[ICache.scala 52:22]
  reg  valid_184_1; // @[ICache.scala 52:22]
  reg  valid_185_0; // @[ICache.scala 52:22]
  reg  valid_185_1; // @[ICache.scala 52:22]
  reg  valid_186_0; // @[ICache.scala 52:22]
  reg  valid_186_1; // @[ICache.scala 52:22]
  reg  valid_187_0; // @[ICache.scala 52:22]
  reg  valid_187_1; // @[ICache.scala 52:22]
  reg  valid_188_0; // @[ICache.scala 52:22]
  reg  valid_188_1; // @[ICache.scala 52:22]
  reg  valid_189_0; // @[ICache.scala 52:22]
  reg  valid_189_1; // @[ICache.scala 52:22]
  reg  valid_190_0; // @[ICache.scala 52:22]
  reg  valid_190_1; // @[ICache.scala 52:22]
  reg  valid_191_0; // @[ICache.scala 52:22]
  reg  valid_191_1; // @[ICache.scala 52:22]
  reg  valid_192_0; // @[ICache.scala 52:22]
  reg  valid_192_1; // @[ICache.scala 52:22]
  reg  valid_193_0; // @[ICache.scala 52:22]
  reg  valid_193_1; // @[ICache.scala 52:22]
  reg  valid_194_0; // @[ICache.scala 52:22]
  reg  valid_194_1; // @[ICache.scala 52:22]
  reg  valid_195_0; // @[ICache.scala 52:22]
  reg  valid_195_1; // @[ICache.scala 52:22]
  reg  valid_196_0; // @[ICache.scala 52:22]
  reg  valid_196_1; // @[ICache.scala 52:22]
  reg  valid_197_0; // @[ICache.scala 52:22]
  reg  valid_197_1; // @[ICache.scala 52:22]
  reg  valid_198_0; // @[ICache.scala 52:22]
  reg  valid_198_1; // @[ICache.scala 52:22]
  reg  valid_199_0; // @[ICache.scala 52:22]
  reg  valid_199_1; // @[ICache.scala 52:22]
  reg  valid_200_0; // @[ICache.scala 52:22]
  reg  valid_200_1; // @[ICache.scala 52:22]
  reg  valid_201_0; // @[ICache.scala 52:22]
  reg  valid_201_1; // @[ICache.scala 52:22]
  reg  valid_202_0; // @[ICache.scala 52:22]
  reg  valid_202_1; // @[ICache.scala 52:22]
  reg  valid_203_0; // @[ICache.scala 52:22]
  reg  valid_203_1; // @[ICache.scala 52:22]
  reg  valid_204_0; // @[ICache.scala 52:22]
  reg  valid_204_1; // @[ICache.scala 52:22]
  reg  valid_205_0; // @[ICache.scala 52:22]
  reg  valid_205_1; // @[ICache.scala 52:22]
  reg  valid_206_0; // @[ICache.scala 52:22]
  reg  valid_206_1; // @[ICache.scala 52:22]
  reg  valid_207_0; // @[ICache.scala 52:22]
  reg  valid_207_1; // @[ICache.scala 52:22]
  reg  valid_208_0; // @[ICache.scala 52:22]
  reg  valid_208_1; // @[ICache.scala 52:22]
  reg  valid_209_0; // @[ICache.scala 52:22]
  reg  valid_209_1; // @[ICache.scala 52:22]
  reg  valid_210_0; // @[ICache.scala 52:22]
  reg  valid_210_1; // @[ICache.scala 52:22]
  reg  valid_211_0; // @[ICache.scala 52:22]
  reg  valid_211_1; // @[ICache.scala 52:22]
  reg  valid_212_0; // @[ICache.scala 52:22]
  reg  valid_212_1; // @[ICache.scala 52:22]
  reg  valid_213_0; // @[ICache.scala 52:22]
  reg  valid_213_1; // @[ICache.scala 52:22]
  reg  valid_214_0; // @[ICache.scala 52:22]
  reg  valid_214_1; // @[ICache.scala 52:22]
  reg  valid_215_0; // @[ICache.scala 52:22]
  reg  valid_215_1; // @[ICache.scala 52:22]
  reg  valid_216_0; // @[ICache.scala 52:22]
  reg  valid_216_1; // @[ICache.scala 52:22]
  reg  valid_217_0; // @[ICache.scala 52:22]
  reg  valid_217_1; // @[ICache.scala 52:22]
  reg  valid_218_0; // @[ICache.scala 52:22]
  reg  valid_218_1; // @[ICache.scala 52:22]
  reg  valid_219_0; // @[ICache.scala 52:22]
  reg  valid_219_1; // @[ICache.scala 52:22]
  reg  valid_220_0; // @[ICache.scala 52:22]
  reg  valid_220_1; // @[ICache.scala 52:22]
  reg  valid_221_0; // @[ICache.scala 52:22]
  reg  valid_221_1; // @[ICache.scala 52:22]
  reg  valid_222_0; // @[ICache.scala 52:22]
  reg  valid_222_1; // @[ICache.scala 52:22]
  reg  valid_223_0; // @[ICache.scala 52:22]
  reg  valid_223_1; // @[ICache.scala 52:22]
  reg  valid_224_0; // @[ICache.scala 52:22]
  reg  valid_224_1; // @[ICache.scala 52:22]
  reg  valid_225_0; // @[ICache.scala 52:22]
  reg  valid_225_1; // @[ICache.scala 52:22]
  reg  valid_226_0; // @[ICache.scala 52:22]
  reg  valid_226_1; // @[ICache.scala 52:22]
  reg  valid_227_0; // @[ICache.scala 52:22]
  reg  valid_227_1; // @[ICache.scala 52:22]
  reg  valid_228_0; // @[ICache.scala 52:22]
  reg  valid_228_1; // @[ICache.scala 52:22]
  reg  valid_229_0; // @[ICache.scala 52:22]
  reg  valid_229_1; // @[ICache.scala 52:22]
  reg  valid_230_0; // @[ICache.scala 52:22]
  reg  valid_230_1; // @[ICache.scala 52:22]
  reg  valid_231_0; // @[ICache.scala 52:22]
  reg  valid_231_1; // @[ICache.scala 52:22]
  reg  valid_232_0; // @[ICache.scala 52:22]
  reg  valid_232_1; // @[ICache.scala 52:22]
  reg  valid_233_0; // @[ICache.scala 52:22]
  reg  valid_233_1; // @[ICache.scala 52:22]
  reg  valid_234_0; // @[ICache.scala 52:22]
  reg  valid_234_1; // @[ICache.scala 52:22]
  reg  valid_235_0; // @[ICache.scala 52:22]
  reg  valid_235_1; // @[ICache.scala 52:22]
  reg  valid_236_0; // @[ICache.scala 52:22]
  reg  valid_236_1; // @[ICache.scala 52:22]
  reg  valid_237_0; // @[ICache.scala 52:22]
  reg  valid_237_1; // @[ICache.scala 52:22]
  reg  valid_238_0; // @[ICache.scala 52:22]
  reg  valid_238_1; // @[ICache.scala 52:22]
  reg  valid_239_0; // @[ICache.scala 52:22]
  reg  valid_239_1; // @[ICache.scala 52:22]
  reg  valid_240_0; // @[ICache.scala 52:22]
  reg  valid_240_1; // @[ICache.scala 52:22]
  reg  valid_241_0; // @[ICache.scala 52:22]
  reg  valid_241_1; // @[ICache.scala 52:22]
  reg  valid_242_0; // @[ICache.scala 52:22]
  reg  valid_242_1; // @[ICache.scala 52:22]
  reg  valid_243_0; // @[ICache.scala 52:22]
  reg  valid_243_1; // @[ICache.scala 52:22]
  reg  valid_244_0; // @[ICache.scala 52:22]
  reg  valid_244_1; // @[ICache.scala 52:22]
  reg  valid_245_0; // @[ICache.scala 52:22]
  reg  valid_245_1; // @[ICache.scala 52:22]
  reg  valid_246_0; // @[ICache.scala 52:22]
  reg  valid_246_1; // @[ICache.scala 52:22]
  reg  valid_247_0; // @[ICache.scala 52:22]
  reg  valid_247_1; // @[ICache.scala 52:22]
  reg  valid_248_0; // @[ICache.scala 52:22]
  reg  valid_248_1; // @[ICache.scala 52:22]
  reg  valid_249_0; // @[ICache.scala 52:22]
  reg  valid_249_1; // @[ICache.scala 52:22]
  reg  valid_250_0; // @[ICache.scala 52:22]
  reg  valid_250_1; // @[ICache.scala 52:22]
  reg  valid_251_0; // @[ICache.scala 52:22]
  reg  valid_251_1; // @[ICache.scala 52:22]
  reg  valid_252_0; // @[ICache.scala 52:22]
  reg  valid_252_1; // @[ICache.scala 52:22]
  reg  valid_253_0; // @[ICache.scala 52:22]
  reg  valid_253_1; // @[ICache.scala 52:22]
  reg  valid_254_0; // @[ICache.scala 52:22]
  reg  valid_254_1; // @[ICache.scala 52:22]
  reg  valid_255_0; // @[ICache.scala 52:22]
  reg  valid_255_1; // @[ICache.scala 52:22]
  reg  valid_256_0; // @[ICache.scala 52:22]
  reg  valid_256_1; // @[ICache.scala 52:22]
  reg  valid_257_0; // @[ICache.scala 52:22]
  reg  valid_257_1; // @[ICache.scala 52:22]
  reg  valid_258_0; // @[ICache.scala 52:22]
  reg  valid_258_1; // @[ICache.scala 52:22]
  reg  valid_259_0; // @[ICache.scala 52:22]
  reg  valid_259_1; // @[ICache.scala 52:22]
  reg  valid_260_0; // @[ICache.scala 52:22]
  reg  valid_260_1; // @[ICache.scala 52:22]
  reg  valid_261_0; // @[ICache.scala 52:22]
  reg  valid_261_1; // @[ICache.scala 52:22]
  reg  valid_262_0; // @[ICache.scala 52:22]
  reg  valid_262_1; // @[ICache.scala 52:22]
  reg  valid_263_0; // @[ICache.scala 52:22]
  reg  valid_263_1; // @[ICache.scala 52:22]
  reg  valid_264_0; // @[ICache.scala 52:22]
  reg  valid_264_1; // @[ICache.scala 52:22]
  reg  valid_265_0; // @[ICache.scala 52:22]
  reg  valid_265_1; // @[ICache.scala 52:22]
  reg  valid_266_0; // @[ICache.scala 52:22]
  reg  valid_266_1; // @[ICache.scala 52:22]
  reg  valid_267_0; // @[ICache.scala 52:22]
  reg  valid_267_1; // @[ICache.scala 52:22]
  reg  valid_268_0; // @[ICache.scala 52:22]
  reg  valid_268_1; // @[ICache.scala 52:22]
  reg  valid_269_0; // @[ICache.scala 52:22]
  reg  valid_269_1; // @[ICache.scala 52:22]
  reg  valid_270_0; // @[ICache.scala 52:22]
  reg  valid_270_1; // @[ICache.scala 52:22]
  reg  valid_271_0; // @[ICache.scala 52:22]
  reg  valid_271_1; // @[ICache.scala 52:22]
  reg  valid_272_0; // @[ICache.scala 52:22]
  reg  valid_272_1; // @[ICache.scala 52:22]
  reg  valid_273_0; // @[ICache.scala 52:22]
  reg  valid_273_1; // @[ICache.scala 52:22]
  reg  valid_274_0; // @[ICache.scala 52:22]
  reg  valid_274_1; // @[ICache.scala 52:22]
  reg  valid_275_0; // @[ICache.scala 52:22]
  reg  valid_275_1; // @[ICache.scala 52:22]
  reg  valid_276_0; // @[ICache.scala 52:22]
  reg  valid_276_1; // @[ICache.scala 52:22]
  reg  valid_277_0; // @[ICache.scala 52:22]
  reg  valid_277_1; // @[ICache.scala 52:22]
  reg  valid_278_0; // @[ICache.scala 52:22]
  reg  valid_278_1; // @[ICache.scala 52:22]
  reg  valid_279_0; // @[ICache.scala 52:22]
  reg  valid_279_1; // @[ICache.scala 52:22]
  reg  valid_280_0; // @[ICache.scala 52:22]
  reg  valid_280_1; // @[ICache.scala 52:22]
  reg  valid_281_0; // @[ICache.scala 52:22]
  reg  valid_281_1; // @[ICache.scala 52:22]
  reg  valid_282_0; // @[ICache.scala 52:22]
  reg  valid_282_1; // @[ICache.scala 52:22]
  reg  valid_283_0; // @[ICache.scala 52:22]
  reg  valid_283_1; // @[ICache.scala 52:22]
  reg  valid_284_0; // @[ICache.scala 52:22]
  reg  valid_284_1; // @[ICache.scala 52:22]
  reg  valid_285_0; // @[ICache.scala 52:22]
  reg  valid_285_1; // @[ICache.scala 52:22]
  reg  valid_286_0; // @[ICache.scala 52:22]
  reg  valid_286_1; // @[ICache.scala 52:22]
  reg  valid_287_0; // @[ICache.scala 52:22]
  reg  valid_287_1; // @[ICache.scala 52:22]
  reg  valid_288_0; // @[ICache.scala 52:22]
  reg  valid_288_1; // @[ICache.scala 52:22]
  reg  valid_289_0; // @[ICache.scala 52:22]
  reg  valid_289_1; // @[ICache.scala 52:22]
  reg  valid_290_0; // @[ICache.scala 52:22]
  reg  valid_290_1; // @[ICache.scala 52:22]
  reg  valid_291_0; // @[ICache.scala 52:22]
  reg  valid_291_1; // @[ICache.scala 52:22]
  reg  valid_292_0; // @[ICache.scala 52:22]
  reg  valid_292_1; // @[ICache.scala 52:22]
  reg  valid_293_0; // @[ICache.scala 52:22]
  reg  valid_293_1; // @[ICache.scala 52:22]
  reg  valid_294_0; // @[ICache.scala 52:22]
  reg  valid_294_1; // @[ICache.scala 52:22]
  reg  valid_295_0; // @[ICache.scala 52:22]
  reg  valid_295_1; // @[ICache.scala 52:22]
  reg  valid_296_0; // @[ICache.scala 52:22]
  reg  valid_296_1; // @[ICache.scala 52:22]
  reg  valid_297_0; // @[ICache.scala 52:22]
  reg  valid_297_1; // @[ICache.scala 52:22]
  reg  valid_298_0; // @[ICache.scala 52:22]
  reg  valid_298_1; // @[ICache.scala 52:22]
  reg  valid_299_0; // @[ICache.scala 52:22]
  reg  valid_299_1; // @[ICache.scala 52:22]
  reg  valid_300_0; // @[ICache.scala 52:22]
  reg  valid_300_1; // @[ICache.scala 52:22]
  reg  valid_301_0; // @[ICache.scala 52:22]
  reg  valid_301_1; // @[ICache.scala 52:22]
  reg  valid_302_0; // @[ICache.scala 52:22]
  reg  valid_302_1; // @[ICache.scala 52:22]
  reg  valid_303_0; // @[ICache.scala 52:22]
  reg  valid_303_1; // @[ICache.scala 52:22]
  reg  valid_304_0; // @[ICache.scala 52:22]
  reg  valid_304_1; // @[ICache.scala 52:22]
  reg  valid_305_0; // @[ICache.scala 52:22]
  reg  valid_305_1; // @[ICache.scala 52:22]
  reg  valid_306_0; // @[ICache.scala 52:22]
  reg  valid_306_1; // @[ICache.scala 52:22]
  reg  valid_307_0; // @[ICache.scala 52:22]
  reg  valid_307_1; // @[ICache.scala 52:22]
  reg  valid_308_0; // @[ICache.scala 52:22]
  reg  valid_308_1; // @[ICache.scala 52:22]
  reg  valid_309_0; // @[ICache.scala 52:22]
  reg  valid_309_1; // @[ICache.scala 52:22]
  reg  valid_310_0; // @[ICache.scala 52:22]
  reg  valid_310_1; // @[ICache.scala 52:22]
  reg  valid_311_0; // @[ICache.scala 52:22]
  reg  valid_311_1; // @[ICache.scala 52:22]
  reg  valid_312_0; // @[ICache.scala 52:22]
  reg  valid_312_1; // @[ICache.scala 52:22]
  reg  valid_313_0; // @[ICache.scala 52:22]
  reg  valid_313_1; // @[ICache.scala 52:22]
  reg  valid_314_0; // @[ICache.scala 52:22]
  reg  valid_314_1; // @[ICache.scala 52:22]
  reg  valid_315_0; // @[ICache.scala 52:22]
  reg  valid_315_1; // @[ICache.scala 52:22]
  reg  valid_316_0; // @[ICache.scala 52:22]
  reg  valid_316_1; // @[ICache.scala 52:22]
  reg  valid_317_0; // @[ICache.scala 52:22]
  reg  valid_317_1; // @[ICache.scala 52:22]
  reg  valid_318_0; // @[ICache.scala 52:22]
  reg  valid_318_1; // @[ICache.scala 52:22]
  reg  valid_319_0; // @[ICache.scala 52:22]
  reg  valid_319_1; // @[ICache.scala 52:22]
  reg  valid_320_0; // @[ICache.scala 52:22]
  reg  valid_320_1; // @[ICache.scala 52:22]
  reg  valid_321_0; // @[ICache.scala 52:22]
  reg  valid_321_1; // @[ICache.scala 52:22]
  reg  valid_322_0; // @[ICache.scala 52:22]
  reg  valid_322_1; // @[ICache.scala 52:22]
  reg  valid_323_0; // @[ICache.scala 52:22]
  reg  valid_323_1; // @[ICache.scala 52:22]
  reg  valid_324_0; // @[ICache.scala 52:22]
  reg  valid_324_1; // @[ICache.scala 52:22]
  reg  valid_325_0; // @[ICache.scala 52:22]
  reg  valid_325_1; // @[ICache.scala 52:22]
  reg  valid_326_0; // @[ICache.scala 52:22]
  reg  valid_326_1; // @[ICache.scala 52:22]
  reg  valid_327_0; // @[ICache.scala 52:22]
  reg  valid_327_1; // @[ICache.scala 52:22]
  reg  valid_328_0; // @[ICache.scala 52:22]
  reg  valid_328_1; // @[ICache.scala 52:22]
  reg  valid_329_0; // @[ICache.scala 52:22]
  reg  valid_329_1; // @[ICache.scala 52:22]
  reg  valid_330_0; // @[ICache.scala 52:22]
  reg  valid_330_1; // @[ICache.scala 52:22]
  reg  valid_331_0; // @[ICache.scala 52:22]
  reg  valid_331_1; // @[ICache.scala 52:22]
  reg  valid_332_0; // @[ICache.scala 52:22]
  reg  valid_332_1; // @[ICache.scala 52:22]
  reg  valid_333_0; // @[ICache.scala 52:22]
  reg  valid_333_1; // @[ICache.scala 52:22]
  reg  valid_334_0; // @[ICache.scala 52:22]
  reg  valid_334_1; // @[ICache.scala 52:22]
  reg  valid_335_0; // @[ICache.scala 52:22]
  reg  valid_335_1; // @[ICache.scala 52:22]
  reg  valid_336_0; // @[ICache.scala 52:22]
  reg  valid_336_1; // @[ICache.scala 52:22]
  reg  valid_337_0; // @[ICache.scala 52:22]
  reg  valid_337_1; // @[ICache.scala 52:22]
  reg  valid_338_0; // @[ICache.scala 52:22]
  reg  valid_338_1; // @[ICache.scala 52:22]
  reg  valid_339_0; // @[ICache.scala 52:22]
  reg  valid_339_1; // @[ICache.scala 52:22]
  reg  valid_340_0; // @[ICache.scala 52:22]
  reg  valid_340_1; // @[ICache.scala 52:22]
  reg  valid_341_0; // @[ICache.scala 52:22]
  reg  valid_341_1; // @[ICache.scala 52:22]
  reg  valid_342_0; // @[ICache.scala 52:22]
  reg  valid_342_1; // @[ICache.scala 52:22]
  reg  valid_343_0; // @[ICache.scala 52:22]
  reg  valid_343_1; // @[ICache.scala 52:22]
  reg  valid_344_0; // @[ICache.scala 52:22]
  reg  valid_344_1; // @[ICache.scala 52:22]
  reg  valid_345_0; // @[ICache.scala 52:22]
  reg  valid_345_1; // @[ICache.scala 52:22]
  reg  valid_346_0; // @[ICache.scala 52:22]
  reg  valid_346_1; // @[ICache.scala 52:22]
  reg  valid_347_0; // @[ICache.scala 52:22]
  reg  valid_347_1; // @[ICache.scala 52:22]
  reg  valid_348_0; // @[ICache.scala 52:22]
  reg  valid_348_1; // @[ICache.scala 52:22]
  reg  valid_349_0; // @[ICache.scala 52:22]
  reg  valid_349_1; // @[ICache.scala 52:22]
  reg  valid_350_0; // @[ICache.scala 52:22]
  reg  valid_350_1; // @[ICache.scala 52:22]
  reg  valid_351_0; // @[ICache.scala 52:22]
  reg  valid_351_1; // @[ICache.scala 52:22]
  reg  valid_352_0; // @[ICache.scala 52:22]
  reg  valid_352_1; // @[ICache.scala 52:22]
  reg  valid_353_0; // @[ICache.scala 52:22]
  reg  valid_353_1; // @[ICache.scala 52:22]
  reg  valid_354_0; // @[ICache.scala 52:22]
  reg  valid_354_1; // @[ICache.scala 52:22]
  reg  valid_355_0; // @[ICache.scala 52:22]
  reg  valid_355_1; // @[ICache.scala 52:22]
  reg  valid_356_0; // @[ICache.scala 52:22]
  reg  valid_356_1; // @[ICache.scala 52:22]
  reg  valid_357_0; // @[ICache.scala 52:22]
  reg  valid_357_1; // @[ICache.scala 52:22]
  reg  valid_358_0; // @[ICache.scala 52:22]
  reg  valid_358_1; // @[ICache.scala 52:22]
  reg  valid_359_0; // @[ICache.scala 52:22]
  reg  valid_359_1; // @[ICache.scala 52:22]
  reg  valid_360_0; // @[ICache.scala 52:22]
  reg  valid_360_1; // @[ICache.scala 52:22]
  reg  valid_361_0; // @[ICache.scala 52:22]
  reg  valid_361_1; // @[ICache.scala 52:22]
  reg  valid_362_0; // @[ICache.scala 52:22]
  reg  valid_362_1; // @[ICache.scala 52:22]
  reg  valid_363_0; // @[ICache.scala 52:22]
  reg  valid_363_1; // @[ICache.scala 52:22]
  reg  valid_364_0; // @[ICache.scala 52:22]
  reg  valid_364_1; // @[ICache.scala 52:22]
  reg  valid_365_0; // @[ICache.scala 52:22]
  reg  valid_365_1; // @[ICache.scala 52:22]
  reg  valid_366_0; // @[ICache.scala 52:22]
  reg  valid_366_1; // @[ICache.scala 52:22]
  reg  valid_367_0; // @[ICache.scala 52:22]
  reg  valid_367_1; // @[ICache.scala 52:22]
  reg  valid_368_0; // @[ICache.scala 52:22]
  reg  valid_368_1; // @[ICache.scala 52:22]
  reg  valid_369_0; // @[ICache.scala 52:22]
  reg  valid_369_1; // @[ICache.scala 52:22]
  reg  valid_370_0; // @[ICache.scala 52:22]
  reg  valid_370_1; // @[ICache.scala 52:22]
  reg  valid_371_0; // @[ICache.scala 52:22]
  reg  valid_371_1; // @[ICache.scala 52:22]
  reg  valid_372_0; // @[ICache.scala 52:22]
  reg  valid_372_1; // @[ICache.scala 52:22]
  reg  valid_373_0; // @[ICache.scala 52:22]
  reg  valid_373_1; // @[ICache.scala 52:22]
  reg  valid_374_0; // @[ICache.scala 52:22]
  reg  valid_374_1; // @[ICache.scala 52:22]
  reg  valid_375_0; // @[ICache.scala 52:22]
  reg  valid_375_1; // @[ICache.scala 52:22]
  reg  valid_376_0; // @[ICache.scala 52:22]
  reg  valid_376_1; // @[ICache.scala 52:22]
  reg  valid_377_0; // @[ICache.scala 52:22]
  reg  valid_377_1; // @[ICache.scala 52:22]
  reg  valid_378_0; // @[ICache.scala 52:22]
  reg  valid_378_1; // @[ICache.scala 52:22]
  reg  valid_379_0; // @[ICache.scala 52:22]
  reg  valid_379_1; // @[ICache.scala 52:22]
  reg  valid_380_0; // @[ICache.scala 52:22]
  reg  valid_380_1; // @[ICache.scala 52:22]
  reg  valid_381_0; // @[ICache.scala 52:22]
  reg  valid_381_1; // @[ICache.scala 52:22]
  reg  valid_382_0; // @[ICache.scala 52:22]
  reg  valid_382_1; // @[ICache.scala 52:22]
  reg  valid_383_0; // @[ICache.scala 52:22]
  reg  valid_383_1; // @[ICache.scala 52:22]
  reg  valid_384_0; // @[ICache.scala 52:22]
  reg  valid_384_1; // @[ICache.scala 52:22]
  reg  valid_385_0; // @[ICache.scala 52:22]
  reg  valid_385_1; // @[ICache.scala 52:22]
  reg  valid_386_0; // @[ICache.scala 52:22]
  reg  valid_386_1; // @[ICache.scala 52:22]
  reg  valid_387_0; // @[ICache.scala 52:22]
  reg  valid_387_1; // @[ICache.scala 52:22]
  reg  valid_388_0; // @[ICache.scala 52:22]
  reg  valid_388_1; // @[ICache.scala 52:22]
  reg  valid_389_0; // @[ICache.scala 52:22]
  reg  valid_389_1; // @[ICache.scala 52:22]
  reg  valid_390_0; // @[ICache.scala 52:22]
  reg  valid_390_1; // @[ICache.scala 52:22]
  reg  valid_391_0; // @[ICache.scala 52:22]
  reg  valid_391_1; // @[ICache.scala 52:22]
  reg  valid_392_0; // @[ICache.scala 52:22]
  reg  valid_392_1; // @[ICache.scala 52:22]
  reg  valid_393_0; // @[ICache.scala 52:22]
  reg  valid_393_1; // @[ICache.scala 52:22]
  reg  valid_394_0; // @[ICache.scala 52:22]
  reg  valid_394_1; // @[ICache.scala 52:22]
  reg  valid_395_0; // @[ICache.scala 52:22]
  reg  valid_395_1; // @[ICache.scala 52:22]
  reg  valid_396_0; // @[ICache.scala 52:22]
  reg  valid_396_1; // @[ICache.scala 52:22]
  reg  valid_397_0; // @[ICache.scala 52:22]
  reg  valid_397_1; // @[ICache.scala 52:22]
  reg  valid_398_0; // @[ICache.scala 52:22]
  reg  valid_398_1; // @[ICache.scala 52:22]
  reg  valid_399_0; // @[ICache.scala 52:22]
  reg  valid_399_1; // @[ICache.scala 52:22]
  reg  valid_400_0; // @[ICache.scala 52:22]
  reg  valid_400_1; // @[ICache.scala 52:22]
  reg  valid_401_0; // @[ICache.scala 52:22]
  reg  valid_401_1; // @[ICache.scala 52:22]
  reg  valid_402_0; // @[ICache.scala 52:22]
  reg  valid_402_1; // @[ICache.scala 52:22]
  reg  valid_403_0; // @[ICache.scala 52:22]
  reg  valid_403_1; // @[ICache.scala 52:22]
  reg  valid_404_0; // @[ICache.scala 52:22]
  reg  valid_404_1; // @[ICache.scala 52:22]
  reg  valid_405_0; // @[ICache.scala 52:22]
  reg  valid_405_1; // @[ICache.scala 52:22]
  reg  valid_406_0; // @[ICache.scala 52:22]
  reg  valid_406_1; // @[ICache.scala 52:22]
  reg  valid_407_0; // @[ICache.scala 52:22]
  reg  valid_407_1; // @[ICache.scala 52:22]
  reg  valid_408_0; // @[ICache.scala 52:22]
  reg  valid_408_1; // @[ICache.scala 52:22]
  reg  valid_409_0; // @[ICache.scala 52:22]
  reg  valid_409_1; // @[ICache.scala 52:22]
  reg  valid_410_0; // @[ICache.scala 52:22]
  reg  valid_410_1; // @[ICache.scala 52:22]
  reg  valid_411_0; // @[ICache.scala 52:22]
  reg  valid_411_1; // @[ICache.scala 52:22]
  reg  valid_412_0; // @[ICache.scala 52:22]
  reg  valid_412_1; // @[ICache.scala 52:22]
  reg  valid_413_0; // @[ICache.scala 52:22]
  reg  valid_413_1; // @[ICache.scala 52:22]
  reg  valid_414_0; // @[ICache.scala 52:22]
  reg  valid_414_1; // @[ICache.scala 52:22]
  reg  valid_415_0; // @[ICache.scala 52:22]
  reg  valid_415_1; // @[ICache.scala 52:22]
  reg  valid_416_0; // @[ICache.scala 52:22]
  reg  valid_416_1; // @[ICache.scala 52:22]
  reg  valid_417_0; // @[ICache.scala 52:22]
  reg  valid_417_1; // @[ICache.scala 52:22]
  reg  valid_418_0; // @[ICache.scala 52:22]
  reg  valid_418_1; // @[ICache.scala 52:22]
  reg  valid_419_0; // @[ICache.scala 52:22]
  reg  valid_419_1; // @[ICache.scala 52:22]
  reg  valid_420_0; // @[ICache.scala 52:22]
  reg  valid_420_1; // @[ICache.scala 52:22]
  reg  valid_421_0; // @[ICache.scala 52:22]
  reg  valid_421_1; // @[ICache.scala 52:22]
  reg  valid_422_0; // @[ICache.scala 52:22]
  reg  valid_422_1; // @[ICache.scala 52:22]
  reg  valid_423_0; // @[ICache.scala 52:22]
  reg  valid_423_1; // @[ICache.scala 52:22]
  reg  valid_424_0; // @[ICache.scala 52:22]
  reg  valid_424_1; // @[ICache.scala 52:22]
  reg  valid_425_0; // @[ICache.scala 52:22]
  reg  valid_425_1; // @[ICache.scala 52:22]
  reg  valid_426_0; // @[ICache.scala 52:22]
  reg  valid_426_1; // @[ICache.scala 52:22]
  reg  valid_427_0; // @[ICache.scala 52:22]
  reg  valid_427_1; // @[ICache.scala 52:22]
  reg  valid_428_0; // @[ICache.scala 52:22]
  reg  valid_428_1; // @[ICache.scala 52:22]
  reg  valid_429_0; // @[ICache.scala 52:22]
  reg  valid_429_1; // @[ICache.scala 52:22]
  reg  valid_430_0; // @[ICache.scala 52:22]
  reg  valid_430_1; // @[ICache.scala 52:22]
  reg  valid_431_0; // @[ICache.scala 52:22]
  reg  valid_431_1; // @[ICache.scala 52:22]
  reg  valid_432_0; // @[ICache.scala 52:22]
  reg  valid_432_1; // @[ICache.scala 52:22]
  reg  valid_433_0; // @[ICache.scala 52:22]
  reg  valid_433_1; // @[ICache.scala 52:22]
  reg  valid_434_0; // @[ICache.scala 52:22]
  reg  valid_434_1; // @[ICache.scala 52:22]
  reg  valid_435_0; // @[ICache.scala 52:22]
  reg  valid_435_1; // @[ICache.scala 52:22]
  reg  valid_436_0; // @[ICache.scala 52:22]
  reg  valid_436_1; // @[ICache.scala 52:22]
  reg  valid_437_0; // @[ICache.scala 52:22]
  reg  valid_437_1; // @[ICache.scala 52:22]
  reg  valid_438_0; // @[ICache.scala 52:22]
  reg  valid_438_1; // @[ICache.scala 52:22]
  reg  valid_439_0; // @[ICache.scala 52:22]
  reg  valid_439_1; // @[ICache.scala 52:22]
  reg  valid_440_0; // @[ICache.scala 52:22]
  reg  valid_440_1; // @[ICache.scala 52:22]
  reg  valid_441_0; // @[ICache.scala 52:22]
  reg  valid_441_1; // @[ICache.scala 52:22]
  reg  valid_442_0; // @[ICache.scala 52:22]
  reg  valid_442_1; // @[ICache.scala 52:22]
  reg  valid_443_0; // @[ICache.scala 52:22]
  reg  valid_443_1; // @[ICache.scala 52:22]
  reg  valid_444_0; // @[ICache.scala 52:22]
  reg  valid_444_1; // @[ICache.scala 52:22]
  reg  valid_445_0; // @[ICache.scala 52:22]
  reg  valid_445_1; // @[ICache.scala 52:22]
  reg  valid_446_0; // @[ICache.scala 52:22]
  reg  valid_446_1; // @[ICache.scala 52:22]
  reg  valid_447_0; // @[ICache.scala 52:22]
  reg  valid_447_1; // @[ICache.scala 52:22]
  reg  valid_448_0; // @[ICache.scala 52:22]
  reg  valid_448_1; // @[ICache.scala 52:22]
  reg  valid_449_0; // @[ICache.scala 52:22]
  reg  valid_449_1; // @[ICache.scala 52:22]
  reg  valid_450_0; // @[ICache.scala 52:22]
  reg  valid_450_1; // @[ICache.scala 52:22]
  reg  valid_451_0; // @[ICache.scala 52:22]
  reg  valid_451_1; // @[ICache.scala 52:22]
  reg  valid_452_0; // @[ICache.scala 52:22]
  reg  valid_452_1; // @[ICache.scala 52:22]
  reg  valid_453_0; // @[ICache.scala 52:22]
  reg  valid_453_1; // @[ICache.scala 52:22]
  reg  valid_454_0; // @[ICache.scala 52:22]
  reg  valid_454_1; // @[ICache.scala 52:22]
  reg  valid_455_0; // @[ICache.scala 52:22]
  reg  valid_455_1; // @[ICache.scala 52:22]
  reg  valid_456_0; // @[ICache.scala 52:22]
  reg  valid_456_1; // @[ICache.scala 52:22]
  reg  valid_457_0; // @[ICache.scala 52:22]
  reg  valid_457_1; // @[ICache.scala 52:22]
  reg  valid_458_0; // @[ICache.scala 52:22]
  reg  valid_458_1; // @[ICache.scala 52:22]
  reg  valid_459_0; // @[ICache.scala 52:22]
  reg  valid_459_1; // @[ICache.scala 52:22]
  reg  valid_460_0; // @[ICache.scala 52:22]
  reg  valid_460_1; // @[ICache.scala 52:22]
  reg  valid_461_0; // @[ICache.scala 52:22]
  reg  valid_461_1; // @[ICache.scala 52:22]
  reg  valid_462_0; // @[ICache.scala 52:22]
  reg  valid_462_1; // @[ICache.scala 52:22]
  reg  valid_463_0; // @[ICache.scala 52:22]
  reg  valid_463_1; // @[ICache.scala 52:22]
  reg  valid_464_0; // @[ICache.scala 52:22]
  reg  valid_464_1; // @[ICache.scala 52:22]
  reg  valid_465_0; // @[ICache.scala 52:22]
  reg  valid_465_1; // @[ICache.scala 52:22]
  reg  valid_466_0; // @[ICache.scala 52:22]
  reg  valid_466_1; // @[ICache.scala 52:22]
  reg  valid_467_0; // @[ICache.scala 52:22]
  reg  valid_467_1; // @[ICache.scala 52:22]
  reg  valid_468_0; // @[ICache.scala 52:22]
  reg  valid_468_1; // @[ICache.scala 52:22]
  reg  valid_469_0; // @[ICache.scala 52:22]
  reg  valid_469_1; // @[ICache.scala 52:22]
  reg  valid_470_0; // @[ICache.scala 52:22]
  reg  valid_470_1; // @[ICache.scala 52:22]
  reg  valid_471_0; // @[ICache.scala 52:22]
  reg  valid_471_1; // @[ICache.scala 52:22]
  reg  valid_472_0; // @[ICache.scala 52:22]
  reg  valid_472_1; // @[ICache.scala 52:22]
  reg  valid_473_0; // @[ICache.scala 52:22]
  reg  valid_473_1; // @[ICache.scala 52:22]
  reg  valid_474_0; // @[ICache.scala 52:22]
  reg  valid_474_1; // @[ICache.scala 52:22]
  reg  valid_475_0; // @[ICache.scala 52:22]
  reg  valid_475_1; // @[ICache.scala 52:22]
  reg  valid_476_0; // @[ICache.scala 52:22]
  reg  valid_476_1; // @[ICache.scala 52:22]
  reg  valid_477_0; // @[ICache.scala 52:22]
  reg  valid_477_1; // @[ICache.scala 52:22]
  reg  valid_478_0; // @[ICache.scala 52:22]
  reg  valid_478_1; // @[ICache.scala 52:22]
  reg  valid_479_0; // @[ICache.scala 52:22]
  reg  valid_479_1; // @[ICache.scala 52:22]
  reg  valid_480_0; // @[ICache.scala 52:22]
  reg  valid_480_1; // @[ICache.scala 52:22]
  reg  valid_481_0; // @[ICache.scala 52:22]
  reg  valid_481_1; // @[ICache.scala 52:22]
  reg  valid_482_0; // @[ICache.scala 52:22]
  reg  valid_482_1; // @[ICache.scala 52:22]
  reg  valid_483_0; // @[ICache.scala 52:22]
  reg  valid_483_1; // @[ICache.scala 52:22]
  reg  valid_484_0; // @[ICache.scala 52:22]
  reg  valid_484_1; // @[ICache.scala 52:22]
  reg  valid_485_0; // @[ICache.scala 52:22]
  reg  valid_485_1; // @[ICache.scala 52:22]
  reg  valid_486_0; // @[ICache.scala 52:22]
  reg  valid_486_1; // @[ICache.scala 52:22]
  reg  valid_487_0; // @[ICache.scala 52:22]
  reg  valid_487_1; // @[ICache.scala 52:22]
  reg  valid_488_0; // @[ICache.scala 52:22]
  reg  valid_488_1; // @[ICache.scala 52:22]
  reg  valid_489_0; // @[ICache.scala 52:22]
  reg  valid_489_1; // @[ICache.scala 52:22]
  reg  valid_490_0; // @[ICache.scala 52:22]
  reg  valid_490_1; // @[ICache.scala 52:22]
  reg  valid_491_0; // @[ICache.scala 52:22]
  reg  valid_491_1; // @[ICache.scala 52:22]
  reg  valid_492_0; // @[ICache.scala 52:22]
  reg  valid_492_1; // @[ICache.scala 52:22]
  reg  valid_493_0; // @[ICache.scala 52:22]
  reg  valid_493_1; // @[ICache.scala 52:22]
  reg  valid_494_0; // @[ICache.scala 52:22]
  reg  valid_494_1; // @[ICache.scala 52:22]
  reg  valid_495_0; // @[ICache.scala 52:22]
  reg  valid_495_1; // @[ICache.scala 52:22]
  reg  valid_496_0; // @[ICache.scala 52:22]
  reg  valid_496_1; // @[ICache.scala 52:22]
  reg  valid_497_0; // @[ICache.scala 52:22]
  reg  valid_497_1; // @[ICache.scala 52:22]
  reg  valid_498_0; // @[ICache.scala 52:22]
  reg  valid_498_1; // @[ICache.scala 52:22]
  reg  valid_499_0; // @[ICache.scala 52:22]
  reg  valid_499_1; // @[ICache.scala 52:22]
  reg  valid_500_0; // @[ICache.scala 52:22]
  reg  valid_500_1; // @[ICache.scala 52:22]
  reg  valid_501_0; // @[ICache.scala 52:22]
  reg  valid_501_1; // @[ICache.scala 52:22]
  reg  valid_502_0; // @[ICache.scala 52:22]
  reg  valid_502_1; // @[ICache.scala 52:22]
  reg  valid_503_0; // @[ICache.scala 52:22]
  reg  valid_503_1; // @[ICache.scala 52:22]
  reg  valid_504_0; // @[ICache.scala 52:22]
  reg  valid_504_1; // @[ICache.scala 52:22]
  reg  valid_505_0; // @[ICache.scala 52:22]
  reg  valid_505_1; // @[ICache.scala 52:22]
  reg  valid_506_0; // @[ICache.scala 52:22]
  reg  valid_506_1; // @[ICache.scala 52:22]
  reg  valid_507_0; // @[ICache.scala 52:22]
  reg  valid_507_1; // @[ICache.scala 52:22]
  reg  valid_508_0; // @[ICache.scala 52:22]
  reg  valid_508_1; // @[ICache.scala 52:22]
  reg  valid_509_0; // @[ICache.scala 52:22]
  reg  valid_509_1; // @[ICache.scala 52:22]
  reg  valid_510_0; // @[ICache.scala 52:22]
  reg  valid_510_1; // @[ICache.scala 52:22]
  reg  valid_511_0; // @[ICache.scala 52:22]
  reg  valid_511_1; // @[ICache.scala 52:22]
  wire  _should_next_addr_T = state == 3'h0; // @[ICache.scala 58:33]
  wire  should_next_addr = state == 3'h0 | state == 3'h4; // @[ICache.scala 58:45]
  wire [31:0] _GEN_1 = should_next_addr ? io_cpu_addr_1 : io_cpu_addr_0; // @[ICache.scala 60:{49,49}]
  reg [3:0] data_wstrb_0_0; // @[ICache.scala 61:27]
  reg [3:0] data_wstrb_0_1; // @[ICache.scala 61:27]
  reg [3:0] data_wstrb_1_0; // @[ICache.scala 61:27]
  reg [3:0] data_wstrb_1_1; // @[ICache.scala 61:27]
  reg  tag_wstrb_0; // @[ICache.scala 64:26]
  reg  tag_wstrb_1; // @[ICache.scala 64:26]
  reg [19:0] tag_wdata; // @[ICache.scala 65:26]
  reg  lru_0; // @[ICache.scala 68:20]
  reg  lru_1; // @[ICache.scala 68:20]
  reg  lru_2; // @[ICache.scala 68:20]
  reg  lru_3; // @[ICache.scala 68:20]
  reg  lru_4; // @[ICache.scala 68:20]
  reg  lru_5; // @[ICache.scala 68:20]
  reg  lru_6; // @[ICache.scala 68:20]
  reg  lru_7; // @[ICache.scala 68:20]
  reg  lru_8; // @[ICache.scala 68:20]
  reg  lru_9; // @[ICache.scala 68:20]
  reg  lru_10; // @[ICache.scala 68:20]
  reg  lru_11; // @[ICache.scala 68:20]
  reg  lru_12; // @[ICache.scala 68:20]
  reg  lru_13; // @[ICache.scala 68:20]
  reg  lru_14; // @[ICache.scala 68:20]
  reg  lru_15; // @[ICache.scala 68:20]
  reg  lru_16; // @[ICache.scala 68:20]
  reg  lru_17; // @[ICache.scala 68:20]
  reg  lru_18; // @[ICache.scala 68:20]
  reg  lru_19; // @[ICache.scala 68:20]
  reg  lru_20; // @[ICache.scala 68:20]
  reg  lru_21; // @[ICache.scala 68:20]
  reg  lru_22; // @[ICache.scala 68:20]
  reg  lru_23; // @[ICache.scala 68:20]
  reg  lru_24; // @[ICache.scala 68:20]
  reg  lru_25; // @[ICache.scala 68:20]
  reg  lru_26; // @[ICache.scala 68:20]
  reg  lru_27; // @[ICache.scala 68:20]
  reg  lru_28; // @[ICache.scala 68:20]
  reg  lru_29; // @[ICache.scala 68:20]
  reg  lru_30; // @[ICache.scala 68:20]
  reg  lru_31; // @[ICache.scala 68:20]
  reg  lru_32; // @[ICache.scala 68:20]
  reg  lru_33; // @[ICache.scala 68:20]
  reg  lru_34; // @[ICache.scala 68:20]
  reg  lru_35; // @[ICache.scala 68:20]
  reg  lru_36; // @[ICache.scala 68:20]
  reg  lru_37; // @[ICache.scala 68:20]
  reg  lru_38; // @[ICache.scala 68:20]
  reg  lru_39; // @[ICache.scala 68:20]
  reg  lru_40; // @[ICache.scala 68:20]
  reg  lru_41; // @[ICache.scala 68:20]
  reg  lru_42; // @[ICache.scala 68:20]
  reg  lru_43; // @[ICache.scala 68:20]
  reg  lru_44; // @[ICache.scala 68:20]
  reg  lru_45; // @[ICache.scala 68:20]
  reg  lru_46; // @[ICache.scala 68:20]
  reg  lru_47; // @[ICache.scala 68:20]
  reg  lru_48; // @[ICache.scala 68:20]
  reg  lru_49; // @[ICache.scala 68:20]
  reg  lru_50; // @[ICache.scala 68:20]
  reg  lru_51; // @[ICache.scala 68:20]
  reg  lru_52; // @[ICache.scala 68:20]
  reg  lru_53; // @[ICache.scala 68:20]
  reg  lru_54; // @[ICache.scala 68:20]
  reg  lru_55; // @[ICache.scala 68:20]
  reg  lru_56; // @[ICache.scala 68:20]
  reg  lru_57; // @[ICache.scala 68:20]
  reg  lru_58; // @[ICache.scala 68:20]
  reg  lru_59; // @[ICache.scala 68:20]
  reg  lru_60; // @[ICache.scala 68:20]
  reg  lru_61; // @[ICache.scala 68:20]
  reg  lru_62; // @[ICache.scala 68:20]
  reg  lru_63; // @[ICache.scala 68:20]
  reg  lru_64; // @[ICache.scala 68:20]
  reg  lru_65; // @[ICache.scala 68:20]
  reg  lru_66; // @[ICache.scala 68:20]
  reg  lru_67; // @[ICache.scala 68:20]
  reg  lru_68; // @[ICache.scala 68:20]
  reg  lru_69; // @[ICache.scala 68:20]
  reg  lru_70; // @[ICache.scala 68:20]
  reg  lru_71; // @[ICache.scala 68:20]
  reg  lru_72; // @[ICache.scala 68:20]
  reg  lru_73; // @[ICache.scala 68:20]
  reg  lru_74; // @[ICache.scala 68:20]
  reg  lru_75; // @[ICache.scala 68:20]
  reg  lru_76; // @[ICache.scala 68:20]
  reg  lru_77; // @[ICache.scala 68:20]
  reg  lru_78; // @[ICache.scala 68:20]
  reg  lru_79; // @[ICache.scala 68:20]
  reg  lru_80; // @[ICache.scala 68:20]
  reg  lru_81; // @[ICache.scala 68:20]
  reg  lru_82; // @[ICache.scala 68:20]
  reg  lru_83; // @[ICache.scala 68:20]
  reg  lru_84; // @[ICache.scala 68:20]
  reg  lru_85; // @[ICache.scala 68:20]
  reg  lru_86; // @[ICache.scala 68:20]
  reg  lru_87; // @[ICache.scala 68:20]
  reg  lru_88; // @[ICache.scala 68:20]
  reg  lru_89; // @[ICache.scala 68:20]
  reg  lru_90; // @[ICache.scala 68:20]
  reg  lru_91; // @[ICache.scala 68:20]
  reg  lru_92; // @[ICache.scala 68:20]
  reg  lru_93; // @[ICache.scala 68:20]
  reg  lru_94; // @[ICache.scala 68:20]
  reg  lru_95; // @[ICache.scala 68:20]
  reg  lru_96; // @[ICache.scala 68:20]
  reg  lru_97; // @[ICache.scala 68:20]
  reg  lru_98; // @[ICache.scala 68:20]
  reg  lru_99; // @[ICache.scala 68:20]
  reg  lru_100; // @[ICache.scala 68:20]
  reg  lru_101; // @[ICache.scala 68:20]
  reg  lru_102; // @[ICache.scala 68:20]
  reg  lru_103; // @[ICache.scala 68:20]
  reg  lru_104; // @[ICache.scala 68:20]
  reg  lru_105; // @[ICache.scala 68:20]
  reg  lru_106; // @[ICache.scala 68:20]
  reg  lru_107; // @[ICache.scala 68:20]
  reg  lru_108; // @[ICache.scala 68:20]
  reg  lru_109; // @[ICache.scala 68:20]
  reg  lru_110; // @[ICache.scala 68:20]
  reg  lru_111; // @[ICache.scala 68:20]
  reg  lru_112; // @[ICache.scala 68:20]
  reg  lru_113; // @[ICache.scala 68:20]
  reg  lru_114; // @[ICache.scala 68:20]
  reg  lru_115; // @[ICache.scala 68:20]
  reg  lru_116; // @[ICache.scala 68:20]
  reg  lru_117; // @[ICache.scala 68:20]
  reg  lru_118; // @[ICache.scala 68:20]
  reg  lru_119; // @[ICache.scala 68:20]
  reg  lru_120; // @[ICache.scala 68:20]
  reg  lru_121; // @[ICache.scala 68:20]
  reg  lru_122; // @[ICache.scala 68:20]
  reg  lru_123; // @[ICache.scala 68:20]
  reg  lru_124; // @[ICache.scala 68:20]
  reg  lru_125; // @[ICache.scala 68:20]
  reg  lru_126; // @[ICache.scala 68:20]
  reg  lru_127; // @[ICache.scala 68:20]
  reg  lru_128; // @[ICache.scala 68:20]
  reg  lru_129; // @[ICache.scala 68:20]
  reg  lru_130; // @[ICache.scala 68:20]
  reg  lru_131; // @[ICache.scala 68:20]
  reg  lru_132; // @[ICache.scala 68:20]
  reg  lru_133; // @[ICache.scala 68:20]
  reg  lru_134; // @[ICache.scala 68:20]
  reg  lru_135; // @[ICache.scala 68:20]
  reg  lru_136; // @[ICache.scala 68:20]
  reg  lru_137; // @[ICache.scala 68:20]
  reg  lru_138; // @[ICache.scala 68:20]
  reg  lru_139; // @[ICache.scala 68:20]
  reg  lru_140; // @[ICache.scala 68:20]
  reg  lru_141; // @[ICache.scala 68:20]
  reg  lru_142; // @[ICache.scala 68:20]
  reg  lru_143; // @[ICache.scala 68:20]
  reg  lru_144; // @[ICache.scala 68:20]
  reg  lru_145; // @[ICache.scala 68:20]
  reg  lru_146; // @[ICache.scala 68:20]
  reg  lru_147; // @[ICache.scala 68:20]
  reg  lru_148; // @[ICache.scala 68:20]
  reg  lru_149; // @[ICache.scala 68:20]
  reg  lru_150; // @[ICache.scala 68:20]
  reg  lru_151; // @[ICache.scala 68:20]
  reg  lru_152; // @[ICache.scala 68:20]
  reg  lru_153; // @[ICache.scala 68:20]
  reg  lru_154; // @[ICache.scala 68:20]
  reg  lru_155; // @[ICache.scala 68:20]
  reg  lru_156; // @[ICache.scala 68:20]
  reg  lru_157; // @[ICache.scala 68:20]
  reg  lru_158; // @[ICache.scala 68:20]
  reg  lru_159; // @[ICache.scala 68:20]
  reg  lru_160; // @[ICache.scala 68:20]
  reg  lru_161; // @[ICache.scala 68:20]
  reg  lru_162; // @[ICache.scala 68:20]
  reg  lru_163; // @[ICache.scala 68:20]
  reg  lru_164; // @[ICache.scala 68:20]
  reg  lru_165; // @[ICache.scala 68:20]
  reg  lru_166; // @[ICache.scala 68:20]
  reg  lru_167; // @[ICache.scala 68:20]
  reg  lru_168; // @[ICache.scala 68:20]
  reg  lru_169; // @[ICache.scala 68:20]
  reg  lru_170; // @[ICache.scala 68:20]
  reg  lru_171; // @[ICache.scala 68:20]
  reg  lru_172; // @[ICache.scala 68:20]
  reg  lru_173; // @[ICache.scala 68:20]
  reg  lru_174; // @[ICache.scala 68:20]
  reg  lru_175; // @[ICache.scala 68:20]
  reg  lru_176; // @[ICache.scala 68:20]
  reg  lru_177; // @[ICache.scala 68:20]
  reg  lru_178; // @[ICache.scala 68:20]
  reg  lru_179; // @[ICache.scala 68:20]
  reg  lru_180; // @[ICache.scala 68:20]
  reg  lru_181; // @[ICache.scala 68:20]
  reg  lru_182; // @[ICache.scala 68:20]
  reg  lru_183; // @[ICache.scala 68:20]
  reg  lru_184; // @[ICache.scala 68:20]
  reg  lru_185; // @[ICache.scala 68:20]
  reg  lru_186; // @[ICache.scala 68:20]
  reg  lru_187; // @[ICache.scala 68:20]
  reg  lru_188; // @[ICache.scala 68:20]
  reg  lru_189; // @[ICache.scala 68:20]
  reg  lru_190; // @[ICache.scala 68:20]
  reg  lru_191; // @[ICache.scala 68:20]
  reg  lru_192; // @[ICache.scala 68:20]
  reg  lru_193; // @[ICache.scala 68:20]
  reg  lru_194; // @[ICache.scala 68:20]
  reg  lru_195; // @[ICache.scala 68:20]
  reg  lru_196; // @[ICache.scala 68:20]
  reg  lru_197; // @[ICache.scala 68:20]
  reg  lru_198; // @[ICache.scala 68:20]
  reg  lru_199; // @[ICache.scala 68:20]
  reg  lru_200; // @[ICache.scala 68:20]
  reg  lru_201; // @[ICache.scala 68:20]
  reg  lru_202; // @[ICache.scala 68:20]
  reg  lru_203; // @[ICache.scala 68:20]
  reg  lru_204; // @[ICache.scala 68:20]
  reg  lru_205; // @[ICache.scala 68:20]
  reg  lru_206; // @[ICache.scala 68:20]
  reg  lru_207; // @[ICache.scala 68:20]
  reg  lru_208; // @[ICache.scala 68:20]
  reg  lru_209; // @[ICache.scala 68:20]
  reg  lru_210; // @[ICache.scala 68:20]
  reg  lru_211; // @[ICache.scala 68:20]
  reg  lru_212; // @[ICache.scala 68:20]
  reg  lru_213; // @[ICache.scala 68:20]
  reg  lru_214; // @[ICache.scala 68:20]
  reg  lru_215; // @[ICache.scala 68:20]
  reg  lru_216; // @[ICache.scala 68:20]
  reg  lru_217; // @[ICache.scala 68:20]
  reg  lru_218; // @[ICache.scala 68:20]
  reg  lru_219; // @[ICache.scala 68:20]
  reg  lru_220; // @[ICache.scala 68:20]
  reg  lru_221; // @[ICache.scala 68:20]
  reg  lru_222; // @[ICache.scala 68:20]
  reg  lru_223; // @[ICache.scala 68:20]
  reg  lru_224; // @[ICache.scala 68:20]
  reg  lru_225; // @[ICache.scala 68:20]
  reg  lru_226; // @[ICache.scala 68:20]
  reg  lru_227; // @[ICache.scala 68:20]
  reg  lru_228; // @[ICache.scala 68:20]
  reg  lru_229; // @[ICache.scala 68:20]
  reg  lru_230; // @[ICache.scala 68:20]
  reg  lru_231; // @[ICache.scala 68:20]
  reg  lru_232; // @[ICache.scala 68:20]
  reg  lru_233; // @[ICache.scala 68:20]
  reg  lru_234; // @[ICache.scala 68:20]
  reg  lru_235; // @[ICache.scala 68:20]
  reg  lru_236; // @[ICache.scala 68:20]
  reg  lru_237; // @[ICache.scala 68:20]
  reg  lru_238; // @[ICache.scala 68:20]
  reg  lru_239; // @[ICache.scala 68:20]
  reg  lru_240; // @[ICache.scala 68:20]
  reg  lru_241; // @[ICache.scala 68:20]
  reg  lru_242; // @[ICache.scala 68:20]
  reg  lru_243; // @[ICache.scala 68:20]
  reg  lru_244; // @[ICache.scala 68:20]
  reg  lru_245; // @[ICache.scala 68:20]
  reg  lru_246; // @[ICache.scala 68:20]
  reg  lru_247; // @[ICache.scala 68:20]
  reg  lru_248; // @[ICache.scala 68:20]
  reg  lru_249; // @[ICache.scala 68:20]
  reg  lru_250; // @[ICache.scala 68:20]
  reg  lru_251; // @[ICache.scala 68:20]
  reg  lru_252; // @[ICache.scala 68:20]
  reg  lru_253; // @[ICache.scala 68:20]
  reg  lru_254; // @[ICache.scala 68:20]
  reg  lru_255; // @[ICache.scala 68:20]
  reg  lru_256; // @[ICache.scala 68:20]
  reg  lru_257; // @[ICache.scala 68:20]
  reg  lru_258; // @[ICache.scala 68:20]
  reg  lru_259; // @[ICache.scala 68:20]
  reg  lru_260; // @[ICache.scala 68:20]
  reg  lru_261; // @[ICache.scala 68:20]
  reg  lru_262; // @[ICache.scala 68:20]
  reg  lru_263; // @[ICache.scala 68:20]
  reg  lru_264; // @[ICache.scala 68:20]
  reg  lru_265; // @[ICache.scala 68:20]
  reg  lru_266; // @[ICache.scala 68:20]
  reg  lru_267; // @[ICache.scala 68:20]
  reg  lru_268; // @[ICache.scala 68:20]
  reg  lru_269; // @[ICache.scala 68:20]
  reg  lru_270; // @[ICache.scala 68:20]
  reg  lru_271; // @[ICache.scala 68:20]
  reg  lru_272; // @[ICache.scala 68:20]
  reg  lru_273; // @[ICache.scala 68:20]
  reg  lru_274; // @[ICache.scala 68:20]
  reg  lru_275; // @[ICache.scala 68:20]
  reg  lru_276; // @[ICache.scala 68:20]
  reg  lru_277; // @[ICache.scala 68:20]
  reg  lru_278; // @[ICache.scala 68:20]
  reg  lru_279; // @[ICache.scala 68:20]
  reg  lru_280; // @[ICache.scala 68:20]
  reg  lru_281; // @[ICache.scala 68:20]
  reg  lru_282; // @[ICache.scala 68:20]
  reg  lru_283; // @[ICache.scala 68:20]
  reg  lru_284; // @[ICache.scala 68:20]
  reg  lru_285; // @[ICache.scala 68:20]
  reg  lru_286; // @[ICache.scala 68:20]
  reg  lru_287; // @[ICache.scala 68:20]
  reg  lru_288; // @[ICache.scala 68:20]
  reg  lru_289; // @[ICache.scala 68:20]
  reg  lru_290; // @[ICache.scala 68:20]
  reg  lru_291; // @[ICache.scala 68:20]
  reg  lru_292; // @[ICache.scala 68:20]
  reg  lru_293; // @[ICache.scala 68:20]
  reg  lru_294; // @[ICache.scala 68:20]
  reg  lru_295; // @[ICache.scala 68:20]
  reg  lru_296; // @[ICache.scala 68:20]
  reg  lru_297; // @[ICache.scala 68:20]
  reg  lru_298; // @[ICache.scala 68:20]
  reg  lru_299; // @[ICache.scala 68:20]
  reg  lru_300; // @[ICache.scala 68:20]
  reg  lru_301; // @[ICache.scala 68:20]
  reg  lru_302; // @[ICache.scala 68:20]
  reg  lru_303; // @[ICache.scala 68:20]
  reg  lru_304; // @[ICache.scala 68:20]
  reg  lru_305; // @[ICache.scala 68:20]
  reg  lru_306; // @[ICache.scala 68:20]
  reg  lru_307; // @[ICache.scala 68:20]
  reg  lru_308; // @[ICache.scala 68:20]
  reg  lru_309; // @[ICache.scala 68:20]
  reg  lru_310; // @[ICache.scala 68:20]
  reg  lru_311; // @[ICache.scala 68:20]
  reg  lru_312; // @[ICache.scala 68:20]
  reg  lru_313; // @[ICache.scala 68:20]
  reg  lru_314; // @[ICache.scala 68:20]
  reg  lru_315; // @[ICache.scala 68:20]
  reg  lru_316; // @[ICache.scala 68:20]
  reg  lru_317; // @[ICache.scala 68:20]
  reg  lru_318; // @[ICache.scala 68:20]
  reg  lru_319; // @[ICache.scala 68:20]
  reg  lru_320; // @[ICache.scala 68:20]
  reg  lru_321; // @[ICache.scala 68:20]
  reg  lru_322; // @[ICache.scala 68:20]
  reg  lru_323; // @[ICache.scala 68:20]
  reg  lru_324; // @[ICache.scala 68:20]
  reg  lru_325; // @[ICache.scala 68:20]
  reg  lru_326; // @[ICache.scala 68:20]
  reg  lru_327; // @[ICache.scala 68:20]
  reg  lru_328; // @[ICache.scala 68:20]
  reg  lru_329; // @[ICache.scala 68:20]
  reg  lru_330; // @[ICache.scala 68:20]
  reg  lru_331; // @[ICache.scala 68:20]
  reg  lru_332; // @[ICache.scala 68:20]
  reg  lru_333; // @[ICache.scala 68:20]
  reg  lru_334; // @[ICache.scala 68:20]
  reg  lru_335; // @[ICache.scala 68:20]
  reg  lru_336; // @[ICache.scala 68:20]
  reg  lru_337; // @[ICache.scala 68:20]
  reg  lru_338; // @[ICache.scala 68:20]
  reg  lru_339; // @[ICache.scala 68:20]
  reg  lru_340; // @[ICache.scala 68:20]
  reg  lru_341; // @[ICache.scala 68:20]
  reg  lru_342; // @[ICache.scala 68:20]
  reg  lru_343; // @[ICache.scala 68:20]
  reg  lru_344; // @[ICache.scala 68:20]
  reg  lru_345; // @[ICache.scala 68:20]
  reg  lru_346; // @[ICache.scala 68:20]
  reg  lru_347; // @[ICache.scala 68:20]
  reg  lru_348; // @[ICache.scala 68:20]
  reg  lru_349; // @[ICache.scala 68:20]
  reg  lru_350; // @[ICache.scala 68:20]
  reg  lru_351; // @[ICache.scala 68:20]
  reg  lru_352; // @[ICache.scala 68:20]
  reg  lru_353; // @[ICache.scala 68:20]
  reg  lru_354; // @[ICache.scala 68:20]
  reg  lru_355; // @[ICache.scala 68:20]
  reg  lru_356; // @[ICache.scala 68:20]
  reg  lru_357; // @[ICache.scala 68:20]
  reg  lru_358; // @[ICache.scala 68:20]
  reg  lru_359; // @[ICache.scala 68:20]
  reg  lru_360; // @[ICache.scala 68:20]
  reg  lru_361; // @[ICache.scala 68:20]
  reg  lru_362; // @[ICache.scala 68:20]
  reg  lru_363; // @[ICache.scala 68:20]
  reg  lru_364; // @[ICache.scala 68:20]
  reg  lru_365; // @[ICache.scala 68:20]
  reg  lru_366; // @[ICache.scala 68:20]
  reg  lru_367; // @[ICache.scala 68:20]
  reg  lru_368; // @[ICache.scala 68:20]
  reg  lru_369; // @[ICache.scala 68:20]
  reg  lru_370; // @[ICache.scala 68:20]
  reg  lru_371; // @[ICache.scala 68:20]
  reg  lru_372; // @[ICache.scala 68:20]
  reg  lru_373; // @[ICache.scala 68:20]
  reg  lru_374; // @[ICache.scala 68:20]
  reg  lru_375; // @[ICache.scala 68:20]
  reg  lru_376; // @[ICache.scala 68:20]
  reg  lru_377; // @[ICache.scala 68:20]
  reg  lru_378; // @[ICache.scala 68:20]
  reg  lru_379; // @[ICache.scala 68:20]
  reg  lru_380; // @[ICache.scala 68:20]
  reg  lru_381; // @[ICache.scala 68:20]
  reg  lru_382; // @[ICache.scala 68:20]
  reg  lru_383; // @[ICache.scala 68:20]
  reg  lru_384; // @[ICache.scala 68:20]
  reg  lru_385; // @[ICache.scala 68:20]
  reg  lru_386; // @[ICache.scala 68:20]
  reg  lru_387; // @[ICache.scala 68:20]
  reg  lru_388; // @[ICache.scala 68:20]
  reg  lru_389; // @[ICache.scala 68:20]
  reg  lru_390; // @[ICache.scala 68:20]
  reg  lru_391; // @[ICache.scala 68:20]
  reg  lru_392; // @[ICache.scala 68:20]
  reg  lru_393; // @[ICache.scala 68:20]
  reg  lru_394; // @[ICache.scala 68:20]
  reg  lru_395; // @[ICache.scala 68:20]
  reg  lru_396; // @[ICache.scala 68:20]
  reg  lru_397; // @[ICache.scala 68:20]
  reg  lru_398; // @[ICache.scala 68:20]
  reg  lru_399; // @[ICache.scala 68:20]
  reg  lru_400; // @[ICache.scala 68:20]
  reg  lru_401; // @[ICache.scala 68:20]
  reg  lru_402; // @[ICache.scala 68:20]
  reg  lru_403; // @[ICache.scala 68:20]
  reg  lru_404; // @[ICache.scala 68:20]
  reg  lru_405; // @[ICache.scala 68:20]
  reg  lru_406; // @[ICache.scala 68:20]
  reg  lru_407; // @[ICache.scala 68:20]
  reg  lru_408; // @[ICache.scala 68:20]
  reg  lru_409; // @[ICache.scala 68:20]
  reg  lru_410; // @[ICache.scala 68:20]
  reg  lru_411; // @[ICache.scala 68:20]
  reg  lru_412; // @[ICache.scala 68:20]
  reg  lru_413; // @[ICache.scala 68:20]
  reg  lru_414; // @[ICache.scala 68:20]
  reg  lru_415; // @[ICache.scala 68:20]
  reg  lru_416; // @[ICache.scala 68:20]
  reg  lru_417; // @[ICache.scala 68:20]
  reg  lru_418; // @[ICache.scala 68:20]
  reg  lru_419; // @[ICache.scala 68:20]
  reg  lru_420; // @[ICache.scala 68:20]
  reg  lru_421; // @[ICache.scala 68:20]
  reg  lru_422; // @[ICache.scala 68:20]
  reg  lru_423; // @[ICache.scala 68:20]
  reg  lru_424; // @[ICache.scala 68:20]
  reg  lru_425; // @[ICache.scala 68:20]
  reg  lru_426; // @[ICache.scala 68:20]
  reg  lru_427; // @[ICache.scala 68:20]
  reg  lru_428; // @[ICache.scala 68:20]
  reg  lru_429; // @[ICache.scala 68:20]
  reg  lru_430; // @[ICache.scala 68:20]
  reg  lru_431; // @[ICache.scala 68:20]
  reg  lru_432; // @[ICache.scala 68:20]
  reg  lru_433; // @[ICache.scala 68:20]
  reg  lru_434; // @[ICache.scala 68:20]
  reg  lru_435; // @[ICache.scala 68:20]
  reg  lru_436; // @[ICache.scala 68:20]
  reg  lru_437; // @[ICache.scala 68:20]
  reg  lru_438; // @[ICache.scala 68:20]
  reg  lru_439; // @[ICache.scala 68:20]
  reg  lru_440; // @[ICache.scala 68:20]
  reg  lru_441; // @[ICache.scala 68:20]
  reg  lru_442; // @[ICache.scala 68:20]
  reg  lru_443; // @[ICache.scala 68:20]
  reg  lru_444; // @[ICache.scala 68:20]
  reg  lru_445; // @[ICache.scala 68:20]
  reg  lru_446; // @[ICache.scala 68:20]
  reg  lru_447; // @[ICache.scala 68:20]
  reg  lru_448; // @[ICache.scala 68:20]
  reg  lru_449; // @[ICache.scala 68:20]
  reg  lru_450; // @[ICache.scala 68:20]
  reg  lru_451; // @[ICache.scala 68:20]
  reg  lru_452; // @[ICache.scala 68:20]
  reg  lru_453; // @[ICache.scala 68:20]
  reg  lru_454; // @[ICache.scala 68:20]
  reg  lru_455; // @[ICache.scala 68:20]
  reg  lru_456; // @[ICache.scala 68:20]
  reg  lru_457; // @[ICache.scala 68:20]
  reg  lru_458; // @[ICache.scala 68:20]
  reg  lru_459; // @[ICache.scala 68:20]
  reg  lru_460; // @[ICache.scala 68:20]
  reg  lru_461; // @[ICache.scala 68:20]
  reg  lru_462; // @[ICache.scala 68:20]
  reg  lru_463; // @[ICache.scala 68:20]
  reg  lru_464; // @[ICache.scala 68:20]
  reg  lru_465; // @[ICache.scala 68:20]
  reg  lru_466; // @[ICache.scala 68:20]
  reg  lru_467; // @[ICache.scala 68:20]
  reg  lru_468; // @[ICache.scala 68:20]
  reg  lru_469; // @[ICache.scala 68:20]
  reg  lru_470; // @[ICache.scala 68:20]
  reg  lru_471; // @[ICache.scala 68:20]
  reg  lru_472; // @[ICache.scala 68:20]
  reg  lru_473; // @[ICache.scala 68:20]
  reg  lru_474; // @[ICache.scala 68:20]
  reg  lru_475; // @[ICache.scala 68:20]
  reg  lru_476; // @[ICache.scala 68:20]
  reg  lru_477; // @[ICache.scala 68:20]
  reg  lru_478; // @[ICache.scala 68:20]
  reg  lru_479; // @[ICache.scala 68:20]
  reg  lru_480; // @[ICache.scala 68:20]
  reg  lru_481; // @[ICache.scala 68:20]
  reg  lru_482; // @[ICache.scala 68:20]
  reg  lru_483; // @[ICache.scala 68:20]
  reg  lru_484; // @[ICache.scala 68:20]
  reg  lru_485; // @[ICache.scala 68:20]
  reg  lru_486; // @[ICache.scala 68:20]
  reg  lru_487; // @[ICache.scala 68:20]
  reg  lru_488; // @[ICache.scala 68:20]
  reg  lru_489; // @[ICache.scala 68:20]
  reg  lru_490; // @[ICache.scala 68:20]
  reg  lru_491; // @[ICache.scala 68:20]
  reg  lru_492; // @[ICache.scala 68:20]
  reg  lru_493; // @[ICache.scala 68:20]
  reg  lru_494; // @[ICache.scala 68:20]
  reg  lru_495; // @[ICache.scala 68:20]
  reg  lru_496; // @[ICache.scala 68:20]
  reg  lru_497; // @[ICache.scala 68:20]
  reg  lru_498; // @[ICache.scala 68:20]
  reg  lru_499; // @[ICache.scala 68:20]
  reg  lru_500; // @[ICache.scala 68:20]
  reg  lru_501; // @[ICache.scala 68:20]
  reg  lru_502; // @[ICache.scala 68:20]
  reg  lru_503; // @[ICache.scala 68:20]
  reg  lru_504; // @[ICache.scala 68:20]
  reg  lru_505; // @[ICache.scala 68:20]
  reg  lru_506; // @[ICache.scala 68:20]
  reg  lru_507; // @[ICache.scala 68:20]
  reg  lru_508; // @[ICache.scala 68:20]
  reg  lru_509; // @[ICache.scala 68:20]
  reg  lru_510; // @[ICache.scala 68:20]
  reg  lru_511; // @[ICache.scala 68:20]
  reg [19:0] tlb_vpn; // @[ICache.scala 71:20]
  reg [19:0] tlb_ppn; // @[ICache.scala 71:20]
  reg  tlb_uncached; // @[ICache.scala 71:20]
  reg  tlb_valid; // @[ICache.scala 71:20]
  wire  direct_mapped = io_cpu_addr_0[31:30] == 2'h2; // @[ICache.scala 79:46]
  wire  uncached = direct_mapped ? io_cpu_addr_0[29] : tlb_uncached; // @[ICache.scala 80:26]
  wire [19:0] _inst_tag_T_1 = {3'h0,io_cpu_addr_0[28:12]}; // @[Cat.scala 33:92]
  wire [19:0] inst_tag = direct_mapped ? _inst_tag_T_1 : tlb_ppn; // @[ICache.scala 81:26]
  wire [19:0] inst_vpn = io_cpu_addr_0[31:12]; // @[ICache.scala 82:37]
  wire [31:0] inst_pa = {inst_tag,io_cpu_addr_0[11:0]}; // @[Cat.scala 33:92]
  wire [5:0] fence_index = io_cpu_fence_addr[11:6]; // @[ICache.scala 86:38]
  wire  _T = ~io_cpu_icache_stall; // @[ICache.scala 87:28]
  wire  _T_2 = ~io_cpu_cpu_stall; // @[ICache.scala 87:52]
  wire  _GEN_2 = io_cpu_fence_tlb & ~io_cpu_icache_stall & ~io_cpu_cpu_stall ? 1'h0 : tlb_valid; // @[ICache.scala 71:20 87:{71,83}]
  wire  _GEN_3 = 6'h0 == fence_index ? 1'h0 : valid_0_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_4 = 6'h1 == fence_index ? 1'h0 : valid_1_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_5 = 6'h2 == fence_index ? 1'h0 : valid_2_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_6 = 6'h3 == fence_index ? 1'h0 : valid_3_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_7 = 6'h4 == fence_index ? 1'h0 : valid_4_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_8 = 6'h5 == fence_index ? 1'h0 : valid_5_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_9 = 6'h6 == fence_index ? 1'h0 : valid_6_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_10 = 6'h7 == fence_index ? 1'h0 : valid_7_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_11 = 6'h8 == fence_index ? 1'h0 : valid_8_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_12 = 6'h9 == fence_index ? 1'h0 : valid_9_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_13 = 6'ha == fence_index ? 1'h0 : valid_10_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_14 = 6'hb == fence_index ? 1'h0 : valid_11_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_15 = 6'hc == fence_index ? 1'h0 : valid_12_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_16 = 6'hd == fence_index ? 1'h0 : valid_13_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_17 = 6'he == fence_index ? 1'h0 : valid_14_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_18 = 6'hf == fence_index ? 1'h0 : valid_15_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_19 = 6'h10 == fence_index ? 1'h0 : valid_16_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_20 = 6'h11 == fence_index ? 1'h0 : valid_17_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_21 = 6'h12 == fence_index ? 1'h0 : valid_18_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_22 = 6'h13 == fence_index ? 1'h0 : valid_19_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_23 = 6'h14 == fence_index ? 1'h0 : valid_20_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_24 = 6'h15 == fence_index ? 1'h0 : valid_21_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_25 = 6'h16 == fence_index ? 1'h0 : valid_22_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_26 = 6'h17 == fence_index ? 1'h0 : valid_23_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_27 = 6'h18 == fence_index ? 1'h0 : valid_24_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_28 = 6'h19 == fence_index ? 1'h0 : valid_25_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_29 = 6'h1a == fence_index ? 1'h0 : valid_26_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_30 = 6'h1b == fence_index ? 1'h0 : valid_27_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_31 = 6'h1c == fence_index ? 1'h0 : valid_28_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_32 = 6'h1d == fence_index ? 1'h0 : valid_29_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_33 = 6'h1e == fence_index ? 1'h0 : valid_30_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_34 = 6'h1f == fence_index ? 1'h0 : valid_31_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_35 = 6'h20 == fence_index ? 1'h0 : valid_32_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_36 = 6'h21 == fence_index ? 1'h0 : valid_33_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_37 = 6'h22 == fence_index ? 1'h0 : valid_34_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_38 = 6'h23 == fence_index ? 1'h0 : valid_35_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_39 = 6'h24 == fence_index ? 1'h0 : valid_36_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_40 = 6'h25 == fence_index ? 1'h0 : valid_37_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_41 = 6'h26 == fence_index ? 1'h0 : valid_38_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_42 = 6'h27 == fence_index ? 1'h0 : valid_39_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_43 = 6'h28 == fence_index ? 1'h0 : valid_40_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_44 = 6'h29 == fence_index ? 1'h0 : valid_41_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_45 = 6'h2a == fence_index ? 1'h0 : valid_42_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_46 = 6'h2b == fence_index ? 1'h0 : valid_43_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_47 = 6'h2c == fence_index ? 1'h0 : valid_44_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_48 = 6'h2d == fence_index ? 1'h0 : valid_45_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_49 = 6'h2e == fence_index ? 1'h0 : valid_46_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_50 = 6'h2f == fence_index ? 1'h0 : valid_47_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_51 = 6'h30 == fence_index ? 1'h0 : valid_48_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_52 = 6'h31 == fence_index ? 1'h0 : valid_49_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_53 = 6'h32 == fence_index ? 1'h0 : valid_50_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_54 = 6'h33 == fence_index ? 1'h0 : valid_51_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_55 = 6'h34 == fence_index ? 1'h0 : valid_52_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_56 = 6'h35 == fence_index ? 1'h0 : valid_53_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_57 = 6'h36 == fence_index ? 1'h0 : valid_54_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_58 = 6'h37 == fence_index ? 1'h0 : valid_55_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_59 = 6'h38 == fence_index ? 1'h0 : valid_56_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_60 = 6'h39 == fence_index ? 1'h0 : valid_57_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_61 = 6'h3a == fence_index ? 1'h0 : valid_58_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_62 = 6'h3b == fence_index ? 1'h0 : valid_59_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_63 = 6'h3c == fence_index ? 1'h0 : valid_60_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_64 = 6'h3d == fence_index ? 1'h0 : valid_61_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_65 = 6'h3e == fence_index ? 1'h0 : valid_62_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_66 = 6'h3f == fence_index ? 1'h0 : valid_63_0; // @[ICache.scala 52:22 89:{24,24}]
  wire [6:0] _GEN_13543 = {{1'd0}, fence_index}; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_67 = 7'h40 == _GEN_13543 ? 1'h0 : valid_64_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_68 = 7'h41 == _GEN_13543 ? 1'h0 : valid_65_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_69 = 7'h42 == _GEN_13543 ? 1'h0 : valid_66_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_70 = 7'h43 == _GEN_13543 ? 1'h0 : valid_67_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_71 = 7'h44 == _GEN_13543 ? 1'h0 : valid_68_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_72 = 7'h45 == _GEN_13543 ? 1'h0 : valid_69_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_73 = 7'h46 == _GEN_13543 ? 1'h0 : valid_70_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_74 = 7'h47 == _GEN_13543 ? 1'h0 : valid_71_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_75 = 7'h48 == _GEN_13543 ? 1'h0 : valid_72_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_76 = 7'h49 == _GEN_13543 ? 1'h0 : valid_73_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_77 = 7'h4a == _GEN_13543 ? 1'h0 : valid_74_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_78 = 7'h4b == _GEN_13543 ? 1'h0 : valid_75_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_79 = 7'h4c == _GEN_13543 ? 1'h0 : valid_76_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_80 = 7'h4d == _GEN_13543 ? 1'h0 : valid_77_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_81 = 7'h4e == _GEN_13543 ? 1'h0 : valid_78_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_82 = 7'h4f == _GEN_13543 ? 1'h0 : valid_79_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_83 = 7'h50 == _GEN_13543 ? 1'h0 : valid_80_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_84 = 7'h51 == _GEN_13543 ? 1'h0 : valid_81_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_85 = 7'h52 == _GEN_13543 ? 1'h0 : valid_82_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_86 = 7'h53 == _GEN_13543 ? 1'h0 : valid_83_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_87 = 7'h54 == _GEN_13543 ? 1'h0 : valid_84_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_88 = 7'h55 == _GEN_13543 ? 1'h0 : valid_85_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_89 = 7'h56 == _GEN_13543 ? 1'h0 : valid_86_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_90 = 7'h57 == _GEN_13543 ? 1'h0 : valid_87_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_91 = 7'h58 == _GEN_13543 ? 1'h0 : valid_88_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_92 = 7'h59 == _GEN_13543 ? 1'h0 : valid_89_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_93 = 7'h5a == _GEN_13543 ? 1'h0 : valid_90_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_94 = 7'h5b == _GEN_13543 ? 1'h0 : valid_91_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_95 = 7'h5c == _GEN_13543 ? 1'h0 : valid_92_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_96 = 7'h5d == _GEN_13543 ? 1'h0 : valid_93_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_97 = 7'h5e == _GEN_13543 ? 1'h0 : valid_94_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_98 = 7'h5f == _GEN_13543 ? 1'h0 : valid_95_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_99 = 7'h60 == _GEN_13543 ? 1'h0 : valid_96_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_100 = 7'h61 == _GEN_13543 ? 1'h0 : valid_97_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_101 = 7'h62 == _GEN_13543 ? 1'h0 : valid_98_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_102 = 7'h63 == _GEN_13543 ? 1'h0 : valid_99_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_103 = 7'h64 == _GEN_13543 ? 1'h0 : valid_100_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_104 = 7'h65 == _GEN_13543 ? 1'h0 : valid_101_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_105 = 7'h66 == _GEN_13543 ? 1'h0 : valid_102_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_106 = 7'h67 == _GEN_13543 ? 1'h0 : valid_103_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_107 = 7'h68 == _GEN_13543 ? 1'h0 : valid_104_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_108 = 7'h69 == _GEN_13543 ? 1'h0 : valid_105_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_109 = 7'h6a == _GEN_13543 ? 1'h0 : valid_106_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_110 = 7'h6b == _GEN_13543 ? 1'h0 : valid_107_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_111 = 7'h6c == _GEN_13543 ? 1'h0 : valid_108_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_112 = 7'h6d == _GEN_13543 ? 1'h0 : valid_109_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_113 = 7'h6e == _GEN_13543 ? 1'h0 : valid_110_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_114 = 7'h6f == _GEN_13543 ? 1'h0 : valid_111_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_115 = 7'h70 == _GEN_13543 ? 1'h0 : valid_112_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_116 = 7'h71 == _GEN_13543 ? 1'h0 : valid_113_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_117 = 7'h72 == _GEN_13543 ? 1'h0 : valid_114_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_118 = 7'h73 == _GEN_13543 ? 1'h0 : valid_115_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_119 = 7'h74 == _GEN_13543 ? 1'h0 : valid_116_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_120 = 7'h75 == _GEN_13543 ? 1'h0 : valid_117_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_121 = 7'h76 == _GEN_13543 ? 1'h0 : valid_118_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_122 = 7'h77 == _GEN_13543 ? 1'h0 : valid_119_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_123 = 7'h78 == _GEN_13543 ? 1'h0 : valid_120_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_124 = 7'h79 == _GEN_13543 ? 1'h0 : valid_121_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_125 = 7'h7a == _GEN_13543 ? 1'h0 : valid_122_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_126 = 7'h7b == _GEN_13543 ? 1'h0 : valid_123_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_127 = 7'h7c == _GEN_13543 ? 1'h0 : valid_124_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_128 = 7'h7d == _GEN_13543 ? 1'h0 : valid_125_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_129 = 7'h7e == _GEN_13543 ? 1'h0 : valid_126_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_130 = 7'h7f == _GEN_13543 ? 1'h0 : valid_127_0; // @[ICache.scala 52:22 89:{24,24}]
  wire [7:0] _GEN_13607 = {{2'd0}, fence_index}; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_131 = 8'h80 == _GEN_13607 ? 1'h0 : valid_128_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_132 = 8'h81 == _GEN_13607 ? 1'h0 : valid_129_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_133 = 8'h82 == _GEN_13607 ? 1'h0 : valid_130_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_134 = 8'h83 == _GEN_13607 ? 1'h0 : valid_131_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_135 = 8'h84 == _GEN_13607 ? 1'h0 : valid_132_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_136 = 8'h85 == _GEN_13607 ? 1'h0 : valid_133_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_137 = 8'h86 == _GEN_13607 ? 1'h0 : valid_134_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_138 = 8'h87 == _GEN_13607 ? 1'h0 : valid_135_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_139 = 8'h88 == _GEN_13607 ? 1'h0 : valid_136_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_140 = 8'h89 == _GEN_13607 ? 1'h0 : valid_137_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_141 = 8'h8a == _GEN_13607 ? 1'h0 : valid_138_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_142 = 8'h8b == _GEN_13607 ? 1'h0 : valid_139_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_143 = 8'h8c == _GEN_13607 ? 1'h0 : valid_140_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_144 = 8'h8d == _GEN_13607 ? 1'h0 : valid_141_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_145 = 8'h8e == _GEN_13607 ? 1'h0 : valid_142_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_146 = 8'h8f == _GEN_13607 ? 1'h0 : valid_143_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_147 = 8'h90 == _GEN_13607 ? 1'h0 : valid_144_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_148 = 8'h91 == _GEN_13607 ? 1'h0 : valid_145_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_149 = 8'h92 == _GEN_13607 ? 1'h0 : valid_146_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_150 = 8'h93 == _GEN_13607 ? 1'h0 : valid_147_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_151 = 8'h94 == _GEN_13607 ? 1'h0 : valid_148_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_152 = 8'h95 == _GEN_13607 ? 1'h0 : valid_149_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_153 = 8'h96 == _GEN_13607 ? 1'h0 : valid_150_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_154 = 8'h97 == _GEN_13607 ? 1'h0 : valid_151_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_155 = 8'h98 == _GEN_13607 ? 1'h0 : valid_152_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_156 = 8'h99 == _GEN_13607 ? 1'h0 : valid_153_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_157 = 8'h9a == _GEN_13607 ? 1'h0 : valid_154_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_158 = 8'h9b == _GEN_13607 ? 1'h0 : valid_155_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_159 = 8'h9c == _GEN_13607 ? 1'h0 : valid_156_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_160 = 8'h9d == _GEN_13607 ? 1'h0 : valid_157_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_161 = 8'h9e == _GEN_13607 ? 1'h0 : valid_158_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_162 = 8'h9f == _GEN_13607 ? 1'h0 : valid_159_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_163 = 8'ha0 == _GEN_13607 ? 1'h0 : valid_160_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_164 = 8'ha1 == _GEN_13607 ? 1'h0 : valid_161_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_165 = 8'ha2 == _GEN_13607 ? 1'h0 : valid_162_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_166 = 8'ha3 == _GEN_13607 ? 1'h0 : valid_163_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_167 = 8'ha4 == _GEN_13607 ? 1'h0 : valid_164_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_168 = 8'ha5 == _GEN_13607 ? 1'h0 : valid_165_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_169 = 8'ha6 == _GEN_13607 ? 1'h0 : valid_166_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_170 = 8'ha7 == _GEN_13607 ? 1'h0 : valid_167_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_171 = 8'ha8 == _GEN_13607 ? 1'h0 : valid_168_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_172 = 8'ha9 == _GEN_13607 ? 1'h0 : valid_169_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_173 = 8'haa == _GEN_13607 ? 1'h0 : valid_170_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_174 = 8'hab == _GEN_13607 ? 1'h0 : valid_171_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_175 = 8'hac == _GEN_13607 ? 1'h0 : valid_172_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_176 = 8'had == _GEN_13607 ? 1'h0 : valid_173_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_177 = 8'hae == _GEN_13607 ? 1'h0 : valid_174_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_178 = 8'haf == _GEN_13607 ? 1'h0 : valid_175_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_179 = 8'hb0 == _GEN_13607 ? 1'h0 : valid_176_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_180 = 8'hb1 == _GEN_13607 ? 1'h0 : valid_177_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_181 = 8'hb2 == _GEN_13607 ? 1'h0 : valid_178_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_182 = 8'hb3 == _GEN_13607 ? 1'h0 : valid_179_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_183 = 8'hb4 == _GEN_13607 ? 1'h0 : valid_180_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_184 = 8'hb5 == _GEN_13607 ? 1'h0 : valid_181_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_185 = 8'hb6 == _GEN_13607 ? 1'h0 : valid_182_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_186 = 8'hb7 == _GEN_13607 ? 1'h0 : valid_183_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_187 = 8'hb8 == _GEN_13607 ? 1'h0 : valid_184_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_188 = 8'hb9 == _GEN_13607 ? 1'h0 : valid_185_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_189 = 8'hba == _GEN_13607 ? 1'h0 : valid_186_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_190 = 8'hbb == _GEN_13607 ? 1'h0 : valid_187_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_191 = 8'hbc == _GEN_13607 ? 1'h0 : valid_188_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_192 = 8'hbd == _GEN_13607 ? 1'h0 : valid_189_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_193 = 8'hbe == _GEN_13607 ? 1'h0 : valid_190_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_194 = 8'hbf == _GEN_13607 ? 1'h0 : valid_191_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_195 = 8'hc0 == _GEN_13607 ? 1'h0 : valid_192_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_196 = 8'hc1 == _GEN_13607 ? 1'h0 : valid_193_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_197 = 8'hc2 == _GEN_13607 ? 1'h0 : valid_194_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_198 = 8'hc3 == _GEN_13607 ? 1'h0 : valid_195_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_199 = 8'hc4 == _GEN_13607 ? 1'h0 : valid_196_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_200 = 8'hc5 == _GEN_13607 ? 1'h0 : valid_197_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_201 = 8'hc6 == _GEN_13607 ? 1'h0 : valid_198_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_202 = 8'hc7 == _GEN_13607 ? 1'h0 : valid_199_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_203 = 8'hc8 == _GEN_13607 ? 1'h0 : valid_200_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_204 = 8'hc9 == _GEN_13607 ? 1'h0 : valid_201_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_205 = 8'hca == _GEN_13607 ? 1'h0 : valid_202_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_206 = 8'hcb == _GEN_13607 ? 1'h0 : valid_203_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_207 = 8'hcc == _GEN_13607 ? 1'h0 : valid_204_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_208 = 8'hcd == _GEN_13607 ? 1'h0 : valid_205_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_209 = 8'hce == _GEN_13607 ? 1'h0 : valid_206_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_210 = 8'hcf == _GEN_13607 ? 1'h0 : valid_207_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_211 = 8'hd0 == _GEN_13607 ? 1'h0 : valid_208_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_212 = 8'hd1 == _GEN_13607 ? 1'h0 : valid_209_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_213 = 8'hd2 == _GEN_13607 ? 1'h0 : valid_210_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_214 = 8'hd3 == _GEN_13607 ? 1'h0 : valid_211_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_215 = 8'hd4 == _GEN_13607 ? 1'h0 : valid_212_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_216 = 8'hd5 == _GEN_13607 ? 1'h0 : valid_213_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_217 = 8'hd6 == _GEN_13607 ? 1'h0 : valid_214_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_218 = 8'hd7 == _GEN_13607 ? 1'h0 : valid_215_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_219 = 8'hd8 == _GEN_13607 ? 1'h0 : valid_216_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_220 = 8'hd9 == _GEN_13607 ? 1'h0 : valid_217_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_221 = 8'hda == _GEN_13607 ? 1'h0 : valid_218_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_222 = 8'hdb == _GEN_13607 ? 1'h0 : valid_219_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_223 = 8'hdc == _GEN_13607 ? 1'h0 : valid_220_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_224 = 8'hdd == _GEN_13607 ? 1'h0 : valid_221_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_225 = 8'hde == _GEN_13607 ? 1'h0 : valid_222_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_226 = 8'hdf == _GEN_13607 ? 1'h0 : valid_223_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_227 = 8'he0 == _GEN_13607 ? 1'h0 : valid_224_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_228 = 8'he1 == _GEN_13607 ? 1'h0 : valid_225_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_229 = 8'he2 == _GEN_13607 ? 1'h0 : valid_226_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_230 = 8'he3 == _GEN_13607 ? 1'h0 : valid_227_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_231 = 8'he4 == _GEN_13607 ? 1'h0 : valid_228_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_232 = 8'he5 == _GEN_13607 ? 1'h0 : valid_229_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_233 = 8'he6 == _GEN_13607 ? 1'h0 : valid_230_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_234 = 8'he7 == _GEN_13607 ? 1'h0 : valid_231_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_235 = 8'he8 == _GEN_13607 ? 1'h0 : valid_232_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_236 = 8'he9 == _GEN_13607 ? 1'h0 : valid_233_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_237 = 8'hea == _GEN_13607 ? 1'h0 : valid_234_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_238 = 8'heb == _GEN_13607 ? 1'h0 : valid_235_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_239 = 8'hec == _GEN_13607 ? 1'h0 : valid_236_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_240 = 8'hed == _GEN_13607 ? 1'h0 : valid_237_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_241 = 8'hee == _GEN_13607 ? 1'h0 : valid_238_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_242 = 8'hef == _GEN_13607 ? 1'h0 : valid_239_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_243 = 8'hf0 == _GEN_13607 ? 1'h0 : valid_240_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_244 = 8'hf1 == _GEN_13607 ? 1'h0 : valid_241_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_245 = 8'hf2 == _GEN_13607 ? 1'h0 : valid_242_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_246 = 8'hf3 == _GEN_13607 ? 1'h0 : valid_243_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_247 = 8'hf4 == _GEN_13607 ? 1'h0 : valid_244_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_248 = 8'hf5 == _GEN_13607 ? 1'h0 : valid_245_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_249 = 8'hf6 == _GEN_13607 ? 1'h0 : valid_246_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_250 = 8'hf7 == _GEN_13607 ? 1'h0 : valid_247_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_251 = 8'hf8 == _GEN_13607 ? 1'h0 : valid_248_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_252 = 8'hf9 == _GEN_13607 ? 1'h0 : valid_249_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_253 = 8'hfa == _GEN_13607 ? 1'h0 : valid_250_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_254 = 8'hfb == _GEN_13607 ? 1'h0 : valid_251_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_255 = 8'hfc == _GEN_13607 ? 1'h0 : valid_252_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_256 = 8'hfd == _GEN_13607 ? 1'h0 : valid_253_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_257 = 8'hfe == _GEN_13607 ? 1'h0 : valid_254_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_258 = 8'hff == _GEN_13607 ? 1'h0 : valid_255_0; // @[ICache.scala 52:22 89:{24,24}]
  wire [8:0] _GEN_13735 = {{3'd0}, fence_index}; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_259 = 9'h100 == _GEN_13735 ? 1'h0 : valid_256_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_260 = 9'h101 == _GEN_13735 ? 1'h0 : valid_257_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_261 = 9'h102 == _GEN_13735 ? 1'h0 : valid_258_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_262 = 9'h103 == _GEN_13735 ? 1'h0 : valid_259_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_263 = 9'h104 == _GEN_13735 ? 1'h0 : valid_260_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_264 = 9'h105 == _GEN_13735 ? 1'h0 : valid_261_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_265 = 9'h106 == _GEN_13735 ? 1'h0 : valid_262_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_266 = 9'h107 == _GEN_13735 ? 1'h0 : valid_263_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_267 = 9'h108 == _GEN_13735 ? 1'h0 : valid_264_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_268 = 9'h109 == _GEN_13735 ? 1'h0 : valid_265_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_269 = 9'h10a == _GEN_13735 ? 1'h0 : valid_266_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_270 = 9'h10b == _GEN_13735 ? 1'h0 : valid_267_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_271 = 9'h10c == _GEN_13735 ? 1'h0 : valid_268_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_272 = 9'h10d == _GEN_13735 ? 1'h0 : valid_269_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_273 = 9'h10e == _GEN_13735 ? 1'h0 : valid_270_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_274 = 9'h10f == _GEN_13735 ? 1'h0 : valid_271_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_275 = 9'h110 == _GEN_13735 ? 1'h0 : valid_272_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_276 = 9'h111 == _GEN_13735 ? 1'h0 : valid_273_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_277 = 9'h112 == _GEN_13735 ? 1'h0 : valid_274_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_278 = 9'h113 == _GEN_13735 ? 1'h0 : valid_275_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_279 = 9'h114 == _GEN_13735 ? 1'h0 : valid_276_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_280 = 9'h115 == _GEN_13735 ? 1'h0 : valid_277_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_281 = 9'h116 == _GEN_13735 ? 1'h0 : valid_278_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_282 = 9'h117 == _GEN_13735 ? 1'h0 : valid_279_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_283 = 9'h118 == _GEN_13735 ? 1'h0 : valid_280_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_284 = 9'h119 == _GEN_13735 ? 1'h0 : valid_281_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_285 = 9'h11a == _GEN_13735 ? 1'h0 : valid_282_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_286 = 9'h11b == _GEN_13735 ? 1'h0 : valid_283_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_287 = 9'h11c == _GEN_13735 ? 1'h0 : valid_284_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_288 = 9'h11d == _GEN_13735 ? 1'h0 : valid_285_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_289 = 9'h11e == _GEN_13735 ? 1'h0 : valid_286_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_290 = 9'h11f == _GEN_13735 ? 1'h0 : valid_287_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_291 = 9'h120 == _GEN_13735 ? 1'h0 : valid_288_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_292 = 9'h121 == _GEN_13735 ? 1'h0 : valid_289_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_293 = 9'h122 == _GEN_13735 ? 1'h0 : valid_290_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_294 = 9'h123 == _GEN_13735 ? 1'h0 : valid_291_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_295 = 9'h124 == _GEN_13735 ? 1'h0 : valid_292_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_296 = 9'h125 == _GEN_13735 ? 1'h0 : valid_293_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_297 = 9'h126 == _GEN_13735 ? 1'h0 : valid_294_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_298 = 9'h127 == _GEN_13735 ? 1'h0 : valid_295_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_299 = 9'h128 == _GEN_13735 ? 1'h0 : valid_296_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_300 = 9'h129 == _GEN_13735 ? 1'h0 : valid_297_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_301 = 9'h12a == _GEN_13735 ? 1'h0 : valid_298_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_302 = 9'h12b == _GEN_13735 ? 1'h0 : valid_299_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_303 = 9'h12c == _GEN_13735 ? 1'h0 : valid_300_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_304 = 9'h12d == _GEN_13735 ? 1'h0 : valid_301_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_305 = 9'h12e == _GEN_13735 ? 1'h0 : valid_302_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_306 = 9'h12f == _GEN_13735 ? 1'h0 : valid_303_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_307 = 9'h130 == _GEN_13735 ? 1'h0 : valid_304_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_308 = 9'h131 == _GEN_13735 ? 1'h0 : valid_305_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_309 = 9'h132 == _GEN_13735 ? 1'h0 : valid_306_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_310 = 9'h133 == _GEN_13735 ? 1'h0 : valid_307_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_311 = 9'h134 == _GEN_13735 ? 1'h0 : valid_308_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_312 = 9'h135 == _GEN_13735 ? 1'h0 : valid_309_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_313 = 9'h136 == _GEN_13735 ? 1'h0 : valid_310_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_314 = 9'h137 == _GEN_13735 ? 1'h0 : valid_311_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_315 = 9'h138 == _GEN_13735 ? 1'h0 : valid_312_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_316 = 9'h139 == _GEN_13735 ? 1'h0 : valid_313_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_317 = 9'h13a == _GEN_13735 ? 1'h0 : valid_314_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_318 = 9'h13b == _GEN_13735 ? 1'h0 : valid_315_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_319 = 9'h13c == _GEN_13735 ? 1'h0 : valid_316_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_320 = 9'h13d == _GEN_13735 ? 1'h0 : valid_317_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_321 = 9'h13e == _GEN_13735 ? 1'h0 : valid_318_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_322 = 9'h13f == _GEN_13735 ? 1'h0 : valid_319_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_323 = 9'h140 == _GEN_13735 ? 1'h0 : valid_320_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_324 = 9'h141 == _GEN_13735 ? 1'h0 : valid_321_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_325 = 9'h142 == _GEN_13735 ? 1'h0 : valid_322_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_326 = 9'h143 == _GEN_13735 ? 1'h0 : valid_323_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_327 = 9'h144 == _GEN_13735 ? 1'h0 : valid_324_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_328 = 9'h145 == _GEN_13735 ? 1'h0 : valid_325_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_329 = 9'h146 == _GEN_13735 ? 1'h0 : valid_326_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_330 = 9'h147 == _GEN_13735 ? 1'h0 : valid_327_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_331 = 9'h148 == _GEN_13735 ? 1'h0 : valid_328_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_332 = 9'h149 == _GEN_13735 ? 1'h0 : valid_329_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_333 = 9'h14a == _GEN_13735 ? 1'h0 : valid_330_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_334 = 9'h14b == _GEN_13735 ? 1'h0 : valid_331_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_335 = 9'h14c == _GEN_13735 ? 1'h0 : valid_332_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_336 = 9'h14d == _GEN_13735 ? 1'h0 : valid_333_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_337 = 9'h14e == _GEN_13735 ? 1'h0 : valid_334_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_338 = 9'h14f == _GEN_13735 ? 1'h0 : valid_335_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_339 = 9'h150 == _GEN_13735 ? 1'h0 : valid_336_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_340 = 9'h151 == _GEN_13735 ? 1'h0 : valid_337_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_341 = 9'h152 == _GEN_13735 ? 1'h0 : valid_338_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_342 = 9'h153 == _GEN_13735 ? 1'h0 : valid_339_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_343 = 9'h154 == _GEN_13735 ? 1'h0 : valid_340_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_344 = 9'h155 == _GEN_13735 ? 1'h0 : valid_341_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_345 = 9'h156 == _GEN_13735 ? 1'h0 : valid_342_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_346 = 9'h157 == _GEN_13735 ? 1'h0 : valid_343_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_347 = 9'h158 == _GEN_13735 ? 1'h0 : valid_344_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_348 = 9'h159 == _GEN_13735 ? 1'h0 : valid_345_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_349 = 9'h15a == _GEN_13735 ? 1'h0 : valid_346_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_350 = 9'h15b == _GEN_13735 ? 1'h0 : valid_347_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_351 = 9'h15c == _GEN_13735 ? 1'h0 : valid_348_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_352 = 9'h15d == _GEN_13735 ? 1'h0 : valid_349_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_353 = 9'h15e == _GEN_13735 ? 1'h0 : valid_350_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_354 = 9'h15f == _GEN_13735 ? 1'h0 : valid_351_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_355 = 9'h160 == _GEN_13735 ? 1'h0 : valid_352_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_356 = 9'h161 == _GEN_13735 ? 1'h0 : valid_353_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_357 = 9'h162 == _GEN_13735 ? 1'h0 : valid_354_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_358 = 9'h163 == _GEN_13735 ? 1'h0 : valid_355_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_359 = 9'h164 == _GEN_13735 ? 1'h0 : valid_356_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_360 = 9'h165 == _GEN_13735 ? 1'h0 : valid_357_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_361 = 9'h166 == _GEN_13735 ? 1'h0 : valid_358_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_362 = 9'h167 == _GEN_13735 ? 1'h0 : valid_359_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_363 = 9'h168 == _GEN_13735 ? 1'h0 : valid_360_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_364 = 9'h169 == _GEN_13735 ? 1'h0 : valid_361_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_365 = 9'h16a == _GEN_13735 ? 1'h0 : valid_362_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_366 = 9'h16b == _GEN_13735 ? 1'h0 : valid_363_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_367 = 9'h16c == _GEN_13735 ? 1'h0 : valid_364_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_368 = 9'h16d == _GEN_13735 ? 1'h0 : valid_365_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_369 = 9'h16e == _GEN_13735 ? 1'h0 : valid_366_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_370 = 9'h16f == _GEN_13735 ? 1'h0 : valid_367_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_371 = 9'h170 == _GEN_13735 ? 1'h0 : valid_368_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_372 = 9'h171 == _GEN_13735 ? 1'h0 : valid_369_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_373 = 9'h172 == _GEN_13735 ? 1'h0 : valid_370_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_374 = 9'h173 == _GEN_13735 ? 1'h0 : valid_371_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_375 = 9'h174 == _GEN_13735 ? 1'h0 : valid_372_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_376 = 9'h175 == _GEN_13735 ? 1'h0 : valid_373_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_377 = 9'h176 == _GEN_13735 ? 1'h0 : valid_374_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_378 = 9'h177 == _GEN_13735 ? 1'h0 : valid_375_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_379 = 9'h178 == _GEN_13735 ? 1'h0 : valid_376_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_380 = 9'h179 == _GEN_13735 ? 1'h0 : valid_377_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_381 = 9'h17a == _GEN_13735 ? 1'h0 : valid_378_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_382 = 9'h17b == _GEN_13735 ? 1'h0 : valid_379_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_383 = 9'h17c == _GEN_13735 ? 1'h0 : valid_380_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_384 = 9'h17d == _GEN_13735 ? 1'h0 : valid_381_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_385 = 9'h17e == _GEN_13735 ? 1'h0 : valid_382_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_386 = 9'h17f == _GEN_13735 ? 1'h0 : valid_383_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_387 = 9'h180 == _GEN_13735 ? 1'h0 : valid_384_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_388 = 9'h181 == _GEN_13735 ? 1'h0 : valid_385_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_389 = 9'h182 == _GEN_13735 ? 1'h0 : valid_386_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_390 = 9'h183 == _GEN_13735 ? 1'h0 : valid_387_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_391 = 9'h184 == _GEN_13735 ? 1'h0 : valid_388_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_392 = 9'h185 == _GEN_13735 ? 1'h0 : valid_389_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_393 = 9'h186 == _GEN_13735 ? 1'h0 : valid_390_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_394 = 9'h187 == _GEN_13735 ? 1'h0 : valid_391_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_395 = 9'h188 == _GEN_13735 ? 1'h0 : valid_392_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_396 = 9'h189 == _GEN_13735 ? 1'h0 : valid_393_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_397 = 9'h18a == _GEN_13735 ? 1'h0 : valid_394_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_398 = 9'h18b == _GEN_13735 ? 1'h0 : valid_395_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_399 = 9'h18c == _GEN_13735 ? 1'h0 : valid_396_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_400 = 9'h18d == _GEN_13735 ? 1'h0 : valid_397_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_401 = 9'h18e == _GEN_13735 ? 1'h0 : valid_398_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_402 = 9'h18f == _GEN_13735 ? 1'h0 : valid_399_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_403 = 9'h190 == _GEN_13735 ? 1'h0 : valid_400_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_404 = 9'h191 == _GEN_13735 ? 1'h0 : valid_401_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_405 = 9'h192 == _GEN_13735 ? 1'h0 : valid_402_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_406 = 9'h193 == _GEN_13735 ? 1'h0 : valid_403_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_407 = 9'h194 == _GEN_13735 ? 1'h0 : valid_404_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_408 = 9'h195 == _GEN_13735 ? 1'h0 : valid_405_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_409 = 9'h196 == _GEN_13735 ? 1'h0 : valid_406_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_410 = 9'h197 == _GEN_13735 ? 1'h0 : valid_407_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_411 = 9'h198 == _GEN_13735 ? 1'h0 : valid_408_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_412 = 9'h199 == _GEN_13735 ? 1'h0 : valid_409_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_413 = 9'h19a == _GEN_13735 ? 1'h0 : valid_410_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_414 = 9'h19b == _GEN_13735 ? 1'h0 : valid_411_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_415 = 9'h19c == _GEN_13735 ? 1'h0 : valid_412_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_416 = 9'h19d == _GEN_13735 ? 1'h0 : valid_413_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_417 = 9'h19e == _GEN_13735 ? 1'h0 : valid_414_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_418 = 9'h19f == _GEN_13735 ? 1'h0 : valid_415_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_419 = 9'h1a0 == _GEN_13735 ? 1'h0 : valid_416_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_420 = 9'h1a1 == _GEN_13735 ? 1'h0 : valid_417_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_421 = 9'h1a2 == _GEN_13735 ? 1'h0 : valid_418_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_422 = 9'h1a3 == _GEN_13735 ? 1'h0 : valid_419_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_423 = 9'h1a4 == _GEN_13735 ? 1'h0 : valid_420_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_424 = 9'h1a5 == _GEN_13735 ? 1'h0 : valid_421_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_425 = 9'h1a6 == _GEN_13735 ? 1'h0 : valid_422_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_426 = 9'h1a7 == _GEN_13735 ? 1'h0 : valid_423_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_427 = 9'h1a8 == _GEN_13735 ? 1'h0 : valid_424_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_428 = 9'h1a9 == _GEN_13735 ? 1'h0 : valid_425_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_429 = 9'h1aa == _GEN_13735 ? 1'h0 : valid_426_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_430 = 9'h1ab == _GEN_13735 ? 1'h0 : valid_427_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_431 = 9'h1ac == _GEN_13735 ? 1'h0 : valid_428_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_432 = 9'h1ad == _GEN_13735 ? 1'h0 : valid_429_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_433 = 9'h1ae == _GEN_13735 ? 1'h0 : valid_430_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_434 = 9'h1af == _GEN_13735 ? 1'h0 : valid_431_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_435 = 9'h1b0 == _GEN_13735 ? 1'h0 : valid_432_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_436 = 9'h1b1 == _GEN_13735 ? 1'h0 : valid_433_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_437 = 9'h1b2 == _GEN_13735 ? 1'h0 : valid_434_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_438 = 9'h1b3 == _GEN_13735 ? 1'h0 : valid_435_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_439 = 9'h1b4 == _GEN_13735 ? 1'h0 : valid_436_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_440 = 9'h1b5 == _GEN_13735 ? 1'h0 : valid_437_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_441 = 9'h1b6 == _GEN_13735 ? 1'h0 : valid_438_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_442 = 9'h1b7 == _GEN_13735 ? 1'h0 : valid_439_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_443 = 9'h1b8 == _GEN_13735 ? 1'h0 : valid_440_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_444 = 9'h1b9 == _GEN_13735 ? 1'h0 : valid_441_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_445 = 9'h1ba == _GEN_13735 ? 1'h0 : valid_442_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_446 = 9'h1bb == _GEN_13735 ? 1'h0 : valid_443_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_447 = 9'h1bc == _GEN_13735 ? 1'h0 : valid_444_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_448 = 9'h1bd == _GEN_13735 ? 1'h0 : valid_445_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_449 = 9'h1be == _GEN_13735 ? 1'h0 : valid_446_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_450 = 9'h1bf == _GEN_13735 ? 1'h0 : valid_447_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_451 = 9'h1c0 == _GEN_13735 ? 1'h0 : valid_448_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_452 = 9'h1c1 == _GEN_13735 ? 1'h0 : valid_449_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_453 = 9'h1c2 == _GEN_13735 ? 1'h0 : valid_450_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_454 = 9'h1c3 == _GEN_13735 ? 1'h0 : valid_451_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_455 = 9'h1c4 == _GEN_13735 ? 1'h0 : valid_452_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_456 = 9'h1c5 == _GEN_13735 ? 1'h0 : valid_453_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_457 = 9'h1c6 == _GEN_13735 ? 1'h0 : valid_454_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_458 = 9'h1c7 == _GEN_13735 ? 1'h0 : valid_455_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_459 = 9'h1c8 == _GEN_13735 ? 1'h0 : valid_456_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_460 = 9'h1c9 == _GEN_13735 ? 1'h0 : valid_457_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_461 = 9'h1ca == _GEN_13735 ? 1'h0 : valid_458_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_462 = 9'h1cb == _GEN_13735 ? 1'h0 : valid_459_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_463 = 9'h1cc == _GEN_13735 ? 1'h0 : valid_460_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_464 = 9'h1cd == _GEN_13735 ? 1'h0 : valid_461_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_465 = 9'h1ce == _GEN_13735 ? 1'h0 : valid_462_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_466 = 9'h1cf == _GEN_13735 ? 1'h0 : valid_463_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_467 = 9'h1d0 == _GEN_13735 ? 1'h0 : valid_464_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_468 = 9'h1d1 == _GEN_13735 ? 1'h0 : valid_465_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_469 = 9'h1d2 == _GEN_13735 ? 1'h0 : valid_466_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_470 = 9'h1d3 == _GEN_13735 ? 1'h0 : valid_467_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_471 = 9'h1d4 == _GEN_13735 ? 1'h0 : valid_468_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_472 = 9'h1d5 == _GEN_13735 ? 1'h0 : valid_469_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_473 = 9'h1d6 == _GEN_13735 ? 1'h0 : valid_470_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_474 = 9'h1d7 == _GEN_13735 ? 1'h0 : valid_471_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_475 = 9'h1d8 == _GEN_13735 ? 1'h0 : valid_472_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_476 = 9'h1d9 == _GEN_13735 ? 1'h0 : valid_473_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_477 = 9'h1da == _GEN_13735 ? 1'h0 : valid_474_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_478 = 9'h1db == _GEN_13735 ? 1'h0 : valid_475_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_479 = 9'h1dc == _GEN_13735 ? 1'h0 : valid_476_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_480 = 9'h1dd == _GEN_13735 ? 1'h0 : valid_477_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_481 = 9'h1de == _GEN_13735 ? 1'h0 : valid_478_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_482 = 9'h1df == _GEN_13735 ? 1'h0 : valid_479_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_483 = 9'h1e0 == _GEN_13735 ? 1'h0 : valid_480_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_484 = 9'h1e1 == _GEN_13735 ? 1'h0 : valid_481_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_485 = 9'h1e2 == _GEN_13735 ? 1'h0 : valid_482_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_486 = 9'h1e3 == _GEN_13735 ? 1'h0 : valid_483_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_487 = 9'h1e4 == _GEN_13735 ? 1'h0 : valid_484_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_488 = 9'h1e5 == _GEN_13735 ? 1'h0 : valid_485_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_489 = 9'h1e6 == _GEN_13735 ? 1'h0 : valid_486_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_490 = 9'h1e7 == _GEN_13735 ? 1'h0 : valid_487_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_491 = 9'h1e8 == _GEN_13735 ? 1'h0 : valid_488_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_492 = 9'h1e9 == _GEN_13735 ? 1'h0 : valid_489_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_493 = 9'h1ea == _GEN_13735 ? 1'h0 : valid_490_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_494 = 9'h1eb == _GEN_13735 ? 1'h0 : valid_491_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_495 = 9'h1ec == _GEN_13735 ? 1'h0 : valid_492_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_496 = 9'h1ed == _GEN_13735 ? 1'h0 : valid_493_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_497 = 9'h1ee == _GEN_13735 ? 1'h0 : valid_494_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_498 = 9'h1ef == _GEN_13735 ? 1'h0 : valid_495_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_499 = 9'h1f0 == _GEN_13735 ? 1'h0 : valid_496_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_500 = 9'h1f1 == _GEN_13735 ? 1'h0 : valid_497_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_501 = 9'h1f2 == _GEN_13735 ? 1'h0 : valid_498_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_502 = 9'h1f3 == _GEN_13735 ? 1'h0 : valid_499_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_503 = 9'h1f4 == _GEN_13735 ? 1'h0 : valid_500_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_504 = 9'h1f5 == _GEN_13735 ? 1'h0 : valid_501_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_505 = 9'h1f6 == _GEN_13735 ? 1'h0 : valid_502_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_506 = 9'h1f7 == _GEN_13735 ? 1'h0 : valid_503_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_507 = 9'h1f8 == _GEN_13735 ? 1'h0 : valid_504_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_508 = 9'h1f9 == _GEN_13735 ? 1'h0 : valid_505_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_509 = 9'h1fa == _GEN_13735 ? 1'h0 : valid_506_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_510 = 9'h1fb == _GEN_13735 ? 1'h0 : valid_507_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_511 = 9'h1fc == _GEN_13735 ? 1'h0 : valid_508_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_512 = 9'h1fd == _GEN_13735 ? 1'h0 : valid_509_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_513 = 9'h1fe == _GEN_13735 ? 1'h0 : valid_510_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_514 = 9'h1ff == _GEN_13735 ? 1'h0 : valid_511_0; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_515 = 6'h0 == fence_index ? 1'h0 : valid_0_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_516 = 6'h1 == fence_index ? 1'h0 : valid_1_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_517 = 6'h2 == fence_index ? 1'h0 : valid_2_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_518 = 6'h3 == fence_index ? 1'h0 : valid_3_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_519 = 6'h4 == fence_index ? 1'h0 : valid_4_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_520 = 6'h5 == fence_index ? 1'h0 : valid_5_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_521 = 6'h6 == fence_index ? 1'h0 : valid_6_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_522 = 6'h7 == fence_index ? 1'h0 : valid_7_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_523 = 6'h8 == fence_index ? 1'h0 : valid_8_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_524 = 6'h9 == fence_index ? 1'h0 : valid_9_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_525 = 6'ha == fence_index ? 1'h0 : valid_10_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_526 = 6'hb == fence_index ? 1'h0 : valid_11_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_527 = 6'hc == fence_index ? 1'h0 : valid_12_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_528 = 6'hd == fence_index ? 1'h0 : valid_13_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_529 = 6'he == fence_index ? 1'h0 : valid_14_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_530 = 6'hf == fence_index ? 1'h0 : valid_15_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_531 = 6'h10 == fence_index ? 1'h0 : valid_16_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_532 = 6'h11 == fence_index ? 1'h0 : valid_17_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_533 = 6'h12 == fence_index ? 1'h0 : valid_18_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_534 = 6'h13 == fence_index ? 1'h0 : valid_19_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_535 = 6'h14 == fence_index ? 1'h0 : valid_20_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_536 = 6'h15 == fence_index ? 1'h0 : valid_21_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_537 = 6'h16 == fence_index ? 1'h0 : valid_22_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_538 = 6'h17 == fence_index ? 1'h0 : valid_23_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_539 = 6'h18 == fence_index ? 1'h0 : valid_24_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_540 = 6'h19 == fence_index ? 1'h0 : valid_25_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_541 = 6'h1a == fence_index ? 1'h0 : valid_26_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_542 = 6'h1b == fence_index ? 1'h0 : valid_27_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_543 = 6'h1c == fence_index ? 1'h0 : valid_28_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_544 = 6'h1d == fence_index ? 1'h0 : valid_29_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_545 = 6'h1e == fence_index ? 1'h0 : valid_30_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_546 = 6'h1f == fence_index ? 1'h0 : valid_31_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_547 = 6'h20 == fence_index ? 1'h0 : valid_32_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_548 = 6'h21 == fence_index ? 1'h0 : valid_33_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_549 = 6'h22 == fence_index ? 1'h0 : valid_34_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_550 = 6'h23 == fence_index ? 1'h0 : valid_35_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_551 = 6'h24 == fence_index ? 1'h0 : valid_36_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_552 = 6'h25 == fence_index ? 1'h0 : valid_37_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_553 = 6'h26 == fence_index ? 1'h0 : valid_38_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_554 = 6'h27 == fence_index ? 1'h0 : valid_39_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_555 = 6'h28 == fence_index ? 1'h0 : valid_40_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_556 = 6'h29 == fence_index ? 1'h0 : valid_41_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_557 = 6'h2a == fence_index ? 1'h0 : valid_42_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_558 = 6'h2b == fence_index ? 1'h0 : valid_43_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_559 = 6'h2c == fence_index ? 1'h0 : valid_44_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_560 = 6'h2d == fence_index ? 1'h0 : valid_45_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_561 = 6'h2e == fence_index ? 1'h0 : valid_46_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_562 = 6'h2f == fence_index ? 1'h0 : valid_47_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_563 = 6'h30 == fence_index ? 1'h0 : valid_48_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_564 = 6'h31 == fence_index ? 1'h0 : valid_49_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_565 = 6'h32 == fence_index ? 1'h0 : valid_50_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_566 = 6'h33 == fence_index ? 1'h0 : valid_51_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_567 = 6'h34 == fence_index ? 1'h0 : valid_52_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_568 = 6'h35 == fence_index ? 1'h0 : valid_53_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_569 = 6'h36 == fence_index ? 1'h0 : valid_54_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_570 = 6'h37 == fence_index ? 1'h0 : valid_55_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_571 = 6'h38 == fence_index ? 1'h0 : valid_56_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_572 = 6'h39 == fence_index ? 1'h0 : valid_57_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_573 = 6'h3a == fence_index ? 1'h0 : valid_58_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_574 = 6'h3b == fence_index ? 1'h0 : valid_59_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_575 = 6'h3c == fence_index ? 1'h0 : valid_60_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_576 = 6'h3d == fence_index ? 1'h0 : valid_61_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_577 = 6'h3e == fence_index ? 1'h0 : valid_62_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_578 = 6'h3f == fence_index ? 1'h0 : valid_63_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_579 = 7'h40 == _GEN_13543 ? 1'h0 : valid_64_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_580 = 7'h41 == _GEN_13543 ? 1'h0 : valid_65_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_581 = 7'h42 == _GEN_13543 ? 1'h0 : valid_66_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_582 = 7'h43 == _GEN_13543 ? 1'h0 : valid_67_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_583 = 7'h44 == _GEN_13543 ? 1'h0 : valid_68_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_584 = 7'h45 == _GEN_13543 ? 1'h0 : valid_69_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_585 = 7'h46 == _GEN_13543 ? 1'h0 : valid_70_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_586 = 7'h47 == _GEN_13543 ? 1'h0 : valid_71_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_587 = 7'h48 == _GEN_13543 ? 1'h0 : valid_72_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_588 = 7'h49 == _GEN_13543 ? 1'h0 : valid_73_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_589 = 7'h4a == _GEN_13543 ? 1'h0 : valid_74_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_590 = 7'h4b == _GEN_13543 ? 1'h0 : valid_75_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_591 = 7'h4c == _GEN_13543 ? 1'h0 : valid_76_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_592 = 7'h4d == _GEN_13543 ? 1'h0 : valid_77_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_593 = 7'h4e == _GEN_13543 ? 1'h0 : valid_78_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_594 = 7'h4f == _GEN_13543 ? 1'h0 : valid_79_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_595 = 7'h50 == _GEN_13543 ? 1'h0 : valid_80_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_596 = 7'h51 == _GEN_13543 ? 1'h0 : valid_81_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_597 = 7'h52 == _GEN_13543 ? 1'h0 : valid_82_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_598 = 7'h53 == _GEN_13543 ? 1'h0 : valid_83_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_599 = 7'h54 == _GEN_13543 ? 1'h0 : valid_84_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_600 = 7'h55 == _GEN_13543 ? 1'h0 : valid_85_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_601 = 7'h56 == _GEN_13543 ? 1'h0 : valid_86_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_602 = 7'h57 == _GEN_13543 ? 1'h0 : valid_87_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_603 = 7'h58 == _GEN_13543 ? 1'h0 : valid_88_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_604 = 7'h59 == _GEN_13543 ? 1'h0 : valid_89_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_605 = 7'h5a == _GEN_13543 ? 1'h0 : valid_90_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_606 = 7'h5b == _GEN_13543 ? 1'h0 : valid_91_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_607 = 7'h5c == _GEN_13543 ? 1'h0 : valid_92_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_608 = 7'h5d == _GEN_13543 ? 1'h0 : valid_93_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_609 = 7'h5e == _GEN_13543 ? 1'h0 : valid_94_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_610 = 7'h5f == _GEN_13543 ? 1'h0 : valid_95_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_611 = 7'h60 == _GEN_13543 ? 1'h0 : valid_96_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_612 = 7'h61 == _GEN_13543 ? 1'h0 : valid_97_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_613 = 7'h62 == _GEN_13543 ? 1'h0 : valid_98_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_614 = 7'h63 == _GEN_13543 ? 1'h0 : valid_99_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_615 = 7'h64 == _GEN_13543 ? 1'h0 : valid_100_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_616 = 7'h65 == _GEN_13543 ? 1'h0 : valid_101_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_617 = 7'h66 == _GEN_13543 ? 1'h0 : valid_102_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_618 = 7'h67 == _GEN_13543 ? 1'h0 : valid_103_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_619 = 7'h68 == _GEN_13543 ? 1'h0 : valid_104_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_620 = 7'h69 == _GEN_13543 ? 1'h0 : valid_105_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_621 = 7'h6a == _GEN_13543 ? 1'h0 : valid_106_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_622 = 7'h6b == _GEN_13543 ? 1'h0 : valid_107_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_623 = 7'h6c == _GEN_13543 ? 1'h0 : valid_108_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_624 = 7'h6d == _GEN_13543 ? 1'h0 : valid_109_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_625 = 7'h6e == _GEN_13543 ? 1'h0 : valid_110_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_626 = 7'h6f == _GEN_13543 ? 1'h0 : valid_111_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_627 = 7'h70 == _GEN_13543 ? 1'h0 : valid_112_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_628 = 7'h71 == _GEN_13543 ? 1'h0 : valid_113_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_629 = 7'h72 == _GEN_13543 ? 1'h0 : valid_114_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_630 = 7'h73 == _GEN_13543 ? 1'h0 : valid_115_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_631 = 7'h74 == _GEN_13543 ? 1'h0 : valid_116_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_632 = 7'h75 == _GEN_13543 ? 1'h0 : valid_117_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_633 = 7'h76 == _GEN_13543 ? 1'h0 : valid_118_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_634 = 7'h77 == _GEN_13543 ? 1'h0 : valid_119_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_635 = 7'h78 == _GEN_13543 ? 1'h0 : valid_120_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_636 = 7'h79 == _GEN_13543 ? 1'h0 : valid_121_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_637 = 7'h7a == _GEN_13543 ? 1'h0 : valid_122_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_638 = 7'h7b == _GEN_13543 ? 1'h0 : valid_123_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_639 = 7'h7c == _GEN_13543 ? 1'h0 : valid_124_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_640 = 7'h7d == _GEN_13543 ? 1'h0 : valid_125_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_641 = 7'h7e == _GEN_13543 ? 1'h0 : valid_126_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_642 = 7'h7f == _GEN_13543 ? 1'h0 : valid_127_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_643 = 8'h80 == _GEN_13607 ? 1'h0 : valid_128_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_644 = 8'h81 == _GEN_13607 ? 1'h0 : valid_129_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_645 = 8'h82 == _GEN_13607 ? 1'h0 : valid_130_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_646 = 8'h83 == _GEN_13607 ? 1'h0 : valid_131_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_647 = 8'h84 == _GEN_13607 ? 1'h0 : valid_132_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_648 = 8'h85 == _GEN_13607 ? 1'h0 : valid_133_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_649 = 8'h86 == _GEN_13607 ? 1'h0 : valid_134_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_650 = 8'h87 == _GEN_13607 ? 1'h0 : valid_135_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_651 = 8'h88 == _GEN_13607 ? 1'h0 : valid_136_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_652 = 8'h89 == _GEN_13607 ? 1'h0 : valid_137_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_653 = 8'h8a == _GEN_13607 ? 1'h0 : valid_138_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_654 = 8'h8b == _GEN_13607 ? 1'h0 : valid_139_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_655 = 8'h8c == _GEN_13607 ? 1'h0 : valid_140_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_656 = 8'h8d == _GEN_13607 ? 1'h0 : valid_141_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_657 = 8'h8e == _GEN_13607 ? 1'h0 : valid_142_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_658 = 8'h8f == _GEN_13607 ? 1'h0 : valid_143_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_659 = 8'h90 == _GEN_13607 ? 1'h0 : valid_144_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_660 = 8'h91 == _GEN_13607 ? 1'h0 : valid_145_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_661 = 8'h92 == _GEN_13607 ? 1'h0 : valid_146_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_662 = 8'h93 == _GEN_13607 ? 1'h0 : valid_147_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_663 = 8'h94 == _GEN_13607 ? 1'h0 : valid_148_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_664 = 8'h95 == _GEN_13607 ? 1'h0 : valid_149_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_665 = 8'h96 == _GEN_13607 ? 1'h0 : valid_150_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_666 = 8'h97 == _GEN_13607 ? 1'h0 : valid_151_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_667 = 8'h98 == _GEN_13607 ? 1'h0 : valid_152_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_668 = 8'h99 == _GEN_13607 ? 1'h0 : valid_153_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_669 = 8'h9a == _GEN_13607 ? 1'h0 : valid_154_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_670 = 8'h9b == _GEN_13607 ? 1'h0 : valid_155_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_671 = 8'h9c == _GEN_13607 ? 1'h0 : valid_156_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_672 = 8'h9d == _GEN_13607 ? 1'h0 : valid_157_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_673 = 8'h9e == _GEN_13607 ? 1'h0 : valid_158_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_674 = 8'h9f == _GEN_13607 ? 1'h0 : valid_159_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_675 = 8'ha0 == _GEN_13607 ? 1'h0 : valid_160_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_676 = 8'ha1 == _GEN_13607 ? 1'h0 : valid_161_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_677 = 8'ha2 == _GEN_13607 ? 1'h0 : valid_162_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_678 = 8'ha3 == _GEN_13607 ? 1'h0 : valid_163_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_679 = 8'ha4 == _GEN_13607 ? 1'h0 : valid_164_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_680 = 8'ha5 == _GEN_13607 ? 1'h0 : valid_165_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_681 = 8'ha6 == _GEN_13607 ? 1'h0 : valid_166_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_682 = 8'ha7 == _GEN_13607 ? 1'h0 : valid_167_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_683 = 8'ha8 == _GEN_13607 ? 1'h0 : valid_168_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_684 = 8'ha9 == _GEN_13607 ? 1'h0 : valid_169_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_685 = 8'haa == _GEN_13607 ? 1'h0 : valid_170_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_686 = 8'hab == _GEN_13607 ? 1'h0 : valid_171_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_687 = 8'hac == _GEN_13607 ? 1'h0 : valid_172_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_688 = 8'had == _GEN_13607 ? 1'h0 : valid_173_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_689 = 8'hae == _GEN_13607 ? 1'h0 : valid_174_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_690 = 8'haf == _GEN_13607 ? 1'h0 : valid_175_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_691 = 8'hb0 == _GEN_13607 ? 1'h0 : valid_176_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_692 = 8'hb1 == _GEN_13607 ? 1'h0 : valid_177_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_693 = 8'hb2 == _GEN_13607 ? 1'h0 : valid_178_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_694 = 8'hb3 == _GEN_13607 ? 1'h0 : valid_179_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_695 = 8'hb4 == _GEN_13607 ? 1'h0 : valid_180_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_696 = 8'hb5 == _GEN_13607 ? 1'h0 : valid_181_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_697 = 8'hb6 == _GEN_13607 ? 1'h0 : valid_182_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_698 = 8'hb7 == _GEN_13607 ? 1'h0 : valid_183_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_699 = 8'hb8 == _GEN_13607 ? 1'h0 : valid_184_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_700 = 8'hb9 == _GEN_13607 ? 1'h0 : valid_185_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_701 = 8'hba == _GEN_13607 ? 1'h0 : valid_186_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_702 = 8'hbb == _GEN_13607 ? 1'h0 : valid_187_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_703 = 8'hbc == _GEN_13607 ? 1'h0 : valid_188_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_704 = 8'hbd == _GEN_13607 ? 1'h0 : valid_189_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_705 = 8'hbe == _GEN_13607 ? 1'h0 : valid_190_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_706 = 8'hbf == _GEN_13607 ? 1'h0 : valid_191_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_707 = 8'hc0 == _GEN_13607 ? 1'h0 : valid_192_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_708 = 8'hc1 == _GEN_13607 ? 1'h0 : valid_193_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_709 = 8'hc2 == _GEN_13607 ? 1'h0 : valid_194_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_710 = 8'hc3 == _GEN_13607 ? 1'h0 : valid_195_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_711 = 8'hc4 == _GEN_13607 ? 1'h0 : valid_196_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_712 = 8'hc5 == _GEN_13607 ? 1'h0 : valid_197_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_713 = 8'hc6 == _GEN_13607 ? 1'h0 : valid_198_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_714 = 8'hc7 == _GEN_13607 ? 1'h0 : valid_199_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_715 = 8'hc8 == _GEN_13607 ? 1'h0 : valid_200_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_716 = 8'hc9 == _GEN_13607 ? 1'h0 : valid_201_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_717 = 8'hca == _GEN_13607 ? 1'h0 : valid_202_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_718 = 8'hcb == _GEN_13607 ? 1'h0 : valid_203_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_719 = 8'hcc == _GEN_13607 ? 1'h0 : valid_204_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_720 = 8'hcd == _GEN_13607 ? 1'h0 : valid_205_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_721 = 8'hce == _GEN_13607 ? 1'h0 : valid_206_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_722 = 8'hcf == _GEN_13607 ? 1'h0 : valid_207_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_723 = 8'hd0 == _GEN_13607 ? 1'h0 : valid_208_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_724 = 8'hd1 == _GEN_13607 ? 1'h0 : valid_209_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_725 = 8'hd2 == _GEN_13607 ? 1'h0 : valid_210_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_726 = 8'hd3 == _GEN_13607 ? 1'h0 : valid_211_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_727 = 8'hd4 == _GEN_13607 ? 1'h0 : valid_212_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_728 = 8'hd5 == _GEN_13607 ? 1'h0 : valid_213_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_729 = 8'hd6 == _GEN_13607 ? 1'h0 : valid_214_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_730 = 8'hd7 == _GEN_13607 ? 1'h0 : valid_215_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_731 = 8'hd8 == _GEN_13607 ? 1'h0 : valid_216_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_732 = 8'hd9 == _GEN_13607 ? 1'h0 : valid_217_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_733 = 8'hda == _GEN_13607 ? 1'h0 : valid_218_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_734 = 8'hdb == _GEN_13607 ? 1'h0 : valid_219_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_735 = 8'hdc == _GEN_13607 ? 1'h0 : valid_220_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_736 = 8'hdd == _GEN_13607 ? 1'h0 : valid_221_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_737 = 8'hde == _GEN_13607 ? 1'h0 : valid_222_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_738 = 8'hdf == _GEN_13607 ? 1'h0 : valid_223_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_739 = 8'he0 == _GEN_13607 ? 1'h0 : valid_224_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_740 = 8'he1 == _GEN_13607 ? 1'h0 : valid_225_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_741 = 8'he2 == _GEN_13607 ? 1'h0 : valid_226_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_742 = 8'he3 == _GEN_13607 ? 1'h0 : valid_227_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_743 = 8'he4 == _GEN_13607 ? 1'h0 : valid_228_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_744 = 8'he5 == _GEN_13607 ? 1'h0 : valid_229_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_745 = 8'he6 == _GEN_13607 ? 1'h0 : valid_230_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_746 = 8'he7 == _GEN_13607 ? 1'h0 : valid_231_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_747 = 8'he8 == _GEN_13607 ? 1'h0 : valid_232_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_748 = 8'he9 == _GEN_13607 ? 1'h0 : valid_233_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_749 = 8'hea == _GEN_13607 ? 1'h0 : valid_234_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_750 = 8'heb == _GEN_13607 ? 1'h0 : valid_235_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_751 = 8'hec == _GEN_13607 ? 1'h0 : valid_236_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_752 = 8'hed == _GEN_13607 ? 1'h0 : valid_237_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_753 = 8'hee == _GEN_13607 ? 1'h0 : valid_238_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_754 = 8'hef == _GEN_13607 ? 1'h0 : valid_239_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_755 = 8'hf0 == _GEN_13607 ? 1'h0 : valid_240_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_756 = 8'hf1 == _GEN_13607 ? 1'h0 : valid_241_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_757 = 8'hf2 == _GEN_13607 ? 1'h0 : valid_242_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_758 = 8'hf3 == _GEN_13607 ? 1'h0 : valid_243_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_759 = 8'hf4 == _GEN_13607 ? 1'h0 : valid_244_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_760 = 8'hf5 == _GEN_13607 ? 1'h0 : valid_245_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_761 = 8'hf6 == _GEN_13607 ? 1'h0 : valid_246_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_762 = 8'hf7 == _GEN_13607 ? 1'h0 : valid_247_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_763 = 8'hf8 == _GEN_13607 ? 1'h0 : valid_248_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_764 = 8'hf9 == _GEN_13607 ? 1'h0 : valid_249_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_765 = 8'hfa == _GEN_13607 ? 1'h0 : valid_250_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_766 = 8'hfb == _GEN_13607 ? 1'h0 : valid_251_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_767 = 8'hfc == _GEN_13607 ? 1'h0 : valid_252_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_768 = 8'hfd == _GEN_13607 ? 1'h0 : valid_253_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_769 = 8'hfe == _GEN_13607 ? 1'h0 : valid_254_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_770 = 8'hff == _GEN_13607 ? 1'h0 : valid_255_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_771 = 9'h100 == _GEN_13735 ? 1'h0 : valid_256_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_772 = 9'h101 == _GEN_13735 ? 1'h0 : valid_257_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_773 = 9'h102 == _GEN_13735 ? 1'h0 : valid_258_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_774 = 9'h103 == _GEN_13735 ? 1'h0 : valid_259_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_775 = 9'h104 == _GEN_13735 ? 1'h0 : valid_260_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_776 = 9'h105 == _GEN_13735 ? 1'h0 : valid_261_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_777 = 9'h106 == _GEN_13735 ? 1'h0 : valid_262_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_778 = 9'h107 == _GEN_13735 ? 1'h0 : valid_263_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_779 = 9'h108 == _GEN_13735 ? 1'h0 : valid_264_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_780 = 9'h109 == _GEN_13735 ? 1'h0 : valid_265_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_781 = 9'h10a == _GEN_13735 ? 1'h0 : valid_266_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_782 = 9'h10b == _GEN_13735 ? 1'h0 : valid_267_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_783 = 9'h10c == _GEN_13735 ? 1'h0 : valid_268_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_784 = 9'h10d == _GEN_13735 ? 1'h0 : valid_269_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_785 = 9'h10e == _GEN_13735 ? 1'h0 : valid_270_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_786 = 9'h10f == _GEN_13735 ? 1'h0 : valid_271_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_787 = 9'h110 == _GEN_13735 ? 1'h0 : valid_272_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_788 = 9'h111 == _GEN_13735 ? 1'h0 : valid_273_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_789 = 9'h112 == _GEN_13735 ? 1'h0 : valid_274_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_790 = 9'h113 == _GEN_13735 ? 1'h0 : valid_275_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_791 = 9'h114 == _GEN_13735 ? 1'h0 : valid_276_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_792 = 9'h115 == _GEN_13735 ? 1'h0 : valid_277_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_793 = 9'h116 == _GEN_13735 ? 1'h0 : valid_278_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_794 = 9'h117 == _GEN_13735 ? 1'h0 : valid_279_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_795 = 9'h118 == _GEN_13735 ? 1'h0 : valid_280_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_796 = 9'h119 == _GEN_13735 ? 1'h0 : valid_281_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_797 = 9'h11a == _GEN_13735 ? 1'h0 : valid_282_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_798 = 9'h11b == _GEN_13735 ? 1'h0 : valid_283_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_799 = 9'h11c == _GEN_13735 ? 1'h0 : valid_284_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_800 = 9'h11d == _GEN_13735 ? 1'h0 : valid_285_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_801 = 9'h11e == _GEN_13735 ? 1'h0 : valid_286_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_802 = 9'h11f == _GEN_13735 ? 1'h0 : valid_287_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_803 = 9'h120 == _GEN_13735 ? 1'h0 : valid_288_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_804 = 9'h121 == _GEN_13735 ? 1'h0 : valid_289_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_805 = 9'h122 == _GEN_13735 ? 1'h0 : valid_290_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_806 = 9'h123 == _GEN_13735 ? 1'h0 : valid_291_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_807 = 9'h124 == _GEN_13735 ? 1'h0 : valid_292_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_808 = 9'h125 == _GEN_13735 ? 1'h0 : valid_293_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_809 = 9'h126 == _GEN_13735 ? 1'h0 : valid_294_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_810 = 9'h127 == _GEN_13735 ? 1'h0 : valid_295_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_811 = 9'h128 == _GEN_13735 ? 1'h0 : valid_296_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_812 = 9'h129 == _GEN_13735 ? 1'h0 : valid_297_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_813 = 9'h12a == _GEN_13735 ? 1'h0 : valid_298_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_814 = 9'h12b == _GEN_13735 ? 1'h0 : valid_299_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_815 = 9'h12c == _GEN_13735 ? 1'h0 : valid_300_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_816 = 9'h12d == _GEN_13735 ? 1'h0 : valid_301_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_817 = 9'h12e == _GEN_13735 ? 1'h0 : valid_302_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_818 = 9'h12f == _GEN_13735 ? 1'h0 : valid_303_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_819 = 9'h130 == _GEN_13735 ? 1'h0 : valid_304_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_820 = 9'h131 == _GEN_13735 ? 1'h0 : valid_305_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_821 = 9'h132 == _GEN_13735 ? 1'h0 : valid_306_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_822 = 9'h133 == _GEN_13735 ? 1'h0 : valid_307_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_823 = 9'h134 == _GEN_13735 ? 1'h0 : valid_308_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_824 = 9'h135 == _GEN_13735 ? 1'h0 : valid_309_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_825 = 9'h136 == _GEN_13735 ? 1'h0 : valid_310_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_826 = 9'h137 == _GEN_13735 ? 1'h0 : valid_311_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_827 = 9'h138 == _GEN_13735 ? 1'h0 : valid_312_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_828 = 9'h139 == _GEN_13735 ? 1'h0 : valid_313_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_829 = 9'h13a == _GEN_13735 ? 1'h0 : valid_314_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_830 = 9'h13b == _GEN_13735 ? 1'h0 : valid_315_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_831 = 9'h13c == _GEN_13735 ? 1'h0 : valid_316_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_832 = 9'h13d == _GEN_13735 ? 1'h0 : valid_317_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_833 = 9'h13e == _GEN_13735 ? 1'h0 : valid_318_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_834 = 9'h13f == _GEN_13735 ? 1'h0 : valid_319_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_835 = 9'h140 == _GEN_13735 ? 1'h0 : valid_320_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_836 = 9'h141 == _GEN_13735 ? 1'h0 : valid_321_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_837 = 9'h142 == _GEN_13735 ? 1'h0 : valid_322_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_838 = 9'h143 == _GEN_13735 ? 1'h0 : valid_323_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_839 = 9'h144 == _GEN_13735 ? 1'h0 : valid_324_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_840 = 9'h145 == _GEN_13735 ? 1'h0 : valid_325_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_841 = 9'h146 == _GEN_13735 ? 1'h0 : valid_326_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_842 = 9'h147 == _GEN_13735 ? 1'h0 : valid_327_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_843 = 9'h148 == _GEN_13735 ? 1'h0 : valid_328_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_844 = 9'h149 == _GEN_13735 ? 1'h0 : valid_329_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_845 = 9'h14a == _GEN_13735 ? 1'h0 : valid_330_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_846 = 9'h14b == _GEN_13735 ? 1'h0 : valid_331_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_847 = 9'h14c == _GEN_13735 ? 1'h0 : valid_332_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_848 = 9'h14d == _GEN_13735 ? 1'h0 : valid_333_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_849 = 9'h14e == _GEN_13735 ? 1'h0 : valid_334_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_850 = 9'h14f == _GEN_13735 ? 1'h0 : valid_335_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_851 = 9'h150 == _GEN_13735 ? 1'h0 : valid_336_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_852 = 9'h151 == _GEN_13735 ? 1'h0 : valid_337_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_853 = 9'h152 == _GEN_13735 ? 1'h0 : valid_338_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_854 = 9'h153 == _GEN_13735 ? 1'h0 : valid_339_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_855 = 9'h154 == _GEN_13735 ? 1'h0 : valid_340_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_856 = 9'h155 == _GEN_13735 ? 1'h0 : valid_341_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_857 = 9'h156 == _GEN_13735 ? 1'h0 : valid_342_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_858 = 9'h157 == _GEN_13735 ? 1'h0 : valid_343_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_859 = 9'h158 == _GEN_13735 ? 1'h0 : valid_344_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_860 = 9'h159 == _GEN_13735 ? 1'h0 : valid_345_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_861 = 9'h15a == _GEN_13735 ? 1'h0 : valid_346_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_862 = 9'h15b == _GEN_13735 ? 1'h0 : valid_347_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_863 = 9'h15c == _GEN_13735 ? 1'h0 : valid_348_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_864 = 9'h15d == _GEN_13735 ? 1'h0 : valid_349_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_865 = 9'h15e == _GEN_13735 ? 1'h0 : valid_350_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_866 = 9'h15f == _GEN_13735 ? 1'h0 : valid_351_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_867 = 9'h160 == _GEN_13735 ? 1'h0 : valid_352_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_868 = 9'h161 == _GEN_13735 ? 1'h0 : valid_353_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_869 = 9'h162 == _GEN_13735 ? 1'h0 : valid_354_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_870 = 9'h163 == _GEN_13735 ? 1'h0 : valid_355_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_871 = 9'h164 == _GEN_13735 ? 1'h0 : valid_356_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_872 = 9'h165 == _GEN_13735 ? 1'h0 : valid_357_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_873 = 9'h166 == _GEN_13735 ? 1'h0 : valid_358_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_874 = 9'h167 == _GEN_13735 ? 1'h0 : valid_359_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_875 = 9'h168 == _GEN_13735 ? 1'h0 : valid_360_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_876 = 9'h169 == _GEN_13735 ? 1'h0 : valid_361_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_877 = 9'h16a == _GEN_13735 ? 1'h0 : valid_362_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_878 = 9'h16b == _GEN_13735 ? 1'h0 : valid_363_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_879 = 9'h16c == _GEN_13735 ? 1'h0 : valid_364_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_880 = 9'h16d == _GEN_13735 ? 1'h0 : valid_365_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_881 = 9'h16e == _GEN_13735 ? 1'h0 : valid_366_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_882 = 9'h16f == _GEN_13735 ? 1'h0 : valid_367_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_883 = 9'h170 == _GEN_13735 ? 1'h0 : valid_368_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_884 = 9'h171 == _GEN_13735 ? 1'h0 : valid_369_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_885 = 9'h172 == _GEN_13735 ? 1'h0 : valid_370_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_886 = 9'h173 == _GEN_13735 ? 1'h0 : valid_371_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_887 = 9'h174 == _GEN_13735 ? 1'h0 : valid_372_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_888 = 9'h175 == _GEN_13735 ? 1'h0 : valid_373_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_889 = 9'h176 == _GEN_13735 ? 1'h0 : valid_374_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_890 = 9'h177 == _GEN_13735 ? 1'h0 : valid_375_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_891 = 9'h178 == _GEN_13735 ? 1'h0 : valid_376_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_892 = 9'h179 == _GEN_13735 ? 1'h0 : valid_377_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_893 = 9'h17a == _GEN_13735 ? 1'h0 : valid_378_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_894 = 9'h17b == _GEN_13735 ? 1'h0 : valid_379_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_895 = 9'h17c == _GEN_13735 ? 1'h0 : valid_380_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_896 = 9'h17d == _GEN_13735 ? 1'h0 : valid_381_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_897 = 9'h17e == _GEN_13735 ? 1'h0 : valid_382_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_898 = 9'h17f == _GEN_13735 ? 1'h0 : valid_383_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_899 = 9'h180 == _GEN_13735 ? 1'h0 : valid_384_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_900 = 9'h181 == _GEN_13735 ? 1'h0 : valid_385_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_901 = 9'h182 == _GEN_13735 ? 1'h0 : valid_386_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_902 = 9'h183 == _GEN_13735 ? 1'h0 : valid_387_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_903 = 9'h184 == _GEN_13735 ? 1'h0 : valid_388_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_904 = 9'h185 == _GEN_13735 ? 1'h0 : valid_389_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_905 = 9'h186 == _GEN_13735 ? 1'h0 : valid_390_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_906 = 9'h187 == _GEN_13735 ? 1'h0 : valid_391_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_907 = 9'h188 == _GEN_13735 ? 1'h0 : valid_392_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_908 = 9'h189 == _GEN_13735 ? 1'h0 : valid_393_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_909 = 9'h18a == _GEN_13735 ? 1'h0 : valid_394_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_910 = 9'h18b == _GEN_13735 ? 1'h0 : valid_395_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_911 = 9'h18c == _GEN_13735 ? 1'h0 : valid_396_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_912 = 9'h18d == _GEN_13735 ? 1'h0 : valid_397_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_913 = 9'h18e == _GEN_13735 ? 1'h0 : valid_398_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_914 = 9'h18f == _GEN_13735 ? 1'h0 : valid_399_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_915 = 9'h190 == _GEN_13735 ? 1'h0 : valid_400_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_916 = 9'h191 == _GEN_13735 ? 1'h0 : valid_401_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_917 = 9'h192 == _GEN_13735 ? 1'h0 : valid_402_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_918 = 9'h193 == _GEN_13735 ? 1'h0 : valid_403_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_919 = 9'h194 == _GEN_13735 ? 1'h0 : valid_404_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_920 = 9'h195 == _GEN_13735 ? 1'h0 : valid_405_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_921 = 9'h196 == _GEN_13735 ? 1'h0 : valid_406_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_922 = 9'h197 == _GEN_13735 ? 1'h0 : valid_407_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_923 = 9'h198 == _GEN_13735 ? 1'h0 : valid_408_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_924 = 9'h199 == _GEN_13735 ? 1'h0 : valid_409_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_925 = 9'h19a == _GEN_13735 ? 1'h0 : valid_410_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_926 = 9'h19b == _GEN_13735 ? 1'h0 : valid_411_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_927 = 9'h19c == _GEN_13735 ? 1'h0 : valid_412_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_928 = 9'h19d == _GEN_13735 ? 1'h0 : valid_413_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_929 = 9'h19e == _GEN_13735 ? 1'h0 : valid_414_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_930 = 9'h19f == _GEN_13735 ? 1'h0 : valid_415_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_931 = 9'h1a0 == _GEN_13735 ? 1'h0 : valid_416_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_932 = 9'h1a1 == _GEN_13735 ? 1'h0 : valid_417_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_933 = 9'h1a2 == _GEN_13735 ? 1'h0 : valid_418_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_934 = 9'h1a3 == _GEN_13735 ? 1'h0 : valid_419_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_935 = 9'h1a4 == _GEN_13735 ? 1'h0 : valid_420_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_936 = 9'h1a5 == _GEN_13735 ? 1'h0 : valid_421_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_937 = 9'h1a6 == _GEN_13735 ? 1'h0 : valid_422_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_938 = 9'h1a7 == _GEN_13735 ? 1'h0 : valid_423_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_939 = 9'h1a8 == _GEN_13735 ? 1'h0 : valid_424_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_940 = 9'h1a9 == _GEN_13735 ? 1'h0 : valid_425_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_941 = 9'h1aa == _GEN_13735 ? 1'h0 : valid_426_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_942 = 9'h1ab == _GEN_13735 ? 1'h0 : valid_427_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_943 = 9'h1ac == _GEN_13735 ? 1'h0 : valid_428_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_944 = 9'h1ad == _GEN_13735 ? 1'h0 : valid_429_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_945 = 9'h1ae == _GEN_13735 ? 1'h0 : valid_430_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_946 = 9'h1af == _GEN_13735 ? 1'h0 : valid_431_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_947 = 9'h1b0 == _GEN_13735 ? 1'h0 : valid_432_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_948 = 9'h1b1 == _GEN_13735 ? 1'h0 : valid_433_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_949 = 9'h1b2 == _GEN_13735 ? 1'h0 : valid_434_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_950 = 9'h1b3 == _GEN_13735 ? 1'h0 : valid_435_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_951 = 9'h1b4 == _GEN_13735 ? 1'h0 : valid_436_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_952 = 9'h1b5 == _GEN_13735 ? 1'h0 : valid_437_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_953 = 9'h1b6 == _GEN_13735 ? 1'h0 : valid_438_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_954 = 9'h1b7 == _GEN_13735 ? 1'h0 : valid_439_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_955 = 9'h1b8 == _GEN_13735 ? 1'h0 : valid_440_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_956 = 9'h1b9 == _GEN_13735 ? 1'h0 : valid_441_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_957 = 9'h1ba == _GEN_13735 ? 1'h0 : valid_442_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_958 = 9'h1bb == _GEN_13735 ? 1'h0 : valid_443_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_959 = 9'h1bc == _GEN_13735 ? 1'h0 : valid_444_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_960 = 9'h1bd == _GEN_13735 ? 1'h0 : valid_445_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_961 = 9'h1be == _GEN_13735 ? 1'h0 : valid_446_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_962 = 9'h1bf == _GEN_13735 ? 1'h0 : valid_447_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_963 = 9'h1c0 == _GEN_13735 ? 1'h0 : valid_448_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_964 = 9'h1c1 == _GEN_13735 ? 1'h0 : valid_449_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_965 = 9'h1c2 == _GEN_13735 ? 1'h0 : valid_450_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_966 = 9'h1c3 == _GEN_13735 ? 1'h0 : valid_451_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_967 = 9'h1c4 == _GEN_13735 ? 1'h0 : valid_452_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_968 = 9'h1c5 == _GEN_13735 ? 1'h0 : valid_453_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_969 = 9'h1c6 == _GEN_13735 ? 1'h0 : valid_454_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_970 = 9'h1c7 == _GEN_13735 ? 1'h0 : valid_455_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_971 = 9'h1c8 == _GEN_13735 ? 1'h0 : valid_456_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_972 = 9'h1c9 == _GEN_13735 ? 1'h0 : valid_457_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_973 = 9'h1ca == _GEN_13735 ? 1'h0 : valid_458_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_974 = 9'h1cb == _GEN_13735 ? 1'h0 : valid_459_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_975 = 9'h1cc == _GEN_13735 ? 1'h0 : valid_460_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_976 = 9'h1cd == _GEN_13735 ? 1'h0 : valid_461_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_977 = 9'h1ce == _GEN_13735 ? 1'h0 : valid_462_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_978 = 9'h1cf == _GEN_13735 ? 1'h0 : valid_463_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_979 = 9'h1d0 == _GEN_13735 ? 1'h0 : valid_464_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_980 = 9'h1d1 == _GEN_13735 ? 1'h0 : valid_465_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_981 = 9'h1d2 == _GEN_13735 ? 1'h0 : valid_466_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_982 = 9'h1d3 == _GEN_13735 ? 1'h0 : valid_467_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_983 = 9'h1d4 == _GEN_13735 ? 1'h0 : valid_468_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_984 = 9'h1d5 == _GEN_13735 ? 1'h0 : valid_469_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_985 = 9'h1d6 == _GEN_13735 ? 1'h0 : valid_470_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_986 = 9'h1d7 == _GEN_13735 ? 1'h0 : valid_471_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_987 = 9'h1d8 == _GEN_13735 ? 1'h0 : valid_472_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_988 = 9'h1d9 == _GEN_13735 ? 1'h0 : valid_473_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_989 = 9'h1da == _GEN_13735 ? 1'h0 : valid_474_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_990 = 9'h1db == _GEN_13735 ? 1'h0 : valid_475_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_991 = 9'h1dc == _GEN_13735 ? 1'h0 : valid_476_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_992 = 9'h1dd == _GEN_13735 ? 1'h0 : valid_477_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_993 = 9'h1de == _GEN_13735 ? 1'h0 : valid_478_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_994 = 9'h1df == _GEN_13735 ? 1'h0 : valid_479_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_995 = 9'h1e0 == _GEN_13735 ? 1'h0 : valid_480_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_996 = 9'h1e1 == _GEN_13735 ? 1'h0 : valid_481_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_997 = 9'h1e2 == _GEN_13735 ? 1'h0 : valid_482_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_998 = 9'h1e3 == _GEN_13735 ? 1'h0 : valid_483_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_999 = 9'h1e4 == _GEN_13735 ? 1'h0 : valid_484_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1000 = 9'h1e5 == _GEN_13735 ? 1'h0 : valid_485_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1001 = 9'h1e6 == _GEN_13735 ? 1'h0 : valid_486_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1002 = 9'h1e7 == _GEN_13735 ? 1'h0 : valid_487_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1003 = 9'h1e8 == _GEN_13735 ? 1'h0 : valid_488_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1004 = 9'h1e9 == _GEN_13735 ? 1'h0 : valid_489_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1005 = 9'h1ea == _GEN_13735 ? 1'h0 : valid_490_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1006 = 9'h1eb == _GEN_13735 ? 1'h0 : valid_491_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1007 = 9'h1ec == _GEN_13735 ? 1'h0 : valid_492_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1008 = 9'h1ed == _GEN_13735 ? 1'h0 : valid_493_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1009 = 9'h1ee == _GEN_13735 ? 1'h0 : valid_494_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1010 = 9'h1ef == _GEN_13735 ? 1'h0 : valid_495_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1011 = 9'h1f0 == _GEN_13735 ? 1'h0 : valid_496_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1012 = 9'h1f1 == _GEN_13735 ? 1'h0 : valid_497_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1013 = 9'h1f2 == _GEN_13735 ? 1'h0 : valid_498_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1014 = 9'h1f3 == _GEN_13735 ? 1'h0 : valid_499_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1015 = 9'h1f4 == _GEN_13735 ? 1'h0 : valid_500_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1016 = 9'h1f5 == _GEN_13735 ? 1'h0 : valid_501_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1017 = 9'h1f6 == _GEN_13735 ? 1'h0 : valid_502_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1018 = 9'h1f7 == _GEN_13735 ? 1'h0 : valid_503_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1019 = 9'h1f8 == _GEN_13735 ? 1'h0 : valid_504_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1020 = 9'h1f9 == _GEN_13735 ? 1'h0 : valid_505_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1021 = 9'h1fa == _GEN_13735 ? 1'h0 : valid_506_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1022 = 9'h1fb == _GEN_13735 ? 1'h0 : valid_507_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1023 = 9'h1fc == _GEN_13735 ? 1'h0 : valid_508_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1024 = 9'h1fd == _GEN_13735 ? 1'h0 : valid_509_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1025 = 9'h1fe == _GEN_13735 ? 1'h0 : valid_510_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1026 = 9'h1ff == _GEN_13735 ? 1'h0 : valid_511_1; // @[ICache.scala 52:22 89:{24,24}]
  wire  _GEN_1027 = io_cpu_fence_value & _T & _T_2 ? _GEN_3 : valid_0_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1028 = io_cpu_fence_value & _T & _T_2 ? _GEN_4 : valid_1_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1029 = io_cpu_fence_value & _T & _T_2 ? _GEN_5 : valid_2_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1030 = io_cpu_fence_value & _T & _T_2 ? _GEN_6 : valid_3_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1031 = io_cpu_fence_value & _T & _T_2 ? _GEN_7 : valid_4_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1032 = io_cpu_fence_value & _T & _T_2 ? _GEN_8 : valid_5_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1033 = io_cpu_fence_value & _T & _T_2 ? _GEN_9 : valid_6_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1034 = io_cpu_fence_value & _T & _T_2 ? _GEN_10 : valid_7_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1035 = io_cpu_fence_value & _T & _T_2 ? _GEN_11 : valid_8_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1036 = io_cpu_fence_value & _T & _T_2 ? _GEN_12 : valid_9_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1037 = io_cpu_fence_value & _T & _T_2 ? _GEN_13 : valid_10_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1038 = io_cpu_fence_value & _T & _T_2 ? _GEN_14 : valid_11_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1039 = io_cpu_fence_value & _T & _T_2 ? _GEN_15 : valid_12_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1040 = io_cpu_fence_value & _T & _T_2 ? _GEN_16 : valid_13_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1041 = io_cpu_fence_value & _T & _T_2 ? _GEN_17 : valid_14_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1042 = io_cpu_fence_value & _T & _T_2 ? _GEN_18 : valid_15_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1043 = io_cpu_fence_value & _T & _T_2 ? _GEN_19 : valid_16_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1044 = io_cpu_fence_value & _T & _T_2 ? _GEN_20 : valid_17_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1045 = io_cpu_fence_value & _T & _T_2 ? _GEN_21 : valid_18_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1046 = io_cpu_fence_value & _T & _T_2 ? _GEN_22 : valid_19_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1047 = io_cpu_fence_value & _T & _T_2 ? _GEN_23 : valid_20_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1048 = io_cpu_fence_value & _T & _T_2 ? _GEN_24 : valid_21_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1049 = io_cpu_fence_value & _T & _T_2 ? _GEN_25 : valid_22_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1050 = io_cpu_fence_value & _T & _T_2 ? _GEN_26 : valid_23_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1051 = io_cpu_fence_value & _T & _T_2 ? _GEN_27 : valid_24_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1052 = io_cpu_fence_value & _T & _T_2 ? _GEN_28 : valid_25_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1053 = io_cpu_fence_value & _T & _T_2 ? _GEN_29 : valid_26_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1054 = io_cpu_fence_value & _T & _T_2 ? _GEN_30 : valid_27_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1055 = io_cpu_fence_value & _T & _T_2 ? _GEN_31 : valid_28_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1056 = io_cpu_fence_value & _T & _T_2 ? _GEN_32 : valid_29_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1057 = io_cpu_fence_value & _T & _T_2 ? _GEN_33 : valid_30_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1058 = io_cpu_fence_value & _T & _T_2 ? _GEN_34 : valid_31_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1059 = io_cpu_fence_value & _T & _T_2 ? _GEN_35 : valid_32_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1060 = io_cpu_fence_value & _T & _T_2 ? _GEN_36 : valid_33_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1061 = io_cpu_fence_value & _T & _T_2 ? _GEN_37 : valid_34_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1062 = io_cpu_fence_value & _T & _T_2 ? _GEN_38 : valid_35_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1063 = io_cpu_fence_value & _T & _T_2 ? _GEN_39 : valid_36_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1064 = io_cpu_fence_value & _T & _T_2 ? _GEN_40 : valid_37_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1065 = io_cpu_fence_value & _T & _T_2 ? _GEN_41 : valid_38_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1066 = io_cpu_fence_value & _T & _T_2 ? _GEN_42 : valid_39_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1067 = io_cpu_fence_value & _T & _T_2 ? _GEN_43 : valid_40_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1068 = io_cpu_fence_value & _T & _T_2 ? _GEN_44 : valid_41_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1069 = io_cpu_fence_value & _T & _T_2 ? _GEN_45 : valid_42_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1070 = io_cpu_fence_value & _T & _T_2 ? _GEN_46 : valid_43_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1071 = io_cpu_fence_value & _T & _T_2 ? _GEN_47 : valid_44_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1072 = io_cpu_fence_value & _T & _T_2 ? _GEN_48 : valid_45_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1073 = io_cpu_fence_value & _T & _T_2 ? _GEN_49 : valid_46_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1074 = io_cpu_fence_value & _T & _T_2 ? _GEN_50 : valid_47_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1075 = io_cpu_fence_value & _T & _T_2 ? _GEN_51 : valid_48_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1076 = io_cpu_fence_value & _T & _T_2 ? _GEN_52 : valid_49_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1077 = io_cpu_fence_value & _T & _T_2 ? _GEN_53 : valid_50_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1078 = io_cpu_fence_value & _T & _T_2 ? _GEN_54 : valid_51_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1079 = io_cpu_fence_value & _T & _T_2 ? _GEN_55 : valid_52_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1080 = io_cpu_fence_value & _T & _T_2 ? _GEN_56 : valid_53_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1081 = io_cpu_fence_value & _T & _T_2 ? _GEN_57 : valid_54_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1082 = io_cpu_fence_value & _T & _T_2 ? _GEN_58 : valid_55_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1083 = io_cpu_fence_value & _T & _T_2 ? _GEN_59 : valid_56_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1084 = io_cpu_fence_value & _T & _T_2 ? _GEN_60 : valid_57_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1085 = io_cpu_fence_value & _T & _T_2 ? _GEN_61 : valid_58_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1086 = io_cpu_fence_value & _T & _T_2 ? _GEN_62 : valid_59_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1087 = io_cpu_fence_value & _T & _T_2 ? _GEN_63 : valid_60_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1088 = io_cpu_fence_value & _T & _T_2 ? _GEN_64 : valid_61_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1089 = io_cpu_fence_value & _T & _T_2 ? _GEN_65 : valid_62_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1090 = io_cpu_fence_value & _T & _T_2 ? _GEN_66 : valid_63_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1091 = io_cpu_fence_value & _T & _T_2 ? _GEN_67 : valid_64_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1092 = io_cpu_fence_value & _T & _T_2 ? _GEN_68 : valid_65_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1093 = io_cpu_fence_value & _T & _T_2 ? _GEN_69 : valid_66_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1094 = io_cpu_fence_value & _T & _T_2 ? _GEN_70 : valid_67_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1095 = io_cpu_fence_value & _T & _T_2 ? _GEN_71 : valid_68_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1096 = io_cpu_fence_value & _T & _T_2 ? _GEN_72 : valid_69_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1097 = io_cpu_fence_value & _T & _T_2 ? _GEN_73 : valid_70_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1098 = io_cpu_fence_value & _T & _T_2 ? _GEN_74 : valid_71_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1099 = io_cpu_fence_value & _T & _T_2 ? _GEN_75 : valid_72_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1100 = io_cpu_fence_value & _T & _T_2 ? _GEN_76 : valid_73_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1101 = io_cpu_fence_value & _T & _T_2 ? _GEN_77 : valid_74_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1102 = io_cpu_fence_value & _T & _T_2 ? _GEN_78 : valid_75_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1103 = io_cpu_fence_value & _T & _T_2 ? _GEN_79 : valid_76_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1104 = io_cpu_fence_value & _T & _T_2 ? _GEN_80 : valid_77_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1105 = io_cpu_fence_value & _T & _T_2 ? _GEN_81 : valid_78_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1106 = io_cpu_fence_value & _T & _T_2 ? _GEN_82 : valid_79_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1107 = io_cpu_fence_value & _T & _T_2 ? _GEN_83 : valid_80_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1108 = io_cpu_fence_value & _T & _T_2 ? _GEN_84 : valid_81_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1109 = io_cpu_fence_value & _T & _T_2 ? _GEN_85 : valid_82_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1110 = io_cpu_fence_value & _T & _T_2 ? _GEN_86 : valid_83_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1111 = io_cpu_fence_value & _T & _T_2 ? _GEN_87 : valid_84_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1112 = io_cpu_fence_value & _T & _T_2 ? _GEN_88 : valid_85_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1113 = io_cpu_fence_value & _T & _T_2 ? _GEN_89 : valid_86_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1114 = io_cpu_fence_value & _T & _T_2 ? _GEN_90 : valid_87_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1115 = io_cpu_fence_value & _T & _T_2 ? _GEN_91 : valid_88_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1116 = io_cpu_fence_value & _T & _T_2 ? _GEN_92 : valid_89_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1117 = io_cpu_fence_value & _T & _T_2 ? _GEN_93 : valid_90_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1118 = io_cpu_fence_value & _T & _T_2 ? _GEN_94 : valid_91_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1119 = io_cpu_fence_value & _T & _T_2 ? _GEN_95 : valid_92_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1120 = io_cpu_fence_value & _T & _T_2 ? _GEN_96 : valid_93_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1121 = io_cpu_fence_value & _T & _T_2 ? _GEN_97 : valid_94_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1122 = io_cpu_fence_value & _T & _T_2 ? _GEN_98 : valid_95_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1123 = io_cpu_fence_value & _T & _T_2 ? _GEN_99 : valid_96_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1124 = io_cpu_fence_value & _T & _T_2 ? _GEN_100 : valid_97_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1125 = io_cpu_fence_value & _T & _T_2 ? _GEN_101 : valid_98_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1126 = io_cpu_fence_value & _T & _T_2 ? _GEN_102 : valid_99_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1127 = io_cpu_fence_value & _T & _T_2 ? _GEN_103 : valid_100_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1128 = io_cpu_fence_value & _T & _T_2 ? _GEN_104 : valid_101_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1129 = io_cpu_fence_value & _T & _T_2 ? _GEN_105 : valid_102_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1130 = io_cpu_fence_value & _T & _T_2 ? _GEN_106 : valid_103_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1131 = io_cpu_fence_value & _T & _T_2 ? _GEN_107 : valid_104_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1132 = io_cpu_fence_value & _T & _T_2 ? _GEN_108 : valid_105_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1133 = io_cpu_fence_value & _T & _T_2 ? _GEN_109 : valid_106_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1134 = io_cpu_fence_value & _T & _T_2 ? _GEN_110 : valid_107_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1135 = io_cpu_fence_value & _T & _T_2 ? _GEN_111 : valid_108_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1136 = io_cpu_fence_value & _T & _T_2 ? _GEN_112 : valid_109_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1137 = io_cpu_fence_value & _T & _T_2 ? _GEN_113 : valid_110_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1138 = io_cpu_fence_value & _T & _T_2 ? _GEN_114 : valid_111_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1139 = io_cpu_fence_value & _T & _T_2 ? _GEN_115 : valid_112_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1140 = io_cpu_fence_value & _T & _T_2 ? _GEN_116 : valid_113_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1141 = io_cpu_fence_value & _T & _T_2 ? _GEN_117 : valid_114_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1142 = io_cpu_fence_value & _T & _T_2 ? _GEN_118 : valid_115_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1143 = io_cpu_fence_value & _T & _T_2 ? _GEN_119 : valid_116_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1144 = io_cpu_fence_value & _T & _T_2 ? _GEN_120 : valid_117_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1145 = io_cpu_fence_value & _T & _T_2 ? _GEN_121 : valid_118_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1146 = io_cpu_fence_value & _T & _T_2 ? _GEN_122 : valid_119_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1147 = io_cpu_fence_value & _T & _T_2 ? _GEN_123 : valid_120_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1148 = io_cpu_fence_value & _T & _T_2 ? _GEN_124 : valid_121_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1149 = io_cpu_fence_value & _T & _T_2 ? _GEN_125 : valid_122_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1150 = io_cpu_fence_value & _T & _T_2 ? _GEN_126 : valid_123_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1151 = io_cpu_fence_value & _T & _T_2 ? _GEN_127 : valid_124_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1152 = io_cpu_fence_value & _T & _T_2 ? _GEN_128 : valid_125_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1153 = io_cpu_fence_value & _T & _T_2 ? _GEN_129 : valid_126_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1154 = io_cpu_fence_value & _T & _T_2 ? _GEN_130 : valid_127_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1155 = io_cpu_fence_value & _T & _T_2 ? _GEN_131 : valid_128_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1156 = io_cpu_fence_value & _T & _T_2 ? _GEN_132 : valid_129_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1157 = io_cpu_fence_value & _T & _T_2 ? _GEN_133 : valid_130_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1158 = io_cpu_fence_value & _T & _T_2 ? _GEN_134 : valid_131_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1159 = io_cpu_fence_value & _T & _T_2 ? _GEN_135 : valid_132_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1160 = io_cpu_fence_value & _T & _T_2 ? _GEN_136 : valid_133_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1161 = io_cpu_fence_value & _T & _T_2 ? _GEN_137 : valid_134_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1162 = io_cpu_fence_value & _T & _T_2 ? _GEN_138 : valid_135_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1163 = io_cpu_fence_value & _T & _T_2 ? _GEN_139 : valid_136_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1164 = io_cpu_fence_value & _T & _T_2 ? _GEN_140 : valid_137_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1165 = io_cpu_fence_value & _T & _T_2 ? _GEN_141 : valid_138_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1166 = io_cpu_fence_value & _T & _T_2 ? _GEN_142 : valid_139_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1167 = io_cpu_fence_value & _T & _T_2 ? _GEN_143 : valid_140_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1168 = io_cpu_fence_value & _T & _T_2 ? _GEN_144 : valid_141_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1169 = io_cpu_fence_value & _T & _T_2 ? _GEN_145 : valid_142_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1170 = io_cpu_fence_value & _T & _T_2 ? _GEN_146 : valid_143_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1171 = io_cpu_fence_value & _T & _T_2 ? _GEN_147 : valid_144_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1172 = io_cpu_fence_value & _T & _T_2 ? _GEN_148 : valid_145_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1173 = io_cpu_fence_value & _T & _T_2 ? _GEN_149 : valid_146_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1174 = io_cpu_fence_value & _T & _T_2 ? _GEN_150 : valid_147_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1175 = io_cpu_fence_value & _T & _T_2 ? _GEN_151 : valid_148_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1176 = io_cpu_fence_value & _T & _T_2 ? _GEN_152 : valid_149_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1177 = io_cpu_fence_value & _T & _T_2 ? _GEN_153 : valid_150_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1178 = io_cpu_fence_value & _T & _T_2 ? _GEN_154 : valid_151_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1179 = io_cpu_fence_value & _T & _T_2 ? _GEN_155 : valid_152_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1180 = io_cpu_fence_value & _T & _T_2 ? _GEN_156 : valid_153_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1181 = io_cpu_fence_value & _T & _T_2 ? _GEN_157 : valid_154_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1182 = io_cpu_fence_value & _T & _T_2 ? _GEN_158 : valid_155_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1183 = io_cpu_fence_value & _T & _T_2 ? _GEN_159 : valid_156_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1184 = io_cpu_fence_value & _T & _T_2 ? _GEN_160 : valid_157_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1185 = io_cpu_fence_value & _T & _T_2 ? _GEN_161 : valid_158_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1186 = io_cpu_fence_value & _T & _T_2 ? _GEN_162 : valid_159_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1187 = io_cpu_fence_value & _T & _T_2 ? _GEN_163 : valid_160_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1188 = io_cpu_fence_value & _T & _T_2 ? _GEN_164 : valid_161_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1189 = io_cpu_fence_value & _T & _T_2 ? _GEN_165 : valid_162_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1190 = io_cpu_fence_value & _T & _T_2 ? _GEN_166 : valid_163_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1191 = io_cpu_fence_value & _T & _T_2 ? _GEN_167 : valid_164_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1192 = io_cpu_fence_value & _T & _T_2 ? _GEN_168 : valid_165_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1193 = io_cpu_fence_value & _T & _T_2 ? _GEN_169 : valid_166_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1194 = io_cpu_fence_value & _T & _T_2 ? _GEN_170 : valid_167_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1195 = io_cpu_fence_value & _T & _T_2 ? _GEN_171 : valid_168_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1196 = io_cpu_fence_value & _T & _T_2 ? _GEN_172 : valid_169_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1197 = io_cpu_fence_value & _T & _T_2 ? _GEN_173 : valid_170_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1198 = io_cpu_fence_value & _T & _T_2 ? _GEN_174 : valid_171_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1199 = io_cpu_fence_value & _T & _T_2 ? _GEN_175 : valid_172_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1200 = io_cpu_fence_value & _T & _T_2 ? _GEN_176 : valid_173_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1201 = io_cpu_fence_value & _T & _T_2 ? _GEN_177 : valid_174_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1202 = io_cpu_fence_value & _T & _T_2 ? _GEN_178 : valid_175_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1203 = io_cpu_fence_value & _T & _T_2 ? _GEN_179 : valid_176_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1204 = io_cpu_fence_value & _T & _T_2 ? _GEN_180 : valid_177_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1205 = io_cpu_fence_value & _T & _T_2 ? _GEN_181 : valid_178_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1206 = io_cpu_fence_value & _T & _T_2 ? _GEN_182 : valid_179_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1207 = io_cpu_fence_value & _T & _T_2 ? _GEN_183 : valid_180_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1208 = io_cpu_fence_value & _T & _T_2 ? _GEN_184 : valid_181_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1209 = io_cpu_fence_value & _T & _T_2 ? _GEN_185 : valid_182_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1210 = io_cpu_fence_value & _T & _T_2 ? _GEN_186 : valid_183_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1211 = io_cpu_fence_value & _T & _T_2 ? _GEN_187 : valid_184_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1212 = io_cpu_fence_value & _T & _T_2 ? _GEN_188 : valid_185_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1213 = io_cpu_fence_value & _T & _T_2 ? _GEN_189 : valid_186_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1214 = io_cpu_fence_value & _T & _T_2 ? _GEN_190 : valid_187_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1215 = io_cpu_fence_value & _T & _T_2 ? _GEN_191 : valid_188_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1216 = io_cpu_fence_value & _T & _T_2 ? _GEN_192 : valid_189_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1217 = io_cpu_fence_value & _T & _T_2 ? _GEN_193 : valid_190_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1218 = io_cpu_fence_value & _T & _T_2 ? _GEN_194 : valid_191_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1219 = io_cpu_fence_value & _T & _T_2 ? _GEN_195 : valid_192_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1220 = io_cpu_fence_value & _T & _T_2 ? _GEN_196 : valid_193_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1221 = io_cpu_fence_value & _T & _T_2 ? _GEN_197 : valid_194_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1222 = io_cpu_fence_value & _T & _T_2 ? _GEN_198 : valid_195_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1223 = io_cpu_fence_value & _T & _T_2 ? _GEN_199 : valid_196_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1224 = io_cpu_fence_value & _T & _T_2 ? _GEN_200 : valid_197_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1225 = io_cpu_fence_value & _T & _T_2 ? _GEN_201 : valid_198_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1226 = io_cpu_fence_value & _T & _T_2 ? _GEN_202 : valid_199_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1227 = io_cpu_fence_value & _T & _T_2 ? _GEN_203 : valid_200_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1228 = io_cpu_fence_value & _T & _T_2 ? _GEN_204 : valid_201_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1229 = io_cpu_fence_value & _T & _T_2 ? _GEN_205 : valid_202_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1230 = io_cpu_fence_value & _T & _T_2 ? _GEN_206 : valid_203_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1231 = io_cpu_fence_value & _T & _T_2 ? _GEN_207 : valid_204_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1232 = io_cpu_fence_value & _T & _T_2 ? _GEN_208 : valid_205_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1233 = io_cpu_fence_value & _T & _T_2 ? _GEN_209 : valid_206_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1234 = io_cpu_fence_value & _T & _T_2 ? _GEN_210 : valid_207_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1235 = io_cpu_fence_value & _T & _T_2 ? _GEN_211 : valid_208_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1236 = io_cpu_fence_value & _T & _T_2 ? _GEN_212 : valid_209_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1237 = io_cpu_fence_value & _T & _T_2 ? _GEN_213 : valid_210_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1238 = io_cpu_fence_value & _T & _T_2 ? _GEN_214 : valid_211_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1239 = io_cpu_fence_value & _T & _T_2 ? _GEN_215 : valid_212_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1240 = io_cpu_fence_value & _T & _T_2 ? _GEN_216 : valid_213_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1241 = io_cpu_fence_value & _T & _T_2 ? _GEN_217 : valid_214_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1242 = io_cpu_fence_value & _T & _T_2 ? _GEN_218 : valid_215_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1243 = io_cpu_fence_value & _T & _T_2 ? _GEN_219 : valid_216_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1244 = io_cpu_fence_value & _T & _T_2 ? _GEN_220 : valid_217_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1245 = io_cpu_fence_value & _T & _T_2 ? _GEN_221 : valid_218_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1246 = io_cpu_fence_value & _T & _T_2 ? _GEN_222 : valid_219_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1247 = io_cpu_fence_value & _T & _T_2 ? _GEN_223 : valid_220_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1248 = io_cpu_fence_value & _T & _T_2 ? _GEN_224 : valid_221_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1249 = io_cpu_fence_value & _T & _T_2 ? _GEN_225 : valid_222_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1250 = io_cpu_fence_value & _T & _T_2 ? _GEN_226 : valid_223_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1251 = io_cpu_fence_value & _T & _T_2 ? _GEN_227 : valid_224_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1252 = io_cpu_fence_value & _T & _T_2 ? _GEN_228 : valid_225_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1253 = io_cpu_fence_value & _T & _T_2 ? _GEN_229 : valid_226_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1254 = io_cpu_fence_value & _T & _T_2 ? _GEN_230 : valid_227_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1255 = io_cpu_fence_value & _T & _T_2 ? _GEN_231 : valid_228_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1256 = io_cpu_fence_value & _T & _T_2 ? _GEN_232 : valid_229_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1257 = io_cpu_fence_value & _T & _T_2 ? _GEN_233 : valid_230_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1258 = io_cpu_fence_value & _T & _T_2 ? _GEN_234 : valid_231_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1259 = io_cpu_fence_value & _T & _T_2 ? _GEN_235 : valid_232_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1260 = io_cpu_fence_value & _T & _T_2 ? _GEN_236 : valid_233_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1261 = io_cpu_fence_value & _T & _T_2 ? _GEN_237 : valid_234_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1262 = io_cpu_fence_value & _T & _T_2 ? _GEN_238 : valid_235_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1263 = io_cpu_fence_value & _T & _T_2 ? _GEN_239 : valid_236_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1264 = io_cpu_fence_value & _T & _T_2 ? _GEN_240 : valid_237_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1265 = io_cpu_fence_value & _T & _T_2 ? _GEN_241 : valid_238_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1266 = io_cpu_fence_value & _T & _T_2 ? _GEN_242 : valid_239_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1267 = io_cpu_fence_value & _T & _T_2 ? _GEN_243 : valid_240_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1268 = io_cpu_fence_value & _T & _T_2 ? _GEN_244 : valid_241_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1269 = io_cpu_fence_value & _T & _T_2 ? _GEN_245 : valid_242_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1270 = io_cpu_fence_value & _T & _T_2 ? _GEN_246 : valid_243_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1271 = io_cpu_fence_value & _T & _T_2 ? _GEN_247 : valid_244_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1272 = io_cpu_fence_value & _T & _T_2 ? _GEN_248 : valid_245_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1273 = io_cpu_fence_value & _T & _T_2 ? _GEN_249 : valid_246_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1274 = io_cpu_fence_value & _T & _T_2 ? _GEN_250 : valid_247_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1275 = io_cpu_fence_value & _T & _T_2 ? _GEN_251 : valid_248_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1276 = io_cpu_fence_value & _T & _T_2 ? _GEN_252 : valid_249_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1277 = io_cpu_fence_value & _T & _T_2 ? _GEN_253 : valid_250_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1278 = io_cpu_fence_value & _T & _T_2 ? _GEN_254 : valid_251_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1279 = io_cpu_fence_value & _T & _T_2 ? _GEN_255 : valid_252_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1280 = io_cpu_fence_value & _T & _T_2 ? _GEN_256 : valid_253_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1281 = io_cpu_fence_value & _T & _T_2 ? _GEN_257 : valid_254_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1282 = io_cpu_fence_value & _T & _T_2 ? _GEN_258 : valid_255_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1283 = io_cpu_fence_value & _T & _T_2 ? _GEN_259 : valid_256_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1284 = io_cpu_fence_value & _T & _T_2 ? _GEN_260 : valid_257_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1285 = io_cpu_fence_value & _T & _T_2 ? _GEN_261 : valid_258_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1286 = io_cpu_fence_value & _T & _T_2 ? _GEN_262 : valid_259_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1287 = io_cpu_fence_value & _T & _T_2 ? _GEN_263 : valid_260_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1288 = io_cpu_fence_value & _T & _T_2 ? _GEN_264 : valid_261_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1289 = io_cpu_fence_value & _T & _T_2 ? _GEN_265 : valid_262_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1290 = io_cpu_fence_value & _T & _T_2 ? _GEN_266 : valid_263_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1291 = io_cpu_fence_value & _T & _T_2 ? _GEN_267 : valid_264_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1292 = io_cpu_fence_value & _T & _T_2 ? _GEN_268 : valid_265_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1293 = io_cpu_fence_value & _T & _T_2 ? _GEN_269 : valid_266_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1294 = io_cpu_fence_value & _T & _T_2 ? _GEN_270 : valid_267_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1295 = io_cpu_fence_value & _T & _T_2 ? _GEN_271 : valid_268_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1296 = io_cpu_fence_value & _T & _T_2 ? _GEN_272 : valid_269_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1297 = io_cpu_fence_value & _T & _T_2 ? _GEN_273 : valid_270_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1298 = io_cpu_fence_value & _T & _T_2 ? _GEN_274 : valid_271_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1299 = io_cpu_fence_value & _T & _T_2 ? _GEN_275 : valid_272_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1300 = io_cpu_fence_value & _T & _T_2 ? _GEN_276 : valid_273_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1301 = io_cpu_fence_value & _T & _T_2 ? _GEN_277 : valid_274_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1302 = io_cpu_fence_value & _T & _T_2 ? _GEN_278 : valid_275_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1303 = io_cpu_fence_value & _T & _T_2 ? _GEN_279 : valid_276_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1304 = io_cpu_fence_value & _T & _T_2 ? _GEN_280 : valid_277_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1305 = io_cpu_fence_value & _T & _T_2 ? _GEN_281 : valid_278_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1306 = io_cpu_fence_value & _T & _T_2 ? _GEN_282 : valid_279_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1307 = io_cpu_fence_value & _T & _T_2 ? _GEN_283 : valid_280_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1308 = io_cpu_fence_value & _T & _T_2 ? _GEN_284 : valid_281_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1309 = io_cpu_fence_value & _T & _T_2 ? _GEN_285 : valid_282_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1310 = io_cpu_fence_value & _T & _T_2 ? _GEN_286 : valid_283_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1311 = io_cpu_fence_value & _T & _T_2 ? _GEN_287 : valid_284_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1312 = io_cpu_fence_value & _T & _T_2 ? _GEN_288 : valid_285_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1313 = io_cpu_fence_value & _T & _T_2 ? _GEN_289 : valid_286_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1314 = io_cpu_fence_value & _T & _T_2 ? _GEN_290 : valid_287_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1315 = io_cpu_fence_value & _T & _T_2 ? _GEN_291 : valid_288_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1316 = io_cpu_fence_value & _T & _T_2 ? _GEN_292 : valid_289_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1317 = io_cpu_fence_value & _T & _T_2 ? _GEN_293 : valid_290_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1318 = io_cpu_fence_value & _T & _T_2 ? _GEN_294 : valid_291_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1319 = io_cpu_fence_value & _T & _T_2 ? _GEN_295 : valid_292_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1320 = io_cpu_fence_value & _T & _T_2 ? _GEN_296 : valid_293_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1321 = io_cpu_fence_value & _T & _T_2 ? _GEN_297 : valid_294_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1322 = io_cpu_fence_value & _T & _T_2 ? _GEN_298 : valid_295_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1323 = io_cpu_fence_value & _T & _T_2 ? _GEN_299 : valid_296_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1324 = io_cpu_fence_value & _T & _T_2 ? _GEN_300 : valid_297_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1325 = io_cpu_fence_value & _T & _T_2 ? _GEN_301 : valid_298_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1326 = io_cpu_fence_value & _T & _T_2 ? _GEN_302 : valid_299_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1327 = io_cpu_fence_value & _T & _T_2 ? _GEN_303 : valid_300_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1328 = io_cpu_fence_value & _T & _T_2 ? _GEN_304 : valid_301_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1329 = io_cpu_fence_value & _T & _T_2 ? _GEN_305 : valid_302_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1330 = io_cpu_fence_value & _T & _T_2 ? _GEN_306 : valid_303_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1331 = io_cpu_fence_value & _T & _T_2 ? _GEN_307 : valid_304_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1332 = io_cpu_fence_value & _T & _T_2 ? _GEN_308 : valid_305_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1333 = io_cpu_fence_value & _T & _T_2 ? _GEN_309 : valid_306_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1334 = io_cpu_fence_value & _T & _T_2 ? _GEN_310 : valid_307_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1335 = io_cpu_fence_value & _T & _T_2 ? _GEN_311 : valid_308_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1336 = io_cpu_fence_value & _T & _T_2 ? _GEN_312 : valid_309_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1337 = io_cpu_fence_value & _T & _T_2 ? _GEN_313 : valid_310_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1338 = io_cpu_fence_value & _T & _T_2 ? _GEN_314 : valid_311_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1339 = io_cpu_fence_value & _T & _T_2 ? _GEN_315 : valid_312_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1340 = io_cpu_fence_value & _T & _T_2 ? _GEN_316 : valid_313_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1341 = io_cpu_fence_value & _T & _T_2 ? _GEN_317 : valid_314_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1342 = io_cpu_fence_value & _T & _T_2 ? _GEN_318 : valid_315_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1343 = io_cpu_fence_value & _T & _T_2 ? _GEN_319 : valid_316_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1344 = io_cpu_fence_value & _T & _T_2 ? _GEN_320 : valid_317_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1345 = io_cpu_fence_value & _T & _T_2 ? _GEN_321 : valid_318_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1346 = io_cpu_fence_value & _T & _T_2 ? _GEN_322 : valid_319_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1347 = io_cpu_fence_value & _T & _T_2 ? _GEN_323 : valid_320_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1348 = io_cpu_fence_value & _T & _T_2 ? _GEN_324 : valid_321_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1349 = io_cpu_fence_value & _T & _T_2 ? _GEN_325 : valid_322_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1350 = io_cpu_fence_value & _T & _T_2 ? _GEN_326 : valid_323_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1351 = io_cpu_fence_value & _T & _T_2 ? _GEN_327 : valid_324_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1352 = io_cpu_fence_value & _T & _T_2 ? _GEN_328 : valid_325_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1353 = io_cpu_fence_value & _T & _T_2 ? _GEN_329 : valid_326_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1354 = io_cpu_fence_value & _T & _T_2 ? _GEN_330 : valid_327_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1355 = io_cpu_fence_value & _T & _T_2 ? _GEN_331 : valid_328_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1356 = io_cpu_fence_value & _T & _T_2 ? _GEN_332 : valid_329_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1357 = io_cpu_fence_value & _T & _T_2 ? _GEN_333 : valid_330_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1358 = io_cpu_fence_value & _T & _T_2 ? _GEN_334 : valid_331_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1359 = io_cpu_fence_value & _T & _T_2 ? _GEN_335 : valid_332_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1360 = io_cpu_fence_value & _T & _T_2 ? _GEN_336 : valid_333_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1361 = io_cpu_fence_value & _T & _T_2 ? _GEN_337 : valid_334_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1362 = io_cpu_fence_value & _T & _T_2 ? _GEN_338 : valid_335_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1363 = io_cpu_fence_value & _T & _T_2 ? _GEN_339 : valid_336_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1364 = io_cpu_fence_value & _T & _T_2 ? _GEN_340 : valid_337_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1365 = io_cpu_fence_value & _T & _T_2 ? _GEN_341 : valid_338_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1366 = io_cpu_fence_value & _T & _T_2 ? _GEN_342 : valid_339_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1367 = io_cpu_fence_value & _T & _T_2 ? _GEN_343 : valid_340_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1368 = io_cpu_fence_value & _T & _T_2 ? _GEN_344 : valid_341_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1369 = io_cpu_fence_value & _T & _T_2 ? _GEN_345 : valid_342_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1370 = io_cpu_fence_value & _T & _T_2 ? _GEN_346 : valid_343_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1371 = io_cpu_fence_value & _T & _T_2 ? _GEN_347 : valid_344_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1372 = io_cpu_fence_value & _T & _T_2 ? _GEN_348 : valid_345_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1373 = io_cpu_fence_value & _T & _T_2 ? _GEN_349 : valid_346_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1374 = io_cpu_fence_value & _T & _T_2 ? _GEN_350 : valid_347_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1375 = io_cpu_fence_value & _T & _T_2 ? _GEN_351 : valid_348_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1376 = io_cpu_fence_value & _T & _T_2 ? _GEN_352 : valid_349_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1377 = io_cpu_fence_value & _T & _T_2 ? _GEN_353 : valid_350_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1378 = io_cpu_fence_value & _T & _T_2 ? _GEN_354 : valid_351_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1379 = io_cpu_fence_value & _T & _T_2 ? _GEN_355 : valid_352_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1380 = io_cpu_fence_value & _T & _T_2 ? _GEN_356 : valid_353_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1381 = io_cpu_fence_value & _T & _T_2 ? _GEN_357 : valid_354_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1382 = io_cpu_fence_value & _T & _T_2 ? _GEN_358 : valid_355_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1383 = io_cpu_fence_value & _T & _T_2 ? _GEN_359 : valid_356_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1384 = io_cpu_fence_value & _T & _T_2 ? _GEN_360 : valid_357_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1385 = io_cpu_fence_value & _T & _T_2 ? _GEN_361 : valid_358_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1386 = io_cpu_fence_value & _T & _T_2 ? _GEN_362 : valid_359_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1387 = io_cpu_fence_value & _T & _T_2 ? _GEN_363 : valid_360_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1388 = io_cpu_fence_value & _T & _T_2 ? _GEN_364 : valid_361_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1389 = io_cpu_fence_value & _T & _T_2 ? _GEN_365 : valid_362_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1390 = io_cpu_fence_value & _T & _T_2 ? _GEN_366 : valid_363_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1391 = io_cpu_fence_value & _T & _T_2 ? _GEN_367 : valid_364_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1392 = io_cpu_fence_value & _T & _T_2 ? _GEN_368 : valid_365_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1393 = io_cpu_fence_value & _T & _T_2 ? _GEN_369 : valid_366_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1394 = io_cpu_fence_value & _T & _T_2 ? _GEN_370 : valid_367_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1395 = io_cpu_fence_value & _T & _T_2 ? _GEN_371 : valid_368_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1396 = io_cpu_fence_value & _T & _T_2 ? _GEN_372 : valid_369_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1397 = io_cpu_fence_value & _T & _T_2 ? _GEN_373 : valid_370_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1398 = io_cpu_fence_value & _T & _T_2 ? _GEN_374 : valid_371_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1399 = io_cpu_fence_value & _T & _T_2 ? _GEN_375 : valid_372_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1400 = io_cpu_fence_value & _T & _T_2 ? _GEN_376 : valid_373_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1401 = io_cpu_fence_value & _T & _T_2 ? _GEN_377 : valid_374_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1402 = io_cpu_fence_value & _T & _T_2 ? _GEN_378 : valid_375_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1403 = io_cpu_fence_value & _T & _T_2 ? _GEN_379 : valid_376_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1404 = io_cpu_fence_value & _T & _T_2 ? _GEN_380 : valid_377_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1405 = io_cpu_fence_value & _T & _T_2 ? _GEN_381 : valid_378_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1406 = io_cpu_fence_value & _T & _T_2 ? _GEN_382 : valid_379_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1407 = io_cpu_fence_value & _T & _T_2 ? _GEN_383 : valid_380_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1408 = io_cpu_fence_value & _T & _T_2 ? _GEN_384 : valid_381_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1409 = io_cpu_fence_value & _T & _T_2 ? _GEN_385 : valid_382_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1410 = io_cpu_fence_value & _T & _T_2 ? _GEN_386 : valid_383_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1411 = io_cpu_fence_value & _T & _T_2 ? _GEN_387 : valid_384_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1412 = io_cpu_fence_value & _T & _T_2 ? _GEN_388 : valid_385_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1413 = io_cpu_fence_value & _T & _T_2 ? _GEN_389 : valid_386_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1414 = io_cpu_fence_value & _T & _T_2 ? _GEN_390 : valid_387_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1415 = io_cpu_fence_value & _T & _T_2 ? _GEN_391 : valid_388_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1416 = io_cpu_fence_value & _T & _T_2 ? _GEN_392 : valid_389_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1417 = io_cpu_fence_value & _T & _T_2 ? _GEN_393 : valid_390_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1418 = io_cpu_fence_value & _T & _T_2 ? _GEN_394 : valid_391_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1419 = io_cpu_fence_value & _T & _T_2 ? _GEN_395 : valid_392_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1420 = io_cpu_fence_value & _T & _T_2 ? _GEN_396 : valid_393_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1421 = io_cpu_fence_value & _T & _T_2 ? _GEN_397 : valid_394_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1422 = io_cpu_fence_value & _T & _T_2 ? _GEN_398 : valid_395_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1423 = io_cpu_fence_value & _T & _T_2 ? _GEN_399 : valid_396_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1424 = io_cpu_fence_value & _T & _T_2 ? _GEN_400 : valid_397_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1425 = io_cpu_fence_value & _T & _T_2 ? _GEN_401 : valid_398_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1426 = io_cpu_fence_value & _T & _T_2 ? _GEN_402 : valid_399_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1427 = io_cpu_fence_value & _T & _T_2 ? _GEN_403 : valid_400_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1428 = io_cpu_fence_value & _T & _T_2 ? _GEN_404 : valid_401_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1429 = io_cpu_fence_value & _T & _T_2 ? _GEN_405 : valid_402_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1430 = io_cpu_fence_value & _T & _T_2 ? _GEN_406 : valid_403_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1431 = io_cpu_fence_value & _T & _T_2 ? _GEN_407 : valid_404_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1432 = io_cpu_fence_value & _T & _T_2 ? _GEN_408 : valid_405_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1433 = io_cpu_fence_value & _T & _T_2 ? _GEN_409 : valid_406_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1434 = io_cpu_fence_value & _T & _T_2 ? _GEN_410 : valid_407_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1435 = io_cpu_fence_value & _T & _T_2 ? _GEN_411 : valid_408_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1436 = io_cpu_fence_value & _T & _T_2 ? _GEN_412 : valid_409_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1437 = io_cpu_fence_value & _T & _T_2 ? _GEN_413 : valid_410_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1438 = io_cpu_fence_value & _T & _T_2 ? _GEN_414 : valid_411_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1439 = io_cpu_fence_value & _T & _T_2 ? _GEN_415 : valid_412_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1440 = io_cpu_fence_value & _T & _T_2 ? _GEN_416 : valid_413_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1441 = io_cpu_fence_value & _T & _T_2 ? _GEN_417 : valid_414_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1442 = io_cpu_fence_value & _T & _T_2 ? _GEN_418 : valid_415_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1443 = io_cpu_fence_value & _T & _T_2 ? _GEN_419 : valid_416_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1444 = io_cpu_fence_value & _T & _T_2 ? _GEN_420 : valid_417_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1445 = io_cpu_fence_value & _T & _T_2 ? _GEN_421 : valid_418_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1446 = io_cpu_fence_value & _T & _T_2 ? _GEN_422 : valid_419_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1447 = io_cpu_fence_value & _T & _T_2 ? _GEN_423 : valid_420_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1448 = io_cpu_fence_value & _T & _T_2 ? _GEN_424 : valid_421_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1449 = io_cpu_fence_value & _T & _T_2 ? _GEN_425 : valid_422_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1450 = io_cpu_fence_value & _T & _T_2 ? _GEN_426 : valid_423_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1451 = io_cpu_fence_value & _T & _T_2 ? _GEN_427 : valid_424_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1452 = io_cpu_fence_value & _T & _T_2 ? _GEN_428 : valid_425_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1453 = io_cpu_fence_value & _T & _T_2 ? _GEN_429 : valid_426_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1454 = io_cpu_fence_value & _T & _T_2 ? _GEN_430 : valid_427_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1455 = io_cpu_fence_value & _T & _T_2 ? _GEN_431 : valid_428_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1456 = io_cpu_fence_value & _T & _T_2 ? _GEN_432 : valid_429_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1457 = io_cpu_fence_value & _T & _T_2 ? _GEN_433 : valid_430_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1458 = io_cpu_fence_value & _T & _T_2 ? _GEN_434 : valid_431_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1459 = io_cpu_fence_value & _T & _T_2 ? _GEN_435 : valid_432_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1460 = io_cpu_fence_value & _T & _T_2 ? _GEN_436 : valid_433_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1461 = io_cpu_fence_value & _T & _T_2 ? _GEN_437 : valid_434_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1462 = io_cpu_fence_value & _T & _T_2 ? _GEN_438 : valid_435_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1463 = io_cpu_fence_value & _T & _T_2 ? _GEN_439 : valid_436_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1464 = io_cpu_fence_value & _T & _T_2 ? _GEN_440 : valid_437_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1465 = io_cpu_fence_value & _T & _T_2 ? _GEN_441 : valid_438_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1466 = io_cpu_fence_value & _T & _T_2 ? _GEN_442 : valid_439_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1467 = io_cpu_fence_value & _T & _T_2 ? _GEN_443 : valid_440_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1468 = io_cpu_fence_value & _T & _T_2 ? _GEN_444 : valid_441_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1469 = io_cpu_fence_value & _T & _T_2 ? _GEN_445 : valid_442_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1470 = io_cpu_fence_value & _T & _T_2 ? _GEN_446 : valid_443_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1471 = io_cpu_fence_value & _T & _T_2 ? _GEN_447 : valid_444_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1472 = io_cpu_fence_value & _T & _T_2 ? _GEN_448 : valid_445_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1473 = io_cpu_fence_value & _T & _T_2 ? _GEN_449 : valid_446_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1474 = io_cpu_fence_value & _T & _T_2 ? _GEN_450 : valid_447_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1475 = io_cpu_fence_value & _T & _T_2 ? _GEN_451 : valid_448_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1476 = io_cpu_fence_value & _T & _T_2 ? _GEN_452 : valid_449_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1477 = io_cpu_fence_value & _T & _T_2 ? _GEN_453 : valid_450_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1478 = io_cpu_fence_value & _T & _T_2 ? _GEN_454 : valid_451_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1479 = io_cpu_fence_value & _T & _T_2 ? _GEN_455 : valid_452_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1480 = io_cpu_fence_value & _T & _T_2 ? _GEN_456 : valid_453_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1481 = io_cpu_fence_value & _T & _T_2 ? _GEN_457 : valid_454_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1482 = io_cpu_fence_value & _T & _T_2 ? _GEN_458 : valid_455_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1483 = io_cpu_fence_value & _T & _T_2 ? _GEN_459 : valid_456_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1484 = io_cpu_fence_value & _T & _T_2 ? _GEN_460 : valid_457_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1485 = io_cpu_fence_value & _T & _T_2 ? _GEN_461 : valid_458_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1486 = io_cpu_fence_value & _T & _T_2 ? _GEN_462 : valid_459_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1487 = io_cpu_fence_value & _T & _T_2 ? _GEN_463 : valid_460_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1488 = io_cpu_fence_value & _T & _T_2 ? _GEN_464 : valid_461_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1489 = io_cpu_fence_value & _T & _T_2 ? _GEN_465 : valid_462_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1490 = io_cpu_fence_value & _T & _T_2 ? _GEN_466 : valid_463_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1491 = io_cpu_fence_value & _T & _T_2 ? _GEN_467 : valid_464_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1492 = io_cpu_fence_value & _T & _T_2 ? _GEN_468 : valid_465_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1493 = io_cpu_fence_value & _T & _T_2 ? _GEN_469 : valid_466_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1494 = io_cpu_fence_value & _T & _T_2 ? _GEN_470 : valid_467_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1495 = io_cpu_fence_value & _T & _T_2 ? _GEN_471 : valid_468_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1496 = io_cpu_fence_value & _T & _T_2 ? _GEN_472 : valid_469_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1497 = io_cpu_fence_value & _T & _T_2 ? _GEN_473 : valid_470_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1498 = io_cpu_fence_value & _T & _T_2 ? _GEN_474 : valid_471_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1499 = io_cpu_fence_value & _T & _T_2 ? _GEN_475 : valid_472_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1500 = io_cpu_fence_value & _T & _T_2 ? _GEN_476 : valid_473_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1501 = io_cpu_fence_value & _T & _T_2 ? _GEN_477 : valid_474_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1502 = io_cpu_fence_value & _T & _T_2 ? _GEN_478 : valid_475_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1503 = io_cpu_fence_value & _T & _T_2 ? _GEN_479 : valid_476_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1504 = io_cpu_fence_value & _T & _T_2 ? _GEN_480 : valid_477_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1505 = io_cpu_fence_value & _T & _T_2 ? _GEN_481 : valid_478_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1506 = io_cpu_fence_value & _T & _T_2 ? _GEN_482 : valid_479_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1507 = io_cpu_fence_value & _T & _T_2 ? _GEN_483 : valid_480_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1508 = io_cpu_fence_value & _T & _T_2 ? _GEN_484 : valid_481_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1509 = io_cpu_fence_value & _T & _T_2 ? _GEN_485 : valid_482_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1510 = io_cpu_fence_value & _T & _T_2 ? _GEN_486 : valid_483_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1511 = io_cpu_fence_value & _T & _T_2 ? _GEN_487 : valid_484_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1512 = io_cpu_fence_value & _T & _T_2 ? _GEN_488 : valid_485_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1513 = io_cpu_fence_value & _T & _T_2 ? _GEN_489 : valid_486_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1514 = io_cpu_fence_value & _T & _T_2 ? _GEN_490 : valid_487_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1515 = io_cpu_fence_value & _T & _T_2 ? _GEN_491 : valid_488_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1516 = io_cpu_fence_value & _T & _T_2 ? _GEN_492 : valid_489_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1517 = io_cpu_fence_value & _T & _T_2 ? _GEN_493 : valid_490_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1518 = io_cpu_fence_value & _T & _T_2 ? _GEN_494 : valid_491_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1519 = io_cpu_fence_value & _T & _T_2 ? _GEN_495 : valid_492_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1520 = io_cpu_fence_value & _T & _T_2 ? _GEN_496 : valid_493_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1521 = io_cpu_fence_value & _T & _T_2 ? _GEN_497 : valid_494_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1522 = io_cpu_fence_value & _T & _T_2 ? _GEN_498 : valid_495_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1523 = io_cpu_fence_value & _T & _T_2 ? _GEN_499 : valid_496_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1524 = io_cpu_fence_value & _T & _T_2 ? _GEN_500 : valid_497_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1525 = io_cpu_fence_value & _T & _T_2 ? _GEN_501 : valid_498_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1526 = io_cpu_fence_value & _T & _T_2 ? _GEN_502 : valid_499_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1527 = io_cpu_fence_value & _T & _T_2 ? _GEN_503 : valid_500_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1528 = io_cpu_fence_value & _T & _T_2 ? _GEN_504 : valid_501_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1529 = io_cpu_fence_value & _T & _T_2 ? _GEN_505 : valid_502_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1530 = io_cpu_fence_value & _T & _T_2 ? _GEN_506 : valid_503_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1531 = io_cpu_fence_value & _T & _T_2 ? _GEN_507 : valid_504_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1532 = io_cpu_fence_value & _T & _T_2 ? _GEN_508 : valid_505_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1533 = io_cpu_fence_value & _T & _T_2 ? _GEN_509 : valid_506_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1534 = io_cpu_fence_value & _T & _T_2 ? _GEN_510 : valid_507_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1535 = io_cpu_fence_value & _T & _T_2 ? _GEN_511 : valid_508_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1536 = io_cpu_fence_value & _T & _T_2 ? _GEN_512 : valid_509_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1537 = io_cpu_fence_value & _T & _T_2 ? _GEN_513 : valid_510_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1538 = io_cpu_fence_value & _T & _T_2 ? _GEN_514 : valid_511_0; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1539 = io_cpu_fence_value & _T & _T_2 ? _GEN_515 : valid_0_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1540 = io_cpu_fence_value & _T & _T_2 ? _GEN_516 : valid_1_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1541 = io_cpu_fence_value & _T & _T_2 ? _GEN_517 : valid_2_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1542 = io_cpu_fence_value & _T & _T_2 ? _GEN_518 : valid_3_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1543 = io_cpu_fence_value & _T & _T_2 ? _GEN_519 : valid_4_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1544 = io_cpu_fence_value & _T & _T_2 ? _GEN_520 : valid_5_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1545 = io_cpu_fence_value & _T & _T_2 ? _GEN_521 : valid_6_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1546 = io_cpu_fence_value & _T & _T_2 ? _GEN_522 : valid_7_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1547 = io_cpu_fence_value & _T & _T_2 ? _GEN_523 : valid_8_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1548 = io_cpu_fence_value & _T & _T_2 ? _GEN_524 : valid_9_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1549 = io_cpu_fence_value & _T & _T_2 ? _GEN_525 : valid_10_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1550 = io_cpu_fence_value & _T & _T_2 ? _GEN_526 : valid_11_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1551 = io_cpu_fence_value & _T & _T_2 ? _GEN_527 : valid_12_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1552 = io_cpu_fence_value & _T & _T_2 ? _GEN_528 : valid_13_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1553 = io_cpu_fence_value & _T & _T_2 ? _GEN_529 : valid_14_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1554 = io_cpu_fence_value & _T & _T_2 ? _GEN_530 : valid_15_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1555 = io_cpu_fence_value & _T & _T_2 ? _GEN_531 : valid_16_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1556 = io_cpu_fence_value & _T & _T_2 ? _GEN_532 : valid_17_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1557 = io_cpu_fence_value & _T & _T_2 ? _GEN_533 : valid_18_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1558 = io_cpu_fence_value & _T & _T_2 ? _GEN_534 : valid_19_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1559 = io_cpu_fence_value & _T & _T_2 ? _GEN_535 : valid_20_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1560 = io_cpu_fence_value & _T & _T_2 ? _GEN_536 : valid_21_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1561 = io_cpu_fence_value & _T & _T_2 ? _GEN_537 : valid_22_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1562 = io_cpu_fence_value & _T & _T_2 ? _GEN_538 : valid_23_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1563 = io_cpu_fence_value & _T & _T_2 ? _GEN_539 : valid_24_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1564 = io_cpu_fence_value & _T & _T_2 ? _GEN_540 : valid_25_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1565 = io_cpu_fence_value & _T & _T_2 ? _GEN_541 : valid_26_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1566 = io_cpu_fence_value & _T & _T_2 ? _GEN_542 : valid_27_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1567 = io_cpu_fence_value & _T & _T_2 ? _GEN_543 : valid_28_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1568 = io_cpu_fence_value & _T & _T_2 ? _GEN_544 : valid_29_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1569 = io_cpu_fence_value & _T & _T_2 ? _GEN_545 : valid_30_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1570 = io_cpu_fence_value & _T & _T_2 ? _GEN_546 : valid_31_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1571 = io_cpu_fence_value & _T & _T_2 ? _GEN_547 : valid_32_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1572 = io_cpu_fence_value & _T & _T_2 ? _GEN_548 : valid_33_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1573 = io_cpu_fence_value & _T & _T_2 ? _GEN_549 : valid_34_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1574 = io_cpu_fence_value & _T & _T_2 ? _GEN_550 : valid_35_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1575 = io_cpu_fence_value & _T & _T_2 ? _GEN_551 : valid_36_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1576 = io_cpu_fence_value & _T & _T_2 ? _GEN_552 : valid_37_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1577 = io_cpu_fence_value & _T & _T_2 ? _GEN_553 : valid_38_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1578 = io_cpu_fence_value & _T & _T_2 ? _GEN_554 : valid_39_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1579 = io_cpu_fence_value & _T & _T_2 ? _GEN_555 : valid_40_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1580 = io_cpu_fence_value & _T & _T_2 ? _GEN_556 : valid_41_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1581 = io_cpu_fence_value & _T & _T_2 ? _GEN_557 : valid_42_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1582 = io_cpu_fence_value & _T & _T_2 ? _GEN_558 : valid_43_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1583 = io_cpu_fence_value & _T & _T_2 ? _GEN_559 : valid_44_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1584 = io_cpu_fence_value & _T & _T_2 ? _GEN_560 : valid_45_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1585 = io_cpu_fence_value & _T & _T_2 ? _GEN_561 : valid_46_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1586 = io_cpu_fence_value & _T & _T_2 ? _GEN_562 : valid_47_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1587 = io_cpu_fence_value & _T & _T_2 ? _GEN_563 : valid_48_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1588 = io_cpu_fence_value & _T & _T_2 ? _GEN_564 : valid_49_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1589 = io_cpu_fence_value & _T & _T_2 ? _GEN_565 : valid_50_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1590 = io_cpu_fence_value & _T & _T_2 ? _GEN_566 : valid_51_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1591 = io_cpu_fence_value & _T & _T_2 ? _GEN_567 : valid_52_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1592 = io_cpu_fence_value & _T & _T_2 ? _GEN_568 : valid_53_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1593 = io_cpu_fence_value & _T & _T_2 ? _GEN_569 : valid_54_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1594 = io_cpu_fence_value & _T & _T_2 ? _GEN_570 : valid_55_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1595 = io_cpu_fence_value & _T & _T_2 ? _GEN_571 : valid_56_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1596 = io_cpu_fence_value & _T & _T_2 ? _GEN_572 : valid_57_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1597 = io_cpu_fence_value & _T & _T_2 ? _GEN_573 : valid_58_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1598 = io_cpu_fence_value & _T & _T_2 ? _GEN_574 : valid_59_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1599 = io_cpu_fence_value & _T & _T_2 ? _GEN_575 : valid_60_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1600 = io_cpu_fence_value & _T & _T_2 ? _GEN_576 : valid_61_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1601 = io_cpu_fence_value & _T & _T_2 ? _GEN_577 : valid_62_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1602 = io_cpu_fence_value & _T & _T_2 ? _GEN_578 : valid_63_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1603 = io_cpu_fence_value & _T & _T_2 ? _GEN_579 : valid_64_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1604 = io_cpu_fence_value & _T & _T_2 ? _GEN_580 : valid_65_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1605 = io_cpu_fence_value & _T & _T_2 ? _GEN_581 : valid_66_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1606 = io_cpu_fence_value & _T & _T_2 ? _GEN_582 : valid_67_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1607 = io_cpu_fence_value & _T & _T_2 ? _GEN_583 : valid_68_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1608 = io_cpu_fence_value & _T & _T_2 ? _GEN_584 : valid_69_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1609 = io_cpu_fence_value & _T & _T_2 ? _GEN_585 : valid_70_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1610 = io_cpu_fence_value & _T & _T_2 ? _GEN_586 : valid_71_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1611 = io_cpu_fence_value & _T & _T_2 ? _GEN_587 : valid_72_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1612 = io_cpu_fence_value & _T & _T_2 ? _GEN_588 : valid_73_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1613 = io_cpu_fence_value & _T & _T_2 ? _GEN_589 : valid_74_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1614 = io_cpu_fence_value & _T & _T_2 ? _GEN_590 : valid_75_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1615 = io_cpu_fence_value & _T & _T_2 ? _GEN_591 : valid_76_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1616 = io_cpu_fence_value & _T & _T_2 ? _GEN_592 : valid_77_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1617 = io_cpu_fence_value & _T & _T_2 ? _GEN_593 : valid_78_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1618 = io_cpu_fence_value & _T & _T_2 ? _GEN_594 : valid_79_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1619 = io_cpu_fence_value & _T & _T_2 ? _GEN_595 : valid_80_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1620 = io_cpu_fence_value & _T & _T_2 ? _GEN_596 : valid_81_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1621 = io_cpu_fence_value & _T & _T_2 ? _GEN_597 : valid_82_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1622 = io_cpu_fence_value & _T & _T_2 ? _GEN_598 : valid_83_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1623 = io_cpu_fence_value & _T & _T_2 ? _GEN_599 : valid_84_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1624 = io_cpu_fence_value & _T & _T_2 ? _GEN_600 : valid_85_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1625 = io_cpu_fence_value & _T & _T_2 ? _GEN_601 : valid_86_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1626 = io_cpu_fence_value & _T & _T_2 ? _GEN_602 : valid_87_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1627 = io_cpu_fence_value & _T & _T_2 ? _GEN_603 : valid_88_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1628 = io_cpu_fence_value & _T & _T_2 ? _GEN_604 : valid_89_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1629 = io_cpu_fence_value & _T & _T_2 ? _GEN_605 : valid_90_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1630 = io_cpu_fence_value & _T & _T_2 ? _GEN_606 : valid_91_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1631 = io_cpu_fence_value & _T & _T_2 ? _GEN_607 : valid_92_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1632 = io_cpu_fence_value & _T & _T_2 ? _GEN_608 : valid_93_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1633 = io_cpu_fence_value & _T & _T_2 ? _GEN_609 : valid_94_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1634 = io_cpu_fence_value & _T & _T_2 ? _GEN_610 : valid_95_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1635 = io_cpu_fence_value & _T & _T_2 ? _GEN_611 : valid_96_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1636 = io_cpu_fence_value & _T & _T_2 ? _GEN_612 : valid_97_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1637 = io_cpu_fence_value & _T & _T_2 ? _GEN_613 : valid_98_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1638 = io_cpu_fence_value & _T & _T_2 ? _GEN_614 : valid_99_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1639 = io_cpu_fence_value & _T & _T_2 ? _GEN_615 : valid_100_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1640 = io_cpu_fence_value & _T & _T_2 ? _GEN_616 : valid_101_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1641 = io_cpu_fence_value & _T & _T_2 ? _GEN_617 : valid_102_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1642 = io_cpu_fence_value & _T & _T_2 ? _GEN_618 : valid_103_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1643 = io_cpu_fence_value & _T & _T_2 ? _GEN_619 : valid_104_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1644 = io_cpu_fence_value & _T & _T_2 ? _GEN_620 : valid_105_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1645 = io_cpu_fence_value & _T & _T_2 ? _GEN_621 : valid_106_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1646 = io_cpu_fence_value & _T & _T_2 ? _GEN_622 : valid_107_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1647 = io_cpu_fence_value & _T & _T_2 ? _GEN_623 : valid_108_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1648 = io_cpu_fence_value & _T & _T_2 ? _GEN_624 : valid_109_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1649 = io_cpu_fence_value & _T & _T_2 ? _GEN_625 : valid_110_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1650 = io_cpu_fence_value & _T & _T_2 ? _GEN_626 : valid_111_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1651 = io_cpu_fence_value & _T & _T_2 ? _GEN_627 : valid_112_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1652 = io_cpu_fence_value & _T & _T_2 ? _GEN_628 : valid_113_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1653 = io_cpu_fence_value & _T & _T_2 ? _GEN_629 : valid_114_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1654 = io_cpu_fence_value & _T & _T_2 ? _GEN_630 : valid_115_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1655 = io_cpu_fence_value & _T & _T_2 ? _GEN_631 : valid_116_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1656 = io_cpu_fence_value & _T & _T_2 ? _GEN_632 : valid_117_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1657 = io_cpu_fence_value & _T & _T_2 ? _GEN_633 : valid_118_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1658 = io_cpu_fence_value & _T & _T_2 ? _GEN_634 : valid_119_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1659 = io_cpu_fence_value & _T & _T_2 ? _GEN_635 : valid_120_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1660 = io_cpu_fence_value & _T & _T_2 ? _GEN_636 : valid_121_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1661 = io_cpu_fence_value & _T & _T_2 ? _GEN_637 : valid_122_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1662 = io_cpu_fence_value & _T & _T_2 ? _GEN_638 : valid_123_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1663 = io_cpu_fence_value & _T & _T_2 ? _GEN_639 : valid_124_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1664 = io_cpu_fence_value & _T & _T_2 ? _GEN_640 : valid_125_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1665 = io_cpu_fence_value & _T & _T_2 ? _GEN_641 : valid_126_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1666 = io_cpu_fence_value & _T & _T_2 ? _GEN_642 : valid_127_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1667 = io_cpu_fence_value & _T & _T_2 ? _GEN_643 : valid_128_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1668 = io_cpu_fence_value & _T & _T_2 ? _GEN_644 : valid_129_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1669 = io_cpu_fence_value & _T & _T_2 ? _GEN_645 : valid_130_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1670 = io_cpu_fence_value & _T & _T_2 ? _GEN_646 : valid_131_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1671 = io_cpu_fence_value & _T & _T_2 ? _GEN_647 : valid_132_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1672 = io_cpu_fence_value & _T & _T_2 ? _GEN_648 : valid_133_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1673 = io_cpu_fence_value & _T & _T_2 ? _GEN_649 : valid_134_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1674 = io_cpu_fence_value & _T & _T_2 ? _GEN_650 : valid_135_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1675 = io_cpu_fence_value & _T & _T_2 ? _GEN_651 : valid_136_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1676 = io_cpu_fence_value & _T & _T_2 ? _GEN_652 : valid_137_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1677 = io_cpu_fence_value & _T & _T_2 ? _GEN_653 : valid_138_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1678 = io_cpu_fence_value & _T & _T_2 ? _GEN_654 : valid_139_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1679 = io_cpu_fence_value & _T & _T_2 ? _GEN_655 : valid_140_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1680 = io_cpu_fence_value & _T & _T_2 ? _GEN_656 : valid_141_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1681 = io_cpu_fence_value & _T & _T_2 ? _GEN_657 : valid_142_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1682 = io_cpu_fence_value & _T & _T_2 ? _GEN_658 : valid_143_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1683 = io_cpu_fence_value & _T & _T_2 ? _GEN_659 : valid_144_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1684 = io_cpu_fence_value & _T & _T_2 ? _GEN_660 : valid_145_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1685 = io_cpu_fence_value & _T & _T_2 ? _GEN_661 : valid_146_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1686 = io_cpu_fence_value & _T & _T_2 ? _GEN_662 : valid_147_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1687 = io_cpu_fence_value & _T & _T_2 ? _GEN_663 : valid_148_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1688 = io_cpu_fence_value & _T & _T_2 ? _GEN_664 : valid_149_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1689 = io_cpu_fence_value & _T & _T_2 ? _GEN_665 : valid_150_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1690 = io_cpu_fence_value & _T & _T_2 ? _GEN_666 : valid_151_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1691 = io_cpu_fence_value & _T & _T_2 ? _GEN_667 : valid_152_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1692 = io_cpu_fence_value & _T & _T_2 ? _GEN_668 : valid_153_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1693 = io_cpu_fence_value & _T & _T_2 ? _GEN_669 : valid_154_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1694 = io_cpu_fence_value & _T & _T_2 ? _GEN_670 : valid_155_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1695 = io_cpu_fence_value & _T & _T_2 ? _GEN_671 : valid_156_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1696 = io_cpu_fence_value & _T & _T_2 ? _GEN_672 : valid_157_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1697 = io_cpu_fence_value & _T & _T_2 ? _GEN_673 : valid_158_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1698 = io_cpu_fence_value & _T & _T_2 ? _GEN_674 : valid_159_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1699 = io_cpu_fence_value & _T & _T_2 ? _GEN_675 : valid_160_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1700 = io_cpu_fence_value & _T & _T_2 ? _GEN_676 : valid_161_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1701 = io_cpu_fence_value & _T & _T_2 ? _GEN_677 : valid_162_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1702 = io_cpu_fence_value & _T & _T_2 ? _GEN_678 : valid_163_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1703 = io_cpu_fence_value & _T & _T_2 ? _GEN_679 : valid_164_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1704 = io_cpu_fence_value & _T & _T_2 ? _GEN_680 : valid_165_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1705 = io_cpu_fence_value & _T & _T_2 ? _GEN_681 : valid_166_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1706 = io_cpu_fence_value & _T & _T_2 ? _GEN_682 : valid_167_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1707 = io_cpu_fence_value & _T & _T_2 ? _GEN_683 : valid_168_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1708 = io_cpu_fence_value & _T & _T_2 ? _GEN_684 : valid_169_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1709 = io_cpu_fence_value & _T & _T_2 ? _GEN_685 : valid_170_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1710 = io_cpu_fence_value & _T & _T_2 ? _GEN_686 : valid_171_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1711 = io_cpu_fence_value & _T & _T_2 ? _GEN_687 : valid_172_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1712 = io_cpu_fence_value & _T & _T_2 ? _GEN_688 : valid_173_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1713 = io_cpu_fence_value & _T & _T_2 ? _GEN_689 : valid_174_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1714 = io_cpu_fence_value & _T & _T_2 ? _GEN_690 : valid_175_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1715 = io_cpu_fence_value & _T & _T_2 ? _GEN_691 : valid_176_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1716 = io_cpu_fence_value & _T & _T_2 ? _GEN_692 : valid_177_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1717 = io_cpu_fence_value & _T & _T_2 ? _GEN_693 : valid_178_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1718 = io_cpu_fence_value & _T & _T_2 ? _GEN_694 : valid_179_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1719 = io_cpu_fence_value & _T & _T_2 ? _GEN_695 : valid_180_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1720 = io_cpu_fence_value & _T & _T_2 ? _GEN_696 : valid_181_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1721 = io_cpu_fence_value & _T & _T_2 ? _GEN_697 : valid_182_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1722 = io_cpu_fence_value & _T & _T_2 ? _GEN_698 : valid_183_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1723 = io_cpu_fence_value & _T & _T_2 ? _GEN_699 : valid_184_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1724 = io_cpu_fence_value & _T & _T_2 ? _GEN_700 : valid_185_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1725 = io_cpu_fence_value & _T & _T_2 ? _GEN_701 : valid_186_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1726 = io_cpu_fence_value & _T & _T_2 ? _GEN_702 : valid_187_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1727 = io_cpu_fence_value & _T & _T_2 ? _GEN_703 : valid_188_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1728 = io_cpu_fence_value & _T & _T_2 ? _GEN_704 : valid_189_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1729 = io_cpu_fence_value & _T & _T_2 ? _GEN_705 : valid_190_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1730 = io_cpu_fence_value & _T & _T_2 ? _GEN_706 : valid_191_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1731 = io_cpu_fence_value & _T & _T_2 ? _GEN_707 : valid_192_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1732 = io_cpu_fence_value & _T & _T_2 ? _GEN_708 : valid_193_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1733 = io_cpu_fence_value & _T & _T_2 ? _GEN_709 : valid_194_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1734 = io_cpu_fence_value & _T & _T_2 ? _GEN_710 : valid_195_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1735 = io_cpu_fence_value & _T & _T_2 ? _GEN_711 : valid_196_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1736 = io_cpu_fence_value & _T & _T_2 ? _GEN_712 : valid_197_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1737 = io_cpu_fence_value & _T & _T_2 ? _GEN_713 : valid_198_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1738 = io_cpu_fence_value & _T & _T_2 ? _GEN_714 : valid_199_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1739 = io_cpu_fence_value & _T & _T_2 ? _GEN_715 : valid_200_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1740 = io_cpu_fence_value & _T & _T_2 ? _GEN_716 : valid_201_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1741 = io_cpu_fence_value & _T & _T_2 ? _GEN_717 : valid_202_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1742 = io_cpu_fence_value & _T & _T_2 ? _GEN_718 : valid_203_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1743 = io_cpu_fence_value & _T & _T_2 ? _GEN_719 : valid_204_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1744 = io_cpu_fence_value & _T & _T_2 ? _GEN_720 : valid_205_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1745 = io_cpu_fence_value & _T & _T_2 ? _GEN_721 : valid_206_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1746 = io_cpu_fence_value & _T & _T_2 ? _GEN_722 : valid_207_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1747 = io_cpu_fence_value & _T & _T_2 ? _GEN_723 : valid_208_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1748 = io_cpu_fence_value & _T & _T_2 ? _GEN_724 : valid_209_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1749 = io_cpu_fence_value & _T & _T_2 ? _GEN_725 : valid_210_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1750 = io_cpu_fence_value & _T & _T_2 ? _GEN_726 : valid_211_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1751 = io_cpu_fence_value & _T & _T_2 ? _GEN_727 : valid_212_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1752 = io_cpu_fence_value & _T & _T_2 ? _GEN_728 : valid_213_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1753 = io_cpu_fence_value & _T & _T_2 ? _GEN_729 : valid_214_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1754 = io_cpu_fence_value & _T & _T_2 ? _GEN_730 : valid_215_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1755 = io_cpu_fence_value & _T & _T_2 ? _GEN_731 : valid_216_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1756 = io_cpu_fence_value & _T & _T_2 ? _GEN_732 : valid_217_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1757 = io_cpu_fence_value & _T & _T_2 ? _GEN_733 : valid_218_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1758 = io_cpu_fence_value & _T & _T_2 ? _GEN_734 : valid_219_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1759 = io_cpu_fence_value & _T & _T_2 ? _GEN_735 : valid_220_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1760 = io_cpu_fence_value & _T & _T_2 ? _GEN_736 : valid_221_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1761 = io_cpu_fence_value & _T & _T_2 ? _GEN_737 : valid_222_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1762 = io_cpu_fence_value & _T & _T_2 ? _GEN_738 : valid_223_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1763 = io_cpu_fence_value & _T & _T_2 ? _GEN_739 : valid_224_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1764 = io_cpu_fence_value & _T & _T_2 ? _GEN_740 : valid_225_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1765 = io_cpu_fence_value & _T & _T_2 ? _GEN_741 : valid_226_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1766 = io_cpu_fence_value & _T & _T_2 ? _GEN_742 : valid_227_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1767 = io_cpu_fence_value & _T & _T_2 ? _GEN_743 : valid_228_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1768 = io_cpu_fence_value & _T & _T_2 ? _GEN_744 : valid_229_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1769 = io_cpu_fence_value & _T & _T_2 ? _GEN_745 : valid_230_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1770 = io_cpu_fence_value & _T & _T_2 ? _GEN_746 : valid_231_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1771 = io_cpu_fence_value & _T & _T_2 ? _GEN_747 : valid_232_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1772 = io_cpu_fence_value & _T & _T_2 ? _GEN_748 : valid_233_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1773 = io_cpu_fence_value & _T & _T_2 ? _GEN_749 : valid_234_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1774 = io_cpu_fence_value & _T & _T_2 ? _GEN_750 : valid_235_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1775 = io_cpu_fence_value & _T & _T_2 ? _GEN_751 : valid_236_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1776 = io_cpu_fence_value & _T & _T_2 ? _GEN_752 : valid_237_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1777 = io_cpu_fence_value & _T & _T_2 ? _GEN_753 : valid_238_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1778 = io_cpu_fence_value & _T & _T_2 ? _GEN_754 : valid_239_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1779 = io_cpu_fence_value & _T & _T_2 ? _GEN_755 : valid_240_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1780 = io_cpu_fence_value & _T & _T_2 ? _GEN_756 : valid_241_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1781 = io_cpu_fence_value & _T & _T_2 ? _GEN_757 : valid_242_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1782 = io_cpu_fence_value & _T & _T_2 ? _GEN_758 : valid_243_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1783 = io_cpu_fence_value & _T & _T_2 ? _GEN_759 : valid_244_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1784 = io_cpu_fence_value & _T & _T_2 ? _GEN_760 : valid_245_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1785 = io_cpu_fence_value & _T & _T_2 ? _GEN_761 : valid_246_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1786 = io_cpu_fence_value & _T & _T_2 ? _GEN_762 : valid_247_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1787 = io_cpu_fence_value & _T & _T_2 ? _GEN_763 : valid_248_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1788 = io_cpu_fence_value & _T & _T_2 ? _GEN_764 : valid_249_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1789 = io_cpu_fence_value & _T & _T_2 ? _GEN_765 : valid_250_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1790 = io_cpu_fence_value & _T & _T_2 ? _GEN_766 : valid_251_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1791 = io_cpu_fence_value & _T & _T_2 ? _GEN_767 : valid_252_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1792 = io_cpu_fence_value & _T & _T_2 ? _GEN_768 : valid_253_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1793 = io_cpu_fence_value & _T & _T_2 ? _GEN_769 : valid_254_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1794 = io_cpu_fence_value & _T & _T_2 ? _GEN_770 : valid_255_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1795 = io_cpu_fence_value & _T & _T_2 ? _GEN_771 : valid_256_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1796 = io_cpu_fence_value & _T & _T_2 ? _GEN_772 : valid_257_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1797 = io_cpu_fence_value & _T & _T_2 ? _GEN_773 : valid_258_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1798 = io_cpu_fence_value & _T & _T_2 ? _GEN_774 : valid_259_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1799 = io_cpu_fence_value & _T & _T_2 ? _GEN_775 : valid_260_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1800 = io_cpu_fence_value & _T & _T_2 ? _GEN_776 : valid_261_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1801 = io_cpu_fence_value & _T & _T_2 ? _GEN_777 : valid_262_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1802 = io_cpu_fence_value & _T & _T_2 ? _GEN_778 : valid_263_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1803 = io_cpu_fence_value & _T & _T_2 ? _GEN_779 : valid_264_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1804 = io_cpu_fence_value & _T & _T_2 ? _GEN_780 : valid_265_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1805 = io_cpu_fence_value & _T & _T_2 ? _GEN_781 : valid_266_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1806 = io_cpu_fence_value & _T & _T_2 ? _GEN_782 : valid_267_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1807 = io_cpu_fence_value & _T & _T_2 ? _GEN_783 : valid_268_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1808 = io_cpu_fence_value & _T & _T_2 ? _GEN_784 : valid_269_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1809 = io_cpu_fence_value & _T & _T_2 ? _GEN_785 : valid_270_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1810 = io_cpu_fence_value & _T & _T_2 ? _GEN_786 : valid_271_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1811 = io_cpu_fence_value & _T & _T_2 ? _GEN_787 : valid_272_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1812 = io_cpu_fence_value & _T & _T_2 ? _GEN_788 : valid_273_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1813 = io_cpu_fence_value & _T & _T_2 ? _GEN_789 : valid_274_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1814 = io_cpu_fence_value & _T & _T_2 ? _GEN_790 : valid_275_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1815 = io_cpu_fence_value & _T & _T_2 ? _GEN_791 : valid_276_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1816 = io_cpu_fence_value & _T & _T_2 ? _GEN_792 : valid_277_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1817 = io_cpu_fence_value & _T & _T_2 ? _GEN_793 : valid_278_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1818 = io_cpu_fence_value & _T & _T_2 ? _GEN_794 : valid_279_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1819 = io_cpu_fence_value & _T & _T_2 ? _GEN_795 : valid_280_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1820 = io_cpu_fence_value & _T & _T_2 ? _GEN_796 : valid_281_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1821 = io_cpu_fence_value & _T & _T_2 ? _GEN_797 : valid_282_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1822 = io_cpu_fence_value & _T & _T_2 ? _GEN_798 : valid_283_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1823 = io_cpu_fence_value & _T & _T_2 ? _GEN_799 : valid_284_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1824 = io_cpu_fence_value & _T & _T_2 ? _GEN_800 : valid_285_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1825 = io_cpu_fence_value & _T & _T_2 ? _GEN_801 : valid_286_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1826 = io_cpu_fence_value & _T & _T_2 ? _GEN_802 : valid_287_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1827 = io_cpu_fence_value & _T & _T_2 ? _GEN_803 : valid_288_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1828 = io_cpu_fence_value & _T & _T_2 ? _GEN_804 : valid_289_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1829 = io_cpu_fence_value & _T & _T_2 ? _GEN_805 : valid_290_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1830 = io_cpu_fence_value & _T & _T_2 ? _GEN_806 : valid_291_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1831 = io_cpu_fence_value & _T & _T_2 ? _GEN_807 : valid_292_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1832 = io_cpu_fence_value & _T & _T_2 ? _GEN_808 : valid_293_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1833 = io_cpu_fence_value & _T & _T_2 ? _GEN_809 : valid_294_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1834 = io_cpu_fence_value & _T & _T_2 ? _GEN_810 : valid_295_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1835 = io_cpu_fence_value & _T & _T_2 ? _GEN_811 : valid_296_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1836 = io_cpu_fence_value & _T & _T_2 ? _GEN_812 : valid_297_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1837 = io_cpu_fence_value & _T & _T_2 ? _GEN_813 : valid_298_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1838 = io_cpu_fence_value & _T & _T_2 ? _GEN_814 : valid_299_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1839 = io_cpu_fence_value & _T & _T_2 ? _GEN_815 : valid_300_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1840 = io_cpu_fence_value & _T & _T_2 ? _GEN_816 : valid_301_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1841 = io_cpu_fence_value & _T & _T_2 ? _GEN_817 : valid_302_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1842 = io_cpu_fence_value & _T & _T_2 ? _GEN_818 : valid_303_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1843 = io_cpu_fence_value & _T & _T_2 ? _GEN_819 : valid_304_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1844 = io_cpu_fence_value & _T & _T_2 ? _GEN_820 : valid_305_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1845 = io_cpu_fence_value & _T & _T_2 ? _GEN_821 : valid_306_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1846 = io_cpu_fence_value & _T & _T_2 ? _GEN_822 : valid_307_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1847 = io_cpu_fence_value & _T & _T_2 ? _GEN_823 : valid_308_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1848 = io_cpu_fence_value & _T & _T_2 ? _GEN_824 : valid_309_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1849 = io_cpu_fence_value & _T & _T_2 ? _GEN_825 : valid_310_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1850 = io_cpu_fence_value & _T & _T_2 ? _GEN_826 : valid_311_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1851 = io_cpu_fence_value & _T & _T_2 ? _GEN_827 : valid_312_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1852 = io_cpu_fence_value & _T & _T_2 ? _GEN_828 : valid_313_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1853 = io_cpu_fence_value & _T & _T_2 ? _GEN_829 : valid_314_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1854 = io_cpu_fence_value & _T & _T_2 ? _GEN_830 : valid_315_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1855 = io_cpu_fence_value & _T & _T_2 ? _GEN_831 : valid_316_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1856 = io_cpu_fence_value & _T & _T_2 ? _GEN_832 : valid_317_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1857 = io_cpu_fence_value & _T & _T_2 ? _GEN_833 : valid_318_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1858 = io_cpu_fence_value & _T & _T_2 ? _GEN_834 : valid_319_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1859 = io_cpu_fence_value & _T & _T_2 ? _GEN_835 : valid_320_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1860 = io_cpu_fence_value & _T & _T_2 ? _GEN_836 : valid_321_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1861 = io_cpu_fence_value & _T & _T_2 ? _GEN_837 : valid_322_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1862 = io_cpu_fence_value & _T & _T_2 ? _GEN_838 : valid_323_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1863 = io_cpu_fence_value & _T & _T_2 ? _GEN_839 : valid_324_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1864 = io_cpu_fence_value & _T & _T_2 ? _GEN_840 : valid_325_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1865 = io_cpu_fence_value & _T & _T_2 ? _GEN_841 : valid_326_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1866 = io_cpu_fence_value & _T & _T_2 ? _GEN_842 : valid_327_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1867 = io_cpu_fence_value & _T & _T_2 ? _GEN_843 : valid_328_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1868 = io_cpu_fence_value & _T & _T_2 ? _GEN_844 : valid_329_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1869 = io_cpu_fence_value & _T & _T_2 ? _GEN_845 : valid_330_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1870 = io_cpu_fence_value & _T & _T_2 ? _GEN_846 : valid_331_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1871 = io_cpu_fence_value & _T & _T_2 ? _GEN_847 : valid_332_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1872 = io_cpu_fence_value & _T & _T_2 ? _GEN_848 : valid_333_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1873 = io_cpu_fence_value & _T & _T_2 ? _GEN_849 : valid_334_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1874 = io_cpu_fence_value & _T & _T_2 ? _GEN_850 : valid_335_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1875 = io_cpu_fence_value & _T & _T_2 ? _GEN_851 : valid_336_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1876 = io_cpu_fence_value & _T & _T_2 ? _GEN_852 : valid_337_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1877 = io_cpu_fence_value & _T & _T_2 ? _GEN_853 : valid_338_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1878 = io_cpu_fence_value & _T & _T_2 ? _GEN_854 : valid_339_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1879 = io_cpu_fence_value & _T & _T_2 ? _GEN_855 : valid_340_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1880 = io_cpu_fence_value & _T & _T_2 ? _GEN_856 : valid_341_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1881 = io_cpu_fence_value & _T & _T_2 ? _GEN_857 : valid_342_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1882 = io_cpu_fence_value & _T & _T_2 ? _GEN_858 : valid_343_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1883 = io_cpu_fence_value & _T & _T_2 ? _GEN_859 : valid_344_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1884 = io_cpu_fence_value & _T & _T_2 ? _GEN_860 : valid_345_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1885 = io_cpu_fence_value & _T & _T_2 ? _GEN_861 : valid_346_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1886 = io_cpu_fence_value & _T & _T_2 ? _GEN_862 : valid_347_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1887 = io_cpu_fence_value & _T & _T_2 ? _GEN_863 : valid_348_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1888 = io_cpu_fence_value & _T & _T_2 ? _GEN_864 : valid_349_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1889 = io_cpu_fence_value & _T & _T_2 ? _GEN_865 : valid_350_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1890 = io_cpu_fence_value & _T & _T_2 ? _GEN_866 : valid_351_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1891 = io_cpu_fence_value & _T & _T_2 ? _GEN_867 : valid_352_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1892 = io_cpu_fence_value & _T & _T_2 ? _GEN_868 : valid_353_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1893 = io_cpu_fence_value & _T & _T_2 ? _GEN_869 : valid_354_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1894 = io_cpu_fence_value & _T & _T_2 ? _GEN_870 : valid_355_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1895 = io_cpu_fence_value & _T & _T_2 ? _GEN_871 : valid_356_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1896 = io_cpu_fence_value & _T & _T_2 ? _GEN_872 : valid_357_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1897 = io_cpu_fence_value & _T & _T_2 ? _GEN_873 : valid_358_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1898 = io_cpu_fence_value & _T & _T_2 ? _GEN_874 : valid_359_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1899 = io_cpu_fence_value & _T & _T_2 ? _GEN_875 : valid_360_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1900 = io_cpu_fence_value & _T & _T_2 ? _GEN_876 : valid_361_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1901 = io_cpu_fence_value & _T & _T_2 ? _GEN_877 : valid_362_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1902 = io_cpu_fence_value & _T & _T_2 ? _GEN_878 : valid_363_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1903 = io_cpu_fence_value & _T & _T_2 ? _GEN_879 : valid_364_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1904 = io_cpu_fence_value & _T & _T_2 ? _GEN_880 : valid_365_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1905 = io_cpu_fence_value & _T & _T_2 ? _GEN_881 : valid_366_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1906 = io_cpu_fence_value & _T & _T_2 ? _GEN_882 : valid_367_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1907 = io_cpu_fence_value & _T & _T_2 ? _GEN_883 : valid_368_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1908 = io_cpu_fence_value & _T & _T_2 ? _GEN_884 : valid_369_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1909 = io_cpu_fence_value & _T & _T_2 ? _GEN_885 : valid_370_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1910 = io_cpu_fence_value & _T & _T_2 ? _GEN_886 : valid_371_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1911 = io_cpu_fence_value & _T & _T_2 ? _GEN_887 : valid_372_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1912 = io_cpu_fence_value & _T & _T_2 ? _GEN_888 : valid_373_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1913 = io_cpu_fence_value & _T & _T_2 ? _GEN_889 : valid_374_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1914 = io_cpu_fence_value & _T & _T_2 ? _GEN_890 : valid_375_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1915 = io_cpu_fence_value & _T & _T_2 ? _GEN_891 : valid_376_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1916 = io_cpu_fence_value & _T & _T_2 ? _GEN_892 : valid_377_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1917 = io_cpu_fence_value & _T & _T_2 ? _GEN_893 : valid_378_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1918 = io_cpu_fence_value & _T & _T_2 ? _GEN_894 : valid_379_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1919 = io_cpu_fence_value & _T & _T_2 ? _GEN_895 : valid_380_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1920 = io_cpu_fence_value & _T & _T_2 ? _GEN_896 : valid_381_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1921 = io_cpu_fence_value & _T & _T_2 ? _GEN_897 : valid_382_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1922 = io_cpu_fence_value & _T & _T_2 ? _GEN_898 : valid_383_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1923 = io_cpu_fence_value & _T & _T_2 ? _GEN_899 : valid_384_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1924 = io_cpu_fence_value & _T & _T_2 ? _GEN_900 : valid_385_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1925 = io_cpu_fence_value & _T & _T_2 ? _GEN_901 : valid_386_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1926 = io_cpu_fence_value & _T & _T_2 ? _GEN_902 : valid_387_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1927 = io_cpu_fence_value & _T & _T_2 ? _GEN_903 : valid_388_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1928 = io_cpu_fence_value & _T & _T_2 ? _GEN_904 : valid_389_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1929 = io_cpu_fence_value & _T & _T_2 ? _GEN_905 : valid_390_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1930 = io_cpu_fence_value & _T & _T_2 ? _GEN_906 : valid_391_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1931 = io_cpu_fence_value & _T & _T_2 ? _GEN_907 : valid_392_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1932 = io_cpu_fence_value & _T & _T_2 ? _GEN_908 : valid_393_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1933 = io_cpu_fence_value & _T & _T_2 ? _GEN_909 : valid_394_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1934 = io_cpu_fence_value & _T & _T_2 ? _GEN_910 : valid_395_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1935 = io_cpu_fence_value & _T & _T_2 ? _GEN_911 : valid_396_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1936 = io_cpu_fence_value & _T & _T_2 ? _GEN_912 : valid_397_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1937 = io_cpu_fence_value & _T & _T_2 ? _GEN_913 : valid_398_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1938 = io_cpu_fence_value & _T & _T_2 ? _GEN_914 : valid_399_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1939 = io_cpu_fence_value & _T & _T_2 ? _GEN_915 : valid_400_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1940 = io_cpu_fence_value & _T & _T_2 ? _GEN_916 : valid_401_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1941 = io_cpu_fence_value & _T & _T_2 ? _GEN_917 : valid_402_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1942 = io_cpu_fence_value & _T & _T_2 ? _GEN_918 : valid_403_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1943 = io_cpu_fence_value & _T & _T_2 ? _GEN_919 : valid_404_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1944 = io_cpu_fence_value & _T & _T_2 ? _GEN_920 : valid_405_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1945 = io_cpu_fence_value & _T & _T_2 ? _GEN_921 : valid_406_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1946 = io_cpu_fence_value & _T & _T_2 ? _GEN_922 : valid_407_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1947 = io_cpu_fence_value & _T & _T_2 ? _GEN_923 : valid_408_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1948 = io_cpu_fence_value & _T & _T_2 ? _GEN_924 : valid_409_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1949 = io_cpu_fence_value & _T & _T_2 ? _GEN_925 : valid_410_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1950 = io_cpu_fence_value & _T & _T_2 ? _GEN_926 : valid_411_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1951 = io_cpu_fence_value & _T & _T_2 ? _GEN_927 : valid_412_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1952 = io_cpu_fence_value & _T & _T_2 ? _GEN_928 : valid_413_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1953 = io_cpu_fence_value & _T & _T_2 ? _GEN_929 : valid_414_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1954 = io_cpu_fence_value & _T & _T_2 ? _GEN_930 : valid_415_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1955 = io_cpu_fence_value & _T & _T_2 ? _GEN_931 : valid_416_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1956 = io_cpu_fence_value & _T & _T_2 ? _GEN_932 : valid_417_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1957 = io_cpu_fence_value & _T & _T_2 ? _GEN_933 : valid_418_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1958 = io_cpu_fence_value & _T & _T_2 ? _GEN_934 : valid_419_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1959 = io_cpu_fence_value & _T & _T_2 ? _GEN_935 : valid_420_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1960 = io_cpu_fence_value & _T & _T_2 ? _GEN_936 : valid_421_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1961 = io_cpu_fence_value & _T & _T_2 ? _GEN_937 : valid_422_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1962 = io_cpu_fence_value & _T & _T_2 ? _GEN_938 : valid_423_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1963 = io_cpu_fence_value & _T & _T_2 ? _GEN_939 : valid_424_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1964 = io_cpu_fence_value & _T & _T_2 ? _GEN_940 : valid_425_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1965 = io_cpu_fence_value & _T & _T_2 ? _GEN_941 : valid_426_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1966 = io_cpu_fence_value & _T & _T_2 ? _GEN_942 : valid_427_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1967 = io_cpu_fence_value & _T & _T_2 ? _GEN_943 : valid_428_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1968 = io_cpu_fence_value & _T & _T_2 ? _GEN_944 : valid_429_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1969 = io_cpu_fence_value & _T & _T_2 ? _GEN_945 : valid_430_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1970 = io_cpu_fence_value & _T & _T_2 ? _GEN_946 : valid_431_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1971 = io_cpu_fence_value & _T & _T_2 ? _GEN_947 : valid_432_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1972 = io_cpu_fence_value & _T & _T_2 ? _GEN_948 : valid_433_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1973 = io_cpu_fence_value & _T & _T_2 ? _GEN_949 : valid_434_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1974 = io_cpu_fence_value & _T & _T_2 ? _GEN_950 : valid_435_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1975 = io_cpu_fence_value & _T & _T_2 ? _GEN_951 : valid_436_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1976 = io_cpu_fence_value & _T & _T_2 ? _GEN_952 : valid_437_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1977 = io_cpu_fence_value & _T & _T_2 ? _GEN_953 : valid_438_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1978 = io_cpu_fence_value & _T & _T_2 ? _GEN_954 : valid_439_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1979 = io_cpu_fence_value & _T & _T_2 ? _GEN_955 : valid_440_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1980 = io_cpu_fence_value & _T & _T_2 ? _GEN_956 : valid_441_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1981 = io_cpu_fence_value & _T & _T_2 ? _GEN_957 : valid_442_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1982 = io_cpu_fence_value & _T & _T_2 ? _GEN_958 : valid_443_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1983 = io_cpu_fence_value & _T & _T_2 ? _GEN_959 : valid_444_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1984 = io_cpu_fence_value & _T & _T_2 ? _GEN_960 : valid_445_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1985 = io_cpu_fence_value & _T & _T_2 ? _GEN_961 : valid_446_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1986 = io_cpu_fence_value & _T & _T_2 ? _GEN_962 : valid_447_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1987 = io_cpu_fence_value & _T & _T_2 ? _GEN_963 : valid_448_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1988 = io_cpu_fence_value & _T & _T_2 ? _GEN_964 : valid_449_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1989 = io_cpu_fence_value & _T & _T_2 ? _GEN_965 : valid_450_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1990 = io_cpu_fence_value & _T & _T_2 ? _GEN_966 : valid_451_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1991 = io_cpu_fence_value & _T & _T_2 ? _GEN_967 : valid_452_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1992 = io_cpu_fence_value & _T & _T_2 ? _GEN_968 : valid_453_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1993 = io_cpu_fence_value & _T & _T_2 ? _GEN_969 : valid_454_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1994 = io_cpu_fence_value & _T & _T_2 ? _GEN_970 : valid_455_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1995 = io_cpu_fence_value & _T & _T_2 ? _GEN_971 : valid_456_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1996 = io_cpu_fence_value & _T & _T_2 ? _GEN_972 : valid_457_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1997 = io_cpu_fence_value & _T & _T_2 ? _GEN_973 : valid_458_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1998 = io_cpu_fence_value & _T & _T_2 ? _GEN_974 : valid_459_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_1999 = io_cpu_fence_value & _T & _T_2 ? _GEN_975 : valid_460_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2000 = io_cpu_fence_value & _T & _T_2 ? _GEN_976 : valid_461_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2001 = io_cpu_fence_value & _T & _T_2 ? _GEN_977 : valid_462_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2002 = io_cpu_fence_value & _T & _T_2 ? _GEN_978 : valid_463_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2003 = io_cpu_fence_value & _T & _T_2 ? _GEN_979 : valid_464_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2004 = io_cpu_fence_value & _T & _T_2 ? _GEN_980 : valid_465_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2005 = io_cpu_fence_value & _T & _T_2 ? _GEN_981 : valid_466_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2006 = io_cpu_fence_value & _T & _T_2 ? _GEN_982 : valid_467_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2007 = io_cpu_fence_value & _T & _T_2 ? _GEN_983 : valid_468_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2008 = io_cpu_fence_value & _T & _T_2 ? _GEN_984 : valid_469_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2009 = io_cpu_fence_value & _T & _T_2 ? _GEN_985 : valid_470_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2010 = io_cpu_fence_value & _T & _T_2 ? _GEN_986 : valid_471_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2011 = io_cpu_fence_value & _T & _T_2 ? _GEN_987 : valid_472_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2012 = io_cpu_fence_value & _T & _T_2 ? _GEN_988 : valid_473_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2013 = io_cpu_fence_value & _T & _T_2 ? _GEN_989 : valid_474_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2014 = io_cpu_fence_value & _T & _T_2 ? _GEN_990 : valid_475_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2015 = io_cpu_fence_value & _T & _T_2 ? _GEN_991 : valid_476_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2016 = io_cpu_fence_value & _T & _T_2 ? _GEN_992 : valid_477_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2017 = io_cpu_fence_value & _T & _T_2 ? _GEN_993 : valid_478_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2018 = io_cpu_fence_value & _T & _T_2 ? _GEN_994 : valid_479_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2019 = io_cpu_fence_value & _T & _T_2 ? _GEN_995 : valid_480_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2020 = io_cpu_fence_value & _T & _T_2 ? _GEN_996 : valid_481_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2021 = io_cpu_fence_value & _T & _T_2 ? _GEN_997 : valid_482_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2022 = io_cpu_fence_value & _T & _T_2 ? _GEN_998 : valid_483_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2023 = io_cpu_fence_value & _T & _T_2 ? _GEN_999 : valid_484_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2024 = io_cpu_fence_value & _T & _T_2 ? _GEN_1000 : valid_485_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2025 = io_cpu_fence_value & _T & _T_2 ? _GEN_1001 : valid_486_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2026 = io_cpu_fence_value & _T & _T_2 ? _GEN_1002 : valid_487_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2027 = io_cpu_fence_value & _T & _T_2 ? _GEN_1003 : valid_488_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2028 = io_cpu_fence_value & _T & _T_2 ? _GEN_1004 : valid_489_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2029 = io_cpu_fence_value & _T & _T_2 ? _GEN_1005 : valid_490_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2030 = io_cpu_fence_value & _T & _T_2 ? _GEN_1006 : valid_491_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2031 = io_cpu_fence_value & _T & _T_2 ? _GEN_1007 : valid_492_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2032 = io_cpu_fence_value & _T & _T_2 ? _GEN_1008 : valid_493_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2033 = io_cpu_fence_value & _T & _T_2 ? _GEN_1009 : valid_494_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2034 = io_cpu_fence_value & _T & _T_2 ? _GEN_1010 : valid_495_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2035 = io_cpu_fence_value & _T & _T_2 ? _GEN_1011 : valid_496_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2036 = io_cpu_fence_value & _T & _T_2 ? _GEN_1012 : valid_497_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2037 = io_cpu_fence_value & _T & _T_2 ? _GEN_1013 : valid_498_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2038 = io_cpu_fence_value & _T & _T_2 ? _GEN_1014 : valid_499_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2039 = io_cpu_fence_value & _T & _T_2 ? _GEN_1015 : valid_500_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2040 = io_cpu_fence_value & _T & _T_2 ? _GEN_1016 : valid_501_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2041 = io_cpu_fence_value & _T & _T_2 ? _GEN_1017 : valid_502_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2042 = io_cpu_fence_value & _T & _T_2 ? _GEN_1018 : valid_503_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2043 = io_cpu_fence_value & _T & _T_2 ? _GEN_1019 : valid_504_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2044 = io_cpu_fence_value & _T & _T_2 ? _GEN_1020 : valid_505_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2045 = io_cpu_fence_value & _T & _T_2 ? _GEN_1021 : valid_506_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2046 = io_cpu_fence_value & _T & _T_2 ? _GEN_1022 : valid_507_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2047 = io_cpu_fence_value & _T & _T_2 ? _GEN_1023 : valid_508_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2048 = io_cpu_fence_value & _T & _T_2 ? _GEN_1024 : valid_509_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2049 = io_cpu_fence_value & _T & _T_2 ? _GEN_1025 : valid_510_1; // @[ICache.scala 52:22 88:73]
  wire  _GEN_2050 = io_cpu_fence_value & _T & _T_2 ? _GEN_1026 : valid_511_1; // @[ICache.scala 52:22 88:73]
  wire  translation_ok = direct_mapped | tlb_vpn == inst_vpn & tlb_valid; // @[ICache.scala 92:38]
  reg [5:0] rset; // @[ICache.scala 95:21]
  wire [5:0] vset = io_cpu_addr_0[11:6]; // @[ICache.scala 98:28]
  wire [19:0] tag_0 = tag_bram_1_io_rdata; // @[ICache.scala 55:18 135:23]
  wire  _GEN_2052 = 6'h1 == vset ? valid_1_0 : valid_0_0; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2053 = 6'h2 == vset ? valid_2_0 : _GEN_2052; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2054 = 6'h3 == vset ? valid_3_0 : _GEN_2053; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2055 = 6'h4 == vset ? valid_4_0 : _GEN_2054; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2056 = 6'h5 == vset ? valid_5_0 : _GEN_2055; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2057 = 6'h6 == vset ? valid_6_0 : _GEN_2056; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2058 = 6'h7 == vset ? valid_7_0 : _GEN_2057; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2059 = 6'h8 == vset ? valid_8_0 : _GEN_2058; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2060 = 6'h9 == vset ? valid_9_0 : _GEN_2059; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2061 = 6'ha == vset ? valid_10_0 : _GEN_2060; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2062 = 6'hb == vset ? valid_11_0 : _GEN_2061; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2063 = 6'hc == vset ? valid_12_0 : _GEN_2062; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2064 = 6'hd == vset ? valid_13_0 : _GEN_2063; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2065 = 6'he == vset ? valid_14_0 : _GEN_2064; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2066 = 6'hf == vset ? valid_15_0 : _GEN_2065; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2067 = 6'h10 == vset ? valid_16_0 : _GEN_2066; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2068 = 6'h11 == vset ? valid_17_0 : _GEN_2067; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2069 = 6'h12 == vset ? valid_18_0 : _GEN_2068; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2070 = 6'h13 == vset ? valid_19_0 : _GEN_2069; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2071 = 6'h14 == vset ? valid_20_0 : _GEN_2070; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2072 = 6'h15 == vset ? valid_21_0 : _GEN_2071; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2073 = 6'h16 == vset ? valid_22_0 : _GEN_2072; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2074 = 6'h17 == vset ? valid_23_0 : _GEN_2073; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2075 = 6'h18 == vset ? valid_24_0 : _GEN_2074; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2076 = 6'h19 == vset ? valid_25_0 : _GEN_2075; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2077 = 6'h1a == vset ? valid_26_0 : _GEN_2076; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2078 = 6'h1b == vset ? valid_27_0 : _GEN_2077; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2079 = 6'h1c == vset ? valid_28_0 : _GEN_2078; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2080 = 6'h1d == vset ? valid_29_0 : _GEN_2079; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2081 = 6'h1e == vset ? valid_30_0 : _GEN_2080; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2082 = 6'h1f == vset ? valid_31_0 : _GEN_2081; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2083 = 6'h20 == vset ? valid_32_0 : _GEN_2082; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2084 = 6'h21 == vset ? valid_33_0 : _GEN_2083; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2085 = 6'h22 == vset ? valid_34_0 : _GEN_2084; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2086 = 6'h23 == vset ? valid_35_0 : _GEN_2085; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2087 = 6'h24 == vset ? valid_36_0 : _GEN_2086; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2088 = 6'h25 == vset ? valid_37_0 : _GEN_2087; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2089 = 6'h26 == vset ? valid_38_0 : _GEN_2088; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2090 = 6'h27 == vset ? valid_39_0 : _GEN_2089; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2091 = 6'h28 == vset ? valid_40_0 : _GEN_2090; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2092 = 6'h29 == vset ? valid_41_0 : _GEN_2091; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2093 = 6'h2a == vset ? valid_42_0 : _GEN_2092; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2094 = 6'h2b == vset ? valid_43_0 : _GEN_2093; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2095 = 6'h2c == vset ? valid_44_0 : _GEN_2094; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2096 = 6'h2d == vset ? valid_45_0 : _GEN_2095; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2097 = 6'h2e == vset ? valid_46_0 : _GEN_2096; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2098 = 6'h2f == vset ? valid_47_0 : _GEN_2097; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2099 = 6'h30 == vset ? valid_48_0 : _GEN_2098; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2100 = 6'h31 == vset ? valid_49_0 : _GEN_2099; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2101 = 6'h32 == vset ? valid_50_0 : _GEN_2100; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2102 = 6'h33 == vset ? valid_51_0 : _GEN_2101; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2103 = 6'h34 == vset ? valid_52_0 : _GEN_2102; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2104 = 6'h35 == vset ? valid_53_0 : _GEN_2103; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2105 = 6'h36 == vset ? valid_54_0 : _GEN_2104; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2106 = 6'h37 == vset ? valid_55_0 : _GEN_2105; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2107 = 6'h38 == vset ? valid_56_0 : _GEN_2106; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2108 = 6'h39 == vset ? valid_57_0 : _GEN_2107; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2109 = 6'h3a == vset ? valid_58_0 : _GEN_2108; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2110 = 6'h3b == vset ? valid_59_0 : _GEN_2109; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2111 = 6'h3c == vset ? valid_60_0 : _GEN_2110; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2112 = 6'h3d == vset ? valid_61_0 : _GEN_2111; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2113 = 6'h3e == vset ? valid_62_0 : _GEN_2112; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2114 = 6'h3f == vset ? valid_63_0 : _GEN_2113; // @[ICache.scala 101:{81,81}]
  wire [6:0] _GEN_14439 = {{1'd0}, vset}; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2115 = 7'h40 == _GEN_14439 ? valid_64_0 : _GEN_2114; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2116 = 7'h41 == _GEN_14439 ? valid_65_0 : _GEN_2115; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2117 = 7'h42 == _GEN_14439 ? valid_66_0 : _GEN_2116; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2118 = 7'h43 == _GEN_14439 ? valid_67_0 : _GEN_2117; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2119 = 7'h44 == _GEN_14439 ? valid_68_0 : _GEN_2118; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2120 = 7'h45 == _GEN_14439 ? valid_69_0 : _GEN_2119; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2121 = 7'h46 == _GEN_14439 ? valid_70_0 : _GEN_2120; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2122 = 7'h47 == _GEN_14439 ? valid_71_0 : _GEN_2121; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2123 = 7'h48 == _GEN_14439 ? valid_72_0 : _GEN_2122; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2124 = 7'h49 == _GEN_14439 ? valid_73_0 : _GEN_2123; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2125 = 7'h4a == _GEN_14439 ? valid_74_0 : _GEN_2124; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2126 = 7'h4b == _GEN_14439 ? valid_75_0 : _GEN_2125; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2127 = 7'h4c == _GEN_14439 ? valid_76_0 : _GEN_2126; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2128 = 7'h4d == _GEN_14439 ? valid_77_0 : _GEN_2127; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2129 = 7'h4e == _GEN_14439 ? valid_78_0 : _GEN_2128; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2130 = 7'h4f == _GEN_14439 ? valid_79_0 : _GEN_2129; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2131 = 7'h50 == _GEN_14439 ? valid_80_0 : _GEN_2130; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2132 = 7'h51 == _GEN_14439 ? valid_81_0 : _GEN_2131; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2133 = 7'h52 == _GEN_14439 ? valid_82_0 : _GEN_2132; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2134 = 7'h53 == _GEN_14439 ? valid_83_0 : _GEN_2133; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2135 = 7'h54 == _GEN_14439 ? valid_84_0 : _GEN_2134; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2136 = 7'h55 == _GEN_14439 ? valid_85_0 : _GEN_2135; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2137 = 7'h56 == _GEN_14439 ? valid_86_0 : _GEN_2136; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2138 = 7'h57 == _GEN_14439 ? valid_87_0 : _GEN_2137; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2139 = 7'h58 == _GEN_14439 ? valid_88_0 : _GEN_2138; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2140 = 7'h59 == _GEN_14439 ? valid_89_0 : _GEN_2139; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2141 = 7'h5a == _GEN_14439 ? valid_90_0 : _GEN_2140; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2142 = 7'h5b == _GEN_14439 ? valid_91_0 : _GEN_2141; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2143 = 7'h5c == _GEN_14439 ? valid_92_0 : _GEN_2142; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2144 = 7'h5d == _GEN_14439 ? valid_93_0 : _GEN_2143; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2145 = 7'h5e == _GEN_14439 ? valid_94_0 : _GEN_2144; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2146 = 7'h5f == _GEN_14439 ? valid_95_0 : _GEN_2145; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2147 = 7'h60 == _GEN_14439 ? valid_96_0 : _GEN_2146; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2148 = 7'h61 == _GEN_14439 ? valid_97_0 : _GEN_2147; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2149 = 7'h62 == _GEN_14439 ? valid_98_0 : _GEN_2148; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2150 = 7'h63 == _GEN_14439 ? valid_99_0 : _GEN_2149; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2151 = 7'h64 == _GEN_14439 ? valid_100_0 : _GEN_2150; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2152 = 7'h65 == _GEN_14439 ? valid_101_0 : _GEN_2151; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2153 = 7'h66 == _GEN_14439 ? valid_102_0 : _GEN_2152; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2154 = 7'h67 == _GEN_14439 ? valid_103_0 : _GEN_2153; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2155 = 7'h68 == _GEN_14439 ? valid_104_0 : _GEN_2154; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2156 = 7'h69 == _GEN_14439 ? valid_105_0 : _GEN_2155; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2157 = 7'h6a == _GEN_14439 ? valid_106_0 : _GEN_2156; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2158 = 7'h6b == _GEN_14439 ? valid_107_0 : _GEN_2157; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2159 = 7'h6c == _GEN_14439 ? valid_108_0 : _GEN_2158; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2160 = 7'h6d == _GEN_14439 ? valid_109_0 : _GEN_2159; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2161 = 7'h6e == _GEN_14439 ? valid_110_0 : _GEN_2160; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2162 = 7'h6f == _GEN_14439 ? valid_111_0 : _GEN_2161; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2163 = 7'h70 == _GEN_14439 ? valid_112_0 : _GEN_2162; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2164 = 7'h71 == _GEN_14439 ? valid_113_0 : _GEN_2163; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2165 = 7'h72 == _GEN_14439 ? valid_114_0 : _GEN_2164; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2166 = 7'h73 == _GEN_14439 ? valid_115_0 : _GEN_2165; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2167 = 7'h74 == _GEN_14439 ? valid_116_0 : _GEN_2166; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2168 = 7'h75 == _GEN_14439 ? valid_117_0 : _GEN_2167; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2169 = 7'h76 == _GEN_14439 ? valid_118_0 : _GEN_2168; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2170 = 7'h77 == _GEN_14439 ? valid_119_0 : _GEN_2169; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2171 = 7'h78 == _GEN_14439 ? valid_120_0 : _GEN_2170; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2172 = 7'h79 == _GEN_14439 ? valid_121_0 : _GEN_2171; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2173 = 7'h7a == _GEN_14439 ? valid_122_0 : _GEN_2172; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2174 = 7'h7b == _GEN_14439 ? valid_123_0 : _GEN_2173; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2175 = 7'h7c == _GEN_14439 ? valid_124_0 : _GEN_2174; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2176 = 7'h7d == _GEN_14439 ? valid_125_0 : _GEN_2175; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2177 = 7'h7e == _GEN_14439 ? valid_126_0 : _GEN_2176; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2178 = 7'h7f == _GEN_14439 ? valid_127_0 : _GEN_2177; // @[ICache.scala 101:{81,81}]
  wire [7:0] _GEN_14503 = {{2'd0}, vset}; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2179 = 8'h80 == _GEN_14503 ? valid_128_0 : _GEN_2178; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2180 = 8'h81 == _GEN_14503 ? valid_129_0 : _GEN_2179; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2181 = 8'h82 == _GEN_14503 ? valid_130_0 : _GEN_2180; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2182 = 8'h83 == _GEN_14503 ? valid_131_0 : _GEN_2181; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2183 = 8'h84 == _GEN_14503 ? valid_132_0 : _GEN_2182; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2184 = 8'h85 == _GEN_14503 ? valid_133_0 : _GEN_2183; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2185 = 8'h86 == _GEN_14503 ? valid_134_0 : _GEN_2184; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2186 = 8'h87 == _GEN_14503 ? valid_135_0 : _GEN_2185; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2187 = 8'h88 == _GEN_14503 ? valid_136_0 : _GEN_2186; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2188 = 8'h89 == _GEN_14503 ? valid_137_0 : _GEN_2187; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2189 = 8'h8a == _GEN_14503 ? valid_138_0 : _GEN_2188; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2190 = 8'h8b == _GEN_14503 ? valid_139_0 : _GEN_2189; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2191 = 8'h8c == _GEN_14503 ? valid_140_0 : _GEN_2190; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2192 = 8'h8d == _GEN_14503 ? valid_141_0 : _GEN_2191; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2193 = 8'h8e == _GEN_14503 ? valid_142_0 : _GEN_2192; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2194 = 8'h8f == _GEN_14503 ? valid_143_0 : _GEN_2193; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2195 = 8'h90 == _GEN_14503 ? valid_144_0 : _GEN_2194; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2196 = 8'h91 == _GEN_14503 ? valid_145_0 : _GEN_2195; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2197 = 8'h92 == _GEN_14503 ? valid_146_0 : _GEN_2196; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2198 = 8'h93 == _GEN_14503 ? valid_147_0 : _GEN_2197; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2199 = 8'h94 == _GEN_14503 ? valid_148_0 : _GEN_2198; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2200 = 8'h95 == _GEN_14503 ? valid_149_0 : _GEN_2199; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2201 = 8'h96 == _GEN_14503 ? valid_150_0 : _GEN_2200; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2202 = 8'h97 == _GEN_14503 ? valid_151_0 : _GEN_2201; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2203 = 8'h98 == _GEN_14503 ? valid_152_0 : _GEN_2202; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2204 = 8'h99 == _GEN_14503 ? valid_153_0 : _GEN_2203; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2205 = 8'h9a == _GEN_14503 ? valid_154_0 : _GEN_2204; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2206 = 8'h9b == _GEN_14503 ? valid_155_0 : _GEN_2205; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2207 = 8'h9c == _GEN_14503 ? valid_156_0 : _GEN_2206; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2208 = 8'h9d == _GEN_14503 ? valid_157_0 : _GEN_2207; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2209 = 8'h9e == _GEN_14503 ? valid_158_0 : _GEN_2208; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2210 = 8'h9f == _GEN_14503 ? valid_159_0 : _GEN_2209; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2211 = 8'ha0 == _GEN_14503 ? valid_160_0 : _GEN_2210; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2212 = 8'ha1 == _GEN_14503 ? valid_161_0 : _GEN_2211; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2213 = 8'ha2 == _GEN_14503 ? valid_162_0 : _GEN_2212; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2214 = 8'ha3 == _GEN_14503 ? valid_163_0 : _GEN_2213; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2215 = 8'ha4 == _GEN_14503 ? valid_164_0 : _GEN_2214; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2216 = 8'ha5 == _GEN_14503 ? valid_165_0 : _GEN_2215; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2217 = 8'ha6 == _GEN_14503 ? valid_166_0 : _GEN_2216; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2218 = 8'ha7 == _GEN_14503 ? valid_167_0 : _GEN_2217; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2219 = 8'ha8 == _GEN_14503 ? valid_168_0 : _GEN_2218; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2220 = 8'ha9 == _GEN_14503 ? valid_169_0 : _GEN_2219; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2221 = 8'haa == _GEN_14503 ? valid_170_0 : _GEN_2220; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2222 = 8'hab == _GEN_14503 ? valid_171_0 : _GEN_2221; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2223 = 8'hac == _GEN_14503 ? valid_172_0 : _GEN_2222; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2224 = 8'had == _GEN_14503 ? valid_173_0 : _GEN_2223; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2225 = 8'hae == _GEN_14503 ? valid_174_0 : _GEN_2224; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2226 = 8'haf == _GEN_14503 ? valid_175_0 : _GEN_2225; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2227 = 8'hb0 == _GEN_14503 ? valid_176_0 : _GEN_2226; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2228 = 8'hb1 == _GEN_14503 ? valid_177_0 : _GEN_2227; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2229 = 8'hb2 == _GEN_14503 ? valid_178_0 : _GEN_2228; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2230 = 8'hb3 == _GEN_14503 ? valid_179_0 : _GEN_2229; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2231 = 8'hb4 == _GEN_14503 ? valid_180_0 : _GEN_2230; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2232 = 8'hb5 == _GEN_14503 ? valid_181_0 : _GEN_2231; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2233 = 8'hb6 == _GEN_14503 ? valid_182_0 : _GEN_2232; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2234 = 8'hb7 == _GEN_14503 ? valid_183_0 : _GEN_2233; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2235 = 8'hb8 == _GEN_14503 ? valid_184_0 : _GEN_2234; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2236 = 8'hb9 == _GEN_14503 ? valid_185_0 : _GEN_2235; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2237 = 8'hba == _GEN_14503 ? valid_186_0 : _GEN_2236; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2238 = 8'hbb == _GEN_14503 ? valid_187_0 : _GEN_2237; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2239 = 8'hbc == _GEN_14503 ? valid_188_0 : _GEN_2238; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2240 = 8'hbd == _GEN_14503 ? valid_189_0 : _GEN_2239; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2241 = 8'hbe == _GEN_14503 ? valid_190_0 : _GEN_2240; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2242 = 8'hbf == _GEN_14503 ? valid_191_0 : _GEN_2241; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2243 = 8'hc0 == _GEN_14503 ? valid_192_0 : _GEN_2242; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2244 = 8'hc1 == _GEN_14503 ? valid_193_0 : _GEN_2243; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2245 = 8'hc2 == _GEN_14503 ? valid_194_0 : _GEN_2244; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2246 = 8'hc3 == _GEN_14503 ? valid_195_0 : _GEN_2245; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2247 = 8'hc4 == _GEN_14503 ? valid_196_0 : _GEN_2246; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2248 = 8'hc5 == _GEN_14503 ? valid_197_0 : _GEN_2247; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2249 = 8'hc6 == _GEN_14503 ? valid_198_0 : _GEN_2248; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2250 = 8'hc7 == _GEN_14503 ? valid_199_0 : _GEN_2249; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2251 = 8'hc8 == _GEN_14503 ? valid_200_0 : _GEN_2250; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2252 = 8'hc9 == _GEN_14503 ? valid_201_0 : _GEN_2251; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2253 = 8'hca == _GEN_14503 ? valid_202_0 : _GEN_2252; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2254 = 8'hcb == _GEN_14503 ? valid_203_0 : _GEN_2253; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2255 = 8'hcc == _GEN_14503 ? valid_204_0 : _GEN_2254; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2256 = 8'hcd == _GEN_14503 ? valid_205_0 : _GEN_2255; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2257 = 8'hce == _GEN_14503 ? valid_206_0 : _GEN_2256; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2258 = 8'hcf == _GEN_14503 ? valid_207_0 : _GEN_2257; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2259 = 8'hd0 == _GEN_14503 ? valid_208_0 : _GEN_2258; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2260 = 8'hd1 == _GEN_14503 ? valid_209_0 : _GEN_2259; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2261 = 8'hd2 == _GEN_14503 ? valid_210_0 : _GEN_2260; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2262 = 8'hd3 == _GEN_14503 ? valid_211_0 : _GEN_2261; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2263 = 8'hd4 == _GEN_14503 ? valid_212_0 : _GEN_2262; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2264 = 8'hd5 == _GEN_14503 ? valid_213_0 : _GEN_2263; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2265 = 8'hd6 == _GEN_14503 ? valid_214_0 : _GEN_2264; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2266 = 8'hd7 == _GEN_14503 ? valid_215_0 : _GEN_2265; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2267 = 8'hd8 == _GEN_14503 ? valid_216_0 : _GEN_2266; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2268 = 8'hd9 == _GEN_14503 ? valid_217_0 : _GEN_2267; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2269 = 8'hda == _GEN_14503 ? valid_218_0 : _GEN_2268; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2270 = 8'hdb == _GEN_14503 ? valid_219_0 : _GEN_2269; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2271 = 8'hdc == _GEN_14503 ? valid_220_0 : _GEN_2270; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2272 = 8'hdd == _GEN_14503 ? valid_221_0 : _GEN_2271; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2273 = 8'hde == _GEN_14503 ? valid_222_0 : _GEN_2272; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2274 = 8'hdf == _GEN_14503 ? valid_223_0 : _GEN_2273; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2275 = 8'he0 == _GEN_14503 ? valid_224_0 : _GEN_2274; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2276 = 8'he1 == _GEN_14503 ? valid_225_0 : _GEN_2275; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2277 = 8'he2 == _GEN_14503 ? valid_226_0 : _GEN_2276; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2278 = 8'he3 == _GEN_14503 ? valid_227_0 : _GEN_2277; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2279 = 8'he4 == _GEN_14503 ? valid_228_0 : _GEN_2278; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2280 = 8'he5 == _GEN_14503 ? valid_229_0 : _GEN_2279; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2281 = 8'he6 == _GEN_14503 ? valid_230_0 : _GEN_2280; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2282 = 8'he7 == _GEN_14503 ? valid_231_0 : _GEN_2281; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2283 = 8'he8 == _GEN_14503 ? valid_232_0 : _GEN_2282; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2284 = 8'he9 == _GEN_14503 ? valid_233_0 : _GEN_2283; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2285 = 8'hea == _GEN_14503 ? valid_234_0 : _GEN_2284; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2286 = 8'heb == _GEN_14503 ? valid_235_0 : _GEN_2285; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2287 = 8'hec == _GEN_14503 ? valid_236_0 : _GEN_2286; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2288 = 8'hed == _GEN_14503 ? valid_237_0 : _GEN_2287; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2289 = 8'hee == _GEN_14503 ? valid_238_0 : _GEN_2288; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2290 = 8'hef == _GEN_14503 ? valid_239_0 : _GEN_2289; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2291 = 8'hf0 == _GEN_14503 ? valid_240_0 : _GEN_2290; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2292 = 8'hf1 == _GEN_14503 ? valid_241_0 : _GEN_2291; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2293 = 8'hf2 == _GEN_14503 ? valid_242_0 : _GEN_2292; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2294 = 8'hf3 == _GEN_14503 ? valid_243_0 : _GEN_2293; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2295 = 8'hf4 == _GEN_14503 ? valid_244_0 : _GEN_2294; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2296 = 8'hf5 == _GEN_14503 ? valid_245_0 : _GEN_2295; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2297 = 8'hf6 == _GEN_14503 ? valid_246_0 : _GEN_2296; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2298 = 8'hf7 == _GEN_14503 ? valid_247_0 : _GEN_2297; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2299 = 8'hf8 == _GEN_14503 ? valid_248_0 : _GEN_2298; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2300 = 8'hf9 == _GEN_14503 ? valid_249_0 : _GEN_2299; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2301 = 8'hfa == _GEN_14503 ? valid_250_0 : _GEN_2300; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2302 = 8'hfb == _GEN_14503 ? valid_251_0 : _GEN_2301; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2303 = 8'hfc == _GEN_14503 ? valid_252_0 : _GEN_2302; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2304 = 8'hfd == _GEN_14503 ? valid_253_0 : _GEN_2303; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2305 = 8'hfe == _GEN_14503 ? valid_254_0 : _GEN_2304; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2306 = 8'hff == _GEN_14503 ? valid_255_0 : _GEN_2305; // @[ICache.scala 101:{81,81}]
  wire [8:0] _GEN_14631 = {{3'd0}, vset}; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2307 = 9'h100 == _GEN_14631 ? valid_256_0 : _GEN_2306; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2308 = 9'h101 == _GEN_14631 ? valid_257_0 : _GEN_2307; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2309 = 9'h102 == _GEN_14631 ? valid_258_0 : _GEN_2308; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2310 = 9'h103 == _GEN_14631 ? valid_259_0 : _GEN_2309; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2311 = 9'h104 == _GEN_14631 ? valid_260_0 : _GEN_2310; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2312 = 9'h105 == _GEN_14631 ? valid_261_0 : _GEN_2311; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2313 = 9'h106 == _GEN_14631 ? valid_262_0 : _GEN_2312; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2314 = 9'h107 == _GEN_14631 ? valid_263_0 : _GEN_2313; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2315 = 9'h108 == _GEN_14631 ? valid_264_0 : _GEN_2314; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2316 = 9'h109 == _GEN_14631 ? valid_265_0 : _GEN_2315; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2317 = 9'h10a == _GEN_14631 ? valid_266_0 : _GEN_2316; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2318 = 9'h10b == _GEN_14631 ? valid_267_0 : _GEN_2317; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2319 = 9'h10c == _GEN_14631 ? valid_268_0 : _GEN_2318; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2320 = 9'h10d == _GEN_14631 ? valid_269_0 : _GEN_2319; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2321 = 9'h10e == _GEN_14631 ? valid_270_0 : _GEN_2320; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2322 = 9'h10f == _GEN_14631 ? valid_271_0 : _GEN_2321; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2323 = 9'h110 == _GEN_14631 ? valid_272_0 : _GEN_2322; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2324 = 9'h111 == _GEN_14631 ? valid_273_0 : _GEN_2323; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2325 = 9'h112 == _GEN_14631 ? valid_274_0 : _GEN_2324; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2326 = 9'h113 == _GEN_14631 ? valid_275_0 : _GEN_2325; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2327 = 9'h114 == _GEN_14631 ? valid_276_0 : _GEN_2326; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2328 = 9'h115 == _GEN_14631 ? valid_277_0 : _GEN_2327; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2329 = 9'h116 == _GEN_14631 ? valid_278_0 : _GEN_2328; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2330 = 9'h117 == _GEN_14631 ? valid_279_0 : _GEN_2329; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2331 = 9'h118 == _GEN_14631 ? valid_280_0 : _GEN_2330; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2332 = 9'h119 == _GEN_14631 ? valid_281_0 : _GEN_2331; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2333 = 9'h11a == _GEN_14631 ? valid_282_0 : _GEN_2332; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2334 = 9'h11b == _GEN_14631 ? valid_283_0 : _GEN_2333; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2335 = 9'h11c == _GEN_14631 ? valid_284_0 : _GEN_2334; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2336 = 9'h11d == _GEN_14631 ? valid_285_0 : _GEN_2335; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2337 = 9'h11e == _GEN_14631 ? valid_286_0 : _GEN_2336; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2338 = 9'h11f == _GEN_14631 ? valid_287_0 : _GEN_2337; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2339 = 9'h120 == _GEN_14631 ? valid_288_0 : _GEN_2338; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2340 = 9'h121 == _GEN_14631 ? valid_289_0 : _GEN_2339; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2341 = 9'h122 == _GEN_14631 ? valid_290_0 : _GEN_2340; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2342 = 9'h123 == _GEN_14631 ? valid_291_0 : _GEN_2341; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2343 = 9'h124 == _GEN_14631 ? valid_292_0 : _GEN_2342; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2344 = 9'h125 == _GEN_14631 ? valid_293_0 : _GEN_2343; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2345 = 9'h126 == _GEN_14631 ? valid_294_0 : _GEN_2344; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2346 = 9'h127 == _GEN_14631 ? valid_295_0 : _GEN_2345; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2347 = 9'h128 == _GEN_14631 ? valid_296_0 : _GEN_2346; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2348 = 9'h129 == _GEN_14631 ? valid_297_0 : _GEN_2347; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2349 = 9'h12a == _GEN_14631 ? valid_298_0 : _GEN_2348; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2350 = 9'h12b == _GEN_14631 ? valid_299_0 : _GEN_2349; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2351 = 9'h12c == _GEN_14631 ? valid_300_0 : _GEN_2350; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2352 = 9'h12d == _GEN_14631 ? valid_301_0 : _GEN_2351; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2353 = 9'h12e == _GEN_14631 ? valid_302_0 : _GEN_2352; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2354 = 9'h12f == _GEN_14631 ? valid_303_0 : _GEN_2353; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2355 = 9'h130 == _GEN_14631 ? valid_304_0 : _GEN_2354; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2356 = 9'h131 == _GEN_14631 ? valid_305_0 : _GEN_2355; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2357 = 9'h132 == _GEN_14631 ? valid_306_0 : _GEN_2356; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2358 = 9'h133 == _GEN_14631 ? valid_307_0 : _GEN_2357; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2359 = 9'h134 == _GEN_14631 ? valid_308_0 : _GEN_2358; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2360 = 9'h135 == _GEN_14631 ? valid_309_0 : _GEN_2359; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2361 = 9'h136 == _GEN_14631 ? valid_310_0 : _GEN_2360; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2362 = 9'h137 == _GEN_14631 ? valid_311_0 : _GEN_2361; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2363 = 9'h138 == _GEN_14631 ? valid_312_0 : _GEN_2362; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2364 = 9'h139 == _GEN_14631 ? valid_313_0 : _GEN_2363; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2365 = 9'h13a == _GEN_14631 ? valid_314_0 : _GEN_2364; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2366 = 9'h13b == _GEN_14631 ? valid_315_0 : _GEN_2365; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2367 = 9'h13c == _GEN_14631 ? valid_316_0 : _GEN_2366; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2368 = 9'h13d == _GEN_14631 ? valid_317_0 : _GEN_2367; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2369 = 9'h13e == _GEN_14631 ? valid_318_0 : _GEN_2368; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2370 = 9'h13f == _GEN_14631 ? valid_319_0 : _GEN_2369; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2371 = 9'h140 == _GEN_14631 ? valid_320_0 : _GEN_2370; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2372 = 9'h141 == _GEN_14631 ? valid_321_0 : _GEN_2371; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2373 = 9'h142 == _GEN_14631 ? valid_322_0 : _GEN_2372; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2374 = 9'h143 == _GEN_14631 ? valid_323_0 : _GEN_2373; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2375 = 9'h144 == _GEN_14631 ? valid_324_0 : _GEN_2374; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2376 = 9'h145 == _GEN_14631 ? valid_325_0 : _GEN_2375; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2377 = 9'h146 == _GEN_14631 ? valid_326_0 : _GEN_2376; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2378 = 9'h147 == _GEN_14631 ? valid_327_0 : _GEN_2377; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2379 = 9'h148 == _GEN_14631 ? valid_328_0 : _GEN_2378; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2380 = 9'h149 == _GEN_14631 ? valid_329_0 : _GEN_2379; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2381 = 9'h14a == _GEN_14631 ? valid_330_0 : _GEN_2380; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2382 = 9'h14b == _GEN_14631 ? valid_331_0 : _GEN_2381; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2383 = 9'h14c == _GEN_14631 ? valid_332_0 : _GEN_2382; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2384 = 9'h14d == _GEN_14631 ? valid_333_0 : _GEN_2383; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2385 = 9'h14e == _GEN_14631 ? valid_334_0 : _GEN_2384; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2386 = 9'h14f == _GEN_14631 ? valid_335_0 : _GEN_2385; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2387 = 9'h150 == _GEN_14631 ? valid_336_0 : _GEN_2386; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2388 = 9'h151 == _GEN_14631 ? valid_337_0 : _GEN_2387; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2389 = 9'h152 == _GEN_14631 ? valid_338_0 : _GEN_2388; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2390 = 9'h153 == _GEN_14631 ? valid_339_0 : _GEN_2389; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2391 = 9'h154 == _GEN_14631 ? valid_340_0 : _GEN_2390; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2392 = 9'h155 == _GEN_14631 ? valid_341_0 : _GEN_2391; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2393 = 9'h156 == _GEN_14631 ? valid_342_0 : _GEN_2392; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2394 = 9'h157 == _GEN_14631 ? valid_343_0 : _GEN_2393; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2395 = 9'h158 == _GEN_14631 ? valid_344_0 : _GEN_2394; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2396 = 9'h159 == _GEN_14631 ? valid_345_0 : _GEN_2395; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2397 = 9'h15a == _GEN_14631 ? valid_346_0 : _GEN_2396; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2398 = 9'h15b == _GEN_14631 ? valid_347_0 : _GEN_2397; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2399 = 9'h15c == _GEN_14631 ? valid_348_0 : _GEN_2398; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2400 = 9'h15d == _GEN_14631 ? valid_349_0 : _GEN_2399; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2401 = 9'h15e == _GEN_14631 ? valid_350_0 : _GEN_2400; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2402 = 9'h15f == _GEN_14631 ? valid_351_0 : _GEN_2401; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2403 = 9'h160 == _GEN_14631 ? valid_352_0 : _GEN_2402; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2404 = 9'h161 == _GEN_14631 ? valid_353_0 : _GEN_2403; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2405 = 9'h162 == _GEN_14631 ? valid_354_0 : _GEN_2404; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2406 = 9'h163 == _GEN_14631 ? valid_355_0 : _GEN_2405; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2407 = 9'h164 == _GEN_14631 ? valid_356_0 : _GEN_2406; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2408 = 9'h165 == _GEN_14631 ? valid_357_0 : _GEN_2407; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2409 = 9'h166 == _GEN_14631 ? valid_358_0 : _GEN_2408; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2410 = 9'h167 == _GEN_14631 ? valid_359_0 : _GEN_2409; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2411 = 9'h168 == _GEN_14631 ? valid_360_0 : _GEN_2410; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2412 = 9'h169 == _GEN_14631 ? valid_361_0 : _GEN_2411; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2413 = 9'h16a == _GEN_14631 ? valid_362_0 : _GEN_2412; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2414 = 9'h16b == _GEN_14631 ? valid_363_0 : _GEN_2413; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2415 = 9'h16c == _GEN_14631 ? valid_364_0 : _GEN_2414; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2416 = 9'h16d == _GEN_14631 ? valid_365_0 : _GEN_2415; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2417 = 9'h16e == _GEN_14631 ? valid_366_0 : _GEN_2416; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2418 = 9'h16f == _GEN_14631 ? valid_367_0 : _GEN_2417; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2419 = 9'h170 == _GEN_14631 ? valid_368_0 : _GEN_2418; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2420 = 9'h171 == _GEN_14631 ? valid_369_0 : _GEN_2419; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2421 = 9'h172 == _GEN_14631 ? valid_370_0 : _GEN_2420; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2422 = 9'h173 == _GEN_14631 ? valid_371_0 : _GEN_2421; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2423 = 9'h174 == _GEN_14631 ? valid_372_0 : _GEN_2422; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2424 = 9'h175 == _GEN_14631 ? valid_373_0 : _GEN_2423; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2425 = 9'h176 == _GEN_14631 ? valid_374_0 : _GEN_2424; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2426 = 9'h177 == _GEN_14631 ? valid_375_0 : _GEN_2425; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2427 = 9'h178 == _GEN_14631 ? valid_376_0 : _GEN_2426; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2428 = 9'h179 == _GEN_14631 ? valid_377_0 : _GEN_2427; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2429 = 9'h17a == _GEN_14631 ? valid_378_0 : _GEN_2428; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2430 = 9'h17b == _GEN_14631 ? valid_379_0 : _GEN_2429; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2431 = 9'h17c == _GEN_14631 ? valid_380_0 : _GEN_2430; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2432 = 9'h17d == _GEN_14631 ? valid_381_0 : _GEN_2431; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2433 = 9'h17e == _GEN_14631 ? valid_382_0 : _GEN_2432; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2434 = 9'h17f == _GEN_14631 ? valid_383_0 : _GEN_2433; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2435 = 9'h180 == _GEN_14631 ? valid_384_0 : _GEN_2434; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2436 = 9'h181 == _GEN_14631 ? valid_385_0 : _GEN_2435; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2437 = 9'h182 == _GEN_14631 ? valid_386_0 : _GEN_2436; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2438 = 9'h183 == _GEN_14631 ? valid_387_0 : _GEN_2437; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2439 = 9'h184 == _GEN_14631 ? valid_388_0 : _GEN_2438; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2440 = 9'h185 == _GEN_14631 ? valid_389_0 : _GEN_2439; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2441 = 9'h186 == _GEN_14631 ? valid_390_0 : _GEN_2440; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2442 = 9'h187 == _GEN_14631 ? valid_391_0 : _GEN_2441; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2443 = 9'h188 == _GEN_14631 ? valid_392_0 : _GEN_2442; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2444 = 9'h189 == _GEN_14631 ? valid_393_0 : _GEN_2443; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2445 = 9'h18a == _GEN_14631 ? valid_394_0 : _GEN_2444; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2446 = 9'h18b == _GEN_14631 ? valid_395_0 : _GEN_2445; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2447 = 9'h18c == _GEN_14631 ? valid_396_0 : _GEN_2446; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2448 = 9'h18d == _GEN_14631 ? valid_397_0 : _GEN_2447; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2449 = 9'h18e == _GEN_14631 ? valid_398_0 : _GEN_2448; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2450 = 9'h18f == _GEN_14631 ? valid_399_0 : _GEN_2449; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2451 = 9'h190 == _GEN_14631 ? valid_400_0 : _GEN_2450; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2452 = 9'h191 == _GEN_14631 ? valid_401_0 : _GEN_2451; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2453 = 9'h192 == _GEN_14631 ? valid_402_0 : _GEN_2452; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2454 = 9'h193 == _GEN_14631 ? valid_403_0 : _GEN_2453; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2455 = 9'h194 == _GEN_14631 ? valid_404_0 : _GEN_2454; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2456 = 9'h195 == _GEN_14631 ? valid_405_0 : _GEN_2455; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2457 = 9'h196 == _GEN_14631 ? valid_406_0 : _GEN_2456; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2458 = 9'h197 == _GEN_14631 ? valid_407_0 : _GEN_2457; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2459 = 9'h198 == _GEN_14631 ? valid_408_0 : _GEN_2458; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2460 = 9'h199 == _GEN_14631 ? valid_409_0 : _GEN_2459; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2461 = 9'h19a == _GEN_14631 ? valid_410_0 : _GEN_2460; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2462 = 9'h19b == _GEN_14631 ? valid_411_0 : _GEN_2461; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2463 = 9'h19c == _GEN_14631 ? valid_412_0 : _GEN_2462; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2464 = 9'h19d == _GEN_14631 ? valid_413_0 : _GEN_2463; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2465 = 9'h19e == _GEN_14631 ? valid_414_0 : _GEN_2464; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2466 = 9'h19f == _GEN_14631 ? valid_415_0 : _GEN_2465; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2467 = 9'h1a0 == _GEN_14631 ? valid_416_0 : _GEN_2466; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2468 = 9'h1a1 == _GEN_14631 ? valid_417_0 : _GEN_2467; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2469 = 9'h1a2 == _GEN_14631 ? valid_418_0 : _GEN_2468; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2470 = 9'h1a3 == _GEN_14631 ? valid_419_0 : _GEN_2469; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2471 = 9'h1a4 == _GEN_14631 ? valid_420_0 : _GEN_2470; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2472 = 9'h1a5 == _GEN_14631 ? valid_421_0 : _GEN_2471; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2473 = 9'h1a6 == _GEN_14631 ? valid_422_0 : _GEN_2472; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2474 = 9'h1a7 == _GEN_14631 ? valid_423_0 : _GEN_2473; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2475 = 9'h1a8 == _GEN_14631 ? valid_424_0 : _GEN_2474; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2476 = 9'h1a9 == _GEN_14631 ? valid_425_0 : _GEN_2475; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2477 = 9'h1aa == _GEN_14631 ? valid_426_0 : _GEN_2476; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2478 = 9'h1ab == _GEN_14631 ? valid_427_0 : _GEN_2477; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2479 = 9'h1ac == _GEN_14631 ? valid_428_0 : _GEN_2478; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2480 = 9'h1ad == _GEN_14631 ? valid_429_0 : _GEN_2479; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2481 = 9'h1ae == _GEN_14631 ? valid_430_0 : _GEN_2480; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2482 = 9'h1af == _GEN_14631 ? valid_431_0 : _GEN_2481; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2483 = 9'h1b0 == _GEN_14631 ? valid_432_0 : _GEN_2482; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2484 = 9'h1b1 == _GEN_14631 ? valid_433_0 : _GEN_2483; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2485 = 9'h1b2 == _GEN_14631 ? valid_434_0 : _GEN_2484; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2486 = 9'h1b3 == _GEN_14631 ? valid_435_0 : _GEN_2485; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2487 = 9'h1b4 == _GEN_14631 ? valid_436_0 : _GEN_2486; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2488 = 9'h1b5 == _GEN_14631 ? valid_437_0 : _GEN_2487; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2489 = 9'h1b6 == _GEN_14631 ? valid_438_0 : _GEN_2488; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2490 = 9'h1b7 == _GEN_14631 ? valid_439_0 : _GEN_2489; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2491 = 9'h1b8 == _GEN_14631 ? valid_440_0 : _GEN_2490; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2492 = 9'h1b9 == _GEN_14631 ? valid_441_0 : _GEN_2491; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2493 = 9'h1ba == _GEN_14631 ? valid_442_0 : _GEN_2492; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2494 = 9'h1bb == _GEN_14631 ? valid_443_0 : _GEN_2493; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2495 = 9'h1bc == _GEN_14631 ? valid_444_0 : _GEN_2494; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2496 = 9'h1bd == _GEN_14631 ? valid_445_0 : _GEN_2495; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2497 = 9'h1be == _GEN_14631 ? valid_446_0 : _GEN_2496; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2498 = 9'h1bf == _GEN_14631 ? valid_447_0 : _GEN_2497; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2499 = 9'h1c0 == _GEN_14631 ? valid_448_0 : _GEN_2498; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2500 = 9'h1c1 == _GEN_14631 ? valid_449_0 : _GEN_2499; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2501 = 9'h1c2 == _GEN_14631 ? valid_450_0 : _GEN_2500; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2502 = 9'h1c3 == _GEN_14631 ? valid_451_0 : _GEN_2501; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2503 = 9'h1c4 == _GEN_14631 ? valid_452_0 : _GEN_2502; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2504 = 9'h1c5 == _GEN_14631 ? valid_453_0 : _GEN_2503; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2505 = 9'h1c6 == _GEN_14631 ? valid_454_0 : _GEN_2504; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2506 = 9'h1c7 == _GEN_14631 ? valid_455_0 : _GEN_2505; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2507 = 9'h1c8 == _GEN_14631 ? valid_456_0 : _GEN_2506; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2508 = 9'h1c9 == _GEN_14631 ? valid_457_0 : _GEN_2507; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2509 = 9'h1ca == _GEN_14631 ? valid_458_0 : _GEN_2508; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2510 = 9'h1cb == _GEN_14631 ? valid_459_0 : _GEN_2509; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2511 = 9'h1cc == _GEN_14631 ? valid_460_0 : _GEN_2510; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2512 = 9'h1cd == _GEN_14631 ? valid_461_0 : _GEN_2511; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2513 = 9'h1ce == _GEN_14631 ? valid_462_0 : _GEN_2512; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2514 = 9'h1cf == _GEN_14631 ? valid_463_0 : _GEN_2513; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2515 = 9'h1d0 == _GEN_14631 ? valid_464_0 : _GEN_2514; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2516 = 9'h1d1 == _GEN_14631 ? valid_465_0 : _GEN_2515; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2517 = 9'h1d2 == _GEN_14631 ? valid_466_0 : _GEN_2516; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2518 = 9'h1d3 == _GEN_14631 ? valid_467_0 : _GEN_2517; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2519 = 9'h1d4 == _GEN_14631 ? valid_468_0 : _GEN_2518; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2520 = 9'h1d5 == _GEN_14631 ? valid_469_0 : _GEN_2519; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2521 = 9'h1d6 == _GEN_14631 ? valid_470_0 : _GEN_2520; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2522 = 9'h1d7 == _GEN_14631 ? valid_471_0 : _GEN_2521; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2523 = 9'h1d8 == _GEN_14631 ? valid_472_0 : _GEN_2522; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2524 = 9'h1d9 == _GEN_14631 ? valid_473_0 : _GEN_2523; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2525 = 9'h1da == _GEN_14631 ? valid_474_0 : _GEN_2524; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2526 = 9'h1db == _GEN_14631 ? valid_475_0 : _GEN_2525; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2527 = 9'h1dc == _GEN_14631 ? valid_476_0 : _GEN_2526; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2528 = 9'h1dd == _GEN_14631 ? valid_477_0 : _GEN_2527; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2529 = 9'h1de == _GEN_14631 ? valid_478_0 : _GEN_2528; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2530 = 9'h1df == _GEN_14631 ? valid_479_0 : _GEN_2529; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2531 = 9'h1e0 == _GEN_14631 ? valid_480_0 : _GEN_2530; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2532 = 9'h1e1 == _GEN_14631 ? valid_481_0 : _GEN_2531; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2533 = 9'h1e2 == _GEN_14631 ? valid_482_0 : _GEN_2532; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2534 = 9'h1e3 == _GEN_14631 ? valid_483_0 : _GEN_2533; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2535 = 9'h1e4 == _GEN_14631 ? valid_484_0 : _GEN_2534; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2536 = 9'h1e5 == _GEN_14631 ? valid_485_0 : _GEN_2535; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2537 = 9'h1e6 == _GEN_14631 ? valid_486_0 : _GEN_2536; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2538 = 9'h1e7 == _GEN_14631 ? valid_487_0 : _GEN_2537; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2539 = 9'h1e8 == _GEN_14631 ? valid_488_0 : _GEN_2538; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2540 = 9'h1e9 == _GEN_14631 ? valid_489_0 : _GEN_2539; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2541 = 9'h1ea == _GEN_14631 ? valid_490_0 : _GEN_2540; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2542 = 9'h1eb == _GEN_14631 ? valid_491_0 : _GEN_2541; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2543 = 9'h1ec == _GEN_14631 ? valid_492_0 : _GEN_2542; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2544 = 9'h1ed == _GEN_14631 ? valid_493_0 : _GEN_2543; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2545 = 9'h1ee == _GEN_14631 ? valid_494_0 : _GEN_2544; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2546 = 9'h1ef == _GEN_14631 ? valid_495_0 : _GEN_2545; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2547 = 9'h1f0 == _GEN_14631 ? valid_496_0 : _GEN_2546; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2548 = 9'h1f1 == _GEN_14631 ? valid_497_0 : _GEN_2547; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2549 = 9'h1f2 == _GEN_14631 ? valid_498_0 : _GEN_2548; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2550 = 9'h1f3 == _GEN_14631 ? valid_499_0 : _GEN_2549; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2551 = 9'h1f4 == _GEN_14631 ? valid_500_0 : _GEN_2550; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2552 = 9'h1f5 == _GEN_14631 ? valid_501_0 : _GEN_2551; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2553 = 9'h1f6 == _GEN_14631 ? valid_502_0 : _GEN_2552; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2554 = 9'h1f7 == _GEN_14631 ? valid_503_0 : _GEN_2553; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2555 = 9'h1f8 == _GEN_14631 ? valid_504_0 : _GEN_2554; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2556 = 9'h1f9 == _GEN_14631 ? valid_505_0 : _GEN_2555; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2557 = 9'h1fa == _GEN_14631 ? valid_506_0 : _GEN_2556; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2558 = 9'h1fb == _GEN_14631 ? valid_507_0 : _GEN_2557; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2559 = 9'h1fc == _GEN_14631 ? valid_508_0 : _GEN_2558; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2560 = 9'h1fd == _GEN_14631 ? valid_509_0 : _GEN_2559; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2561 = 9'h1fe == _GEN_14631 ? valid_510_0 : _GEN_2560; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2562 = 9'h1ff == _GEN_14631 ? valid_511_0 : _GEN_2561; // @[ICache.scala 101:{81,81}]
  wire  tag_compare_valid_0 = tag_0 == inst_tag & _GEN_2562; // @[ICache.scala 101:81]
  wire [19:0] tag_1 = tag_bram_3_io_rdata; // @[ICache.scala 55:18 135:23]
  wire  _GEN_2564 = 6'h1 == vset ? valid_1_1 : valid_0_1; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2565 = 6'h2 == vset ? valid_2_1 : _GEN_2564; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2566 = 6'h3 == vset ? valid_3_1 : _GEN_2565; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2567 = 6'h4 == vset ? valid_4_1 : _GEN_2566; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2568 = 6'h5 == vset ? valid_5_1 : _GEN_2567; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2569 = 6'h6 == vset ? valid_6_1 : _GEN_2568; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2570 = 6'h7 == vset ? valid_7_1 : _GEN_2569; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2571 = 6'h8 == vset ? valid_8_1 : _GEN_2570; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2572 = 6'h9 == vset ? valid_9_1 : _GEN_2571; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2573 = 6'ha == vset ? valid_10_1 : _GEN_2572; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2574 = 6'hb == vset ? valid_11_1 : _GEN_2573; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2575 = 6'hc == vset ? valid_12_1 : _GEN_2574; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2576 = 6'hd == vset ? valid_13_1 : _GEN_2575; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2577 = 6'he == vset ? valid_14_1 : _GEN_2576; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2578 = 6'hf == vset ? valid_15_1 : _GEN_2577; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2579 = 6'h10 == vset ? valid_16_1 : _GEN_2578; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2580 = 6'h11 == vset ? valid_17_1 : _GEN_2579; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2581 = 6'h12 == vset ? valid_18_1 : _GEN_2580; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2582 = 6'h13 == vset ? valid_19_1 : _GEN_2581; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2583 = 6'h14 == vset ? valid_20_1 : _GEN_2582; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2584 = 6'h15 == vset ? valid_21_1 : _GEN_2583; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2585 = 6'h16 == vset ? valid_22_1 : _GEN_2584; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2586 = 6'h17 == vset ? valid_23_1 : _GEN_2585; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2587 = 6'h18 == vset ? valid_24_1 : _GEN_2586; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2588 = 6'h19 == vset ? valid_25_1 : _GEN_2587; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2589 = 6'h1a == vset ? valid_26_1 : _GEN_2588; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2590 = 6'h1b == vset ? valid_27_1 : _GEN_2589; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2591 = 6'h1c == vset ? valid_28_1 : _GEN_2590; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2592 = 6'h1d == vset ? valid_29_1 : _GEN_2591; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2593 = 6'h1e == vset ? valid_30_1 : _GEN_2592; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2594 = 6'h1f == vset ? valid_31_1 : _GEN_2593; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2595 = 6'h20 == vset ? valid_32_1 : _GEN_2594; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2596 = 6'h21 == vset ? valid_33_1 : _GEN_2595; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2597 = 6'h22 == vset ? valid_34_1 : _GEN_2596; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2598 = 6'h23 == vset ? valid_35_1 : _GEN_2597; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2599 = 6'h24 == vset ? valid_36_1 : _GEN_2598; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2600 = 6'h25 == vset ? valid_37_1 : _GEN_2599; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2601 = 6'h26 == vset ? valid_38_1 : _GEN_2600; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2602 = 6'h27 == vset ? valid_39_1 : _GEN_2601; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2603 = 6'h28 == vset ? valid_40_1 : _GEN_2602; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2604 = 6'h29 == vset ? valid_41_1 : _GEN_2603; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2605 = 6'h2a == vset ? valid_42_1 : _GEN_2604; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2606 = 6'h2b == vset ? valid_43_1 : _GEN_2605; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2607 = 6'h2c == vset ? valid_44_1 : _GEN_2606; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2608 = 6'h2d == vset ? valid_45_1 : _GEN_2607; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2609 = 6'h2e == vset ? valid_46_1 : _GEN_2608; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2610 = 6'h2f == vset ? valid_47_1 : _GEN_2609; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2611 = 6'h30 == vset ? valid_48_1 : _GEN_2610; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2612 = 6'h31 == vset ? valid_49_1 : _GEN_2611; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2613 = 6'h32 == vset ? valid_50_1 : _GEN_2612; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2614 = 6'h33 == vset ? valid_51_1 : _GEN_2613; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2615 = 6'h34 == vset ? valid_52_1 : _GEN_2614; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2616 = 6'h35 == vset ? valid_53_1 : _GEN_2615; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2617 = 6'h36 == vset ? valid_54_1 : _GEN_2616; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2618 = 6'h37 == vset ? valid_55_1 : _GEN_2617; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2619 = 6'h38 == vset ? valid_56_1 : _GEN_2618; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2620 = 6'h39 == vset ? valid_57_1 : _GEN_2619; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2621 = 6'h3a == vset ? valid_58_1 : _GEN_2620; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2622 = 6'h3b == vset ? valid_59_1 : _GEN_2621; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2623 = 6'h3c == vset ? valid_60_1 : _GEN_2622; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2624 = 6'h3d == vset ? valid_61_1 : _GEN_2623; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2625 = 6'h3e == vset ? valid_62_1 : _GEN_2624; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2626 = 6'h3f == vset ? valid_63_1 : _GEN_2625; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2627 = 7'h40 == _GEN_14439 ? valid_64_1 : _GEN_2626; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2628 = 7'h41 == _GEN_14439 ? valid_65_1 : _GEN_2627; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2629 = 7'h42 == _GEN_14439 ? valid_66_1 : _GEN_2628; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2630 = 7'h43 == _GEN_14439 ? valid_67_1 : _GEN_2629; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2631 = 7'h44 == _GEN_14439 ? valid_68_1 : _GEN_2630; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2632 = 7'h45 == _GEN_14439 ? valid_69_1 : _GEN_2631; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2633 = 7'h46 == _GEN_14439 ? valid_70_1 : _GEN_2632; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2634 = 7'h47 == _GEN_14439 ? valid_71_1 : _GEN_2633; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2635 = 7'h48 == _GEN_14439 ? valid_72_1 : _GEN_2634; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2636 = 7'h49 == _GEN_14439 ? valid_73_1 : _GEN_2635; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2637 = 7'h4a == _GEN_14439 ? valid_74_1 : _GEN_2636; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2638 = 7'h4b == _GEN_14439 ? valid_75_1 : _GEN_2637; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2639 = 7'h4c == _GEN_14439 ? valid_76_1 : _GEN_2638; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2640 = 7'h4d == _GEN_14439 ? valid_77_1 : _GEN_2639; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2641 = 7'h4e == _GEN_14439 ? valid_78_1 : _GEN_2640; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2642 = 7'h4f == _GEN_14439 ? valid_79_1 : _GEN_2641; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2643 = 7'h50 == _GEN_14439 ? valid_80_1 : _GEN_2642; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2644 = 7'h51 == _GEN_14439 ? valid_81_1 : _GEN_2643; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2645 = 7'h52 == _GEN_14439 ? valid_82_1 : _GEN_2644; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2646 = 7'h53 == _GEN_14439 ? valid_83_1 : _GEN_2645; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2647 = 7'h54 == _GEN_14439 ? valid_84_1 : _GEN_2646; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2648 = 7'h55 == _GEN_14439 ? valid_85_1 : _GEN_2647; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2649 = 7'h56 == _GEN_14439 ? valid_86_1 : _GEN_2648; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2650 = 7'h57 == _GEN_14439 ? valid_87_1 : _GEN_2649; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2651 = 7'h58 == _GEN_14439 ? valid_88_1 : _GEN_2650; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2652 = 7'h59 == _GEN_14439 ? valid_89_1 : _GEN_2651; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2653 = 7'h5a == _GEN_14439 ? valid_90_1 : _GEN_2652; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2654 = 7'h5b == _GEN_14439 ? valid_91_1 : _GEN_2653; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2655 = 7'h5c == _GEN_14439 ? valid_92_1 : _GEN_2654; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2656 = 7'h5d == _GEN_14439 ? valid_93_1 : _GEN_2655; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2657 = 7'h5e == _GEN_14439 ? valid_94_1 : _GEN_2656; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2658 = 7'h5f == _GEN_14439 ? valid_95_1 : _GEN_2657; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2659 = 7'h60 == _GEN_14439 ? valid_96_1 : _GEN_2658; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2660 = 7'h61 == _GEN_14439 ? valid_97_1 : _GEN_2659; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2661 = 7'h62 == _GEN_14439 ? valid_98_1 : _GEN_2660; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2662 = 7'h63 == _GEN_14439 ? valid_99_1 : _GEN_2661; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2663 = 7'h64 == _GEN_14439 ? valid_100_1 : _GEN_2662; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2664 = 7'h65 == _GEN_14439 ? valid_101_1 : _GEN_2663; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2665 = 7'h66 == _GEN_14439 ? valid_102_1 : _GEN_2664; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2666 = 7'h67 == _GEN_14439 ? valid_103_1 : _GEN_2665; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2667 = 7'h68 == _GEN_14439 ? valid_104_1 : _GEN_2666; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2668 = 7'h69 == _GEN_14439 ? valid_105_1 : _GEN_2667; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2669 = 7'h6a == _GEN_14439 ? valid_106_1 : _GEN_2668; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2670 = 7'h6b == _GEN_14439 ? valid_107_1 : _GEN_2669; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2671 = 7'h6c == _GEN_14439 ? valid_108_1 : _GEN_2670; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2672 = 7'h6d == _GEN_14439 ? valid_109_1 : _GEN_2671; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2673 = 7'h6e == _GEN_14439 ? valid_110_1 : _GEN_2672; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2674 = 7'h6f == _GEN_14439 ? valid_111_1 : _GEN_2673; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2675 = 7'h70 == _GEN_14439 ? valid_112_1 : _GEN_2674; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2676 = 7'h71 == _GEN_14439 ? valid_113_1 : _GEN_2675; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2677 = 7'h72 == _GEN_14439 ? valid_114_1 : _GEN_2676; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2678 = 7'h73 == _GEN_14439 ? valid_115_1 : _GEN_2677; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2679 = 7'h74 == _GEN_14439 ? valid_116_1 : _GEN_2678; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2680 = 7'h75 == _GEN_14439 ? valid_117_1 : _GEN_2679; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2681 = 7'h76 == _GEN_14439 ? valid_118_1 : _GEN_2680; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2682 = 7'h77 == _GEN_14439 ? valid_119_1 : _GEN_2681; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2683 = 7'h78 == _GEN_14439 ? valid_120_1 : _GEN_2682; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2684 = 7'h79 == _GEN_14439 ? valid_121_1 : _GEN_2683; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2685 = 7'h7a == _GEN_14439 ? valid_122_1 : _GEN_2684; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2686 = 7'h7b == _GEN_14439 ? valid_123_1 : _GEN_2685; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2687 = 7'h7c == _GEN_14439 ? valid_124_1 : _GEN_2686; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2688 = 7'h7d == _GEN_14439 ? valid_125_1 : _GEN_2687; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2689 = 7'h7e == _GEN_14439 ? valid_126_1 : _GEN_2688; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2690 = 7'h7f == _GEN_14439 ? valid_127_1 : _GEN_2689; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2691 = 8'h80 == _GEN_14503 ? valid_128_1 : _GEN_2690; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2692 = 8'h81 == _GEN_14503 ? valid_129_1 : _GEN_2691; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2693 = 8'h82 == _GEN_14503 ? valid_130_1 : _GEN_2692; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2694 = 8'h83 == _GEN_14503 ? valid_131_1 : _GEN_2693; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2695 = 8'h84 == _GEN_14503 ? valid_132_1 : _GEN_2694; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2696 = 8'h85 == _GEN_14503 ? valid_133_1 : _GEN_2695; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2697 = 8'h86 == _GEN_14503 ? valid_134_1 : _GEN_2696; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2698 = 8'h87 == _GEN_14503 ? valid_135_1 : _GEN_2697; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2699 = 8'h88 == _GEN_14503 ? valid_136_1 : _GEN_2698; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2700 = 8'h89 == _GEN_14503 ? valid_137_1 : _GEN_2699; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2701 = 8'h8a == _GEN_14503 ? valid_138_1 : _GEN_2700; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2702 = 8'h8b == _GEN_14503 ? valid_139_1 : _GEN_2701; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2703 = 8'h8c == _GEN_14503 ? valid_140_1 : _GEN_2702; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2704 = 8'h8d == _GEN_14503 ? valid_141_1 : _GEN_2703; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2705 = 8'h8e == _GEN_14503 ? valid_142_1 : _GEN_2704; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2706 = 8'h8f == _GEN_14503 ? valid_143_1 : _GEN_2705; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2707 = 8'h90 == _GEN_14503 ? valid_144_1 : _GEN_2706; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2708 = 8'h91 == _GEN_14503 ? valid_145_1 : _GEN_2707; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2709 = 8'h92 == _GEN_14503 ? valid_146_1 : _GEN_2708; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2710 = 8'h93 == _GEN_14503 ? valid_147_1 : _GEN_2709; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2711 = 8'h94 == _GEN_14503 ? valid_148_1 : _GEN_2710; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2712 = 8'h95 == _GEN_14503 ? valid_149_1 : _GEN_2711; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2713 = 8'h96 == _GEN_14503 ? valid_150_1 : _GEN_2712; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2714 = 8'h97 == _GEN_14503 ? valid_151_1 : _GEN_2713; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2715 = 8'h98 == _GEN_14503 ? valid_152_1 : _GEN_2714; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2716 = 8'h99 == _GEN_14503 ? valid_153_1 : _GEN_2715; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2717 = 8'h9a == _GEN_14503 ? valid_154_1 : _GEN_2716; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2718 = 8'h9b == _GEN_14503 ? valid_155_1 : _GEN_2717; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2719 = 8'h9c == _GEN_14503 ? valid_156_1 : _GEN_2718; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2720 = 8'h9d == _GEN_14503 ? valid_157_1 : _GEN_2719; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2721 = 8'h9e == _GEN_14503 ? valid_158_1 : _GEN_2720; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2722 = 8'h9f == _GEN_14503 ? valid_159_1 : _GEN_2721; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2723 = 8'ha0 == _GEN_14503 ? valid_160_1 : _GEN_2722; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2724 = 8'ha1 == _GEN_14503 ? valid_161_1 : _GEN_2723; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2725 = 8'ha2 == _GEN_14503 ? valid_162_1 : _GEN_2724; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2726 = 8'ha3 == _GEN_14503 ? valid_163_1 : _GEN_2725; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2727 = 8'ha4 == _GEN_14503 ? valid_164_1 : _GEN_2726; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2728 = 8'ha5 == _GEN_14503 ? valid_165_1 : _GEN_2727; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2729 = 8'ha6 == _GEN_14503 ? valid_166_1 : _GEN_2728; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2730 = 8'ha7 == _GEN_14503 ? valid_167_1 : _GEN_2729; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2731 = 8'ha8 == _GEN_14503 ? valid_168_1 : _GEN_2730; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2732 = 8'ha9 == _GEN_14503 ? valid_169_1 : _GEN_2731; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2733 = 8'haa == _GEN_14503 ? valid_170_1 : _GEN_2732; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2734 = 8'hab == _GEN_14503 ? valid_171_1 : _GEN_2733; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2735 = 8'hac == _GEN_14503 ? valid_172_1 : _GEN_2734; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2736 = 8'had == _GEN_14503 ? valid_173_1 : _GEN_2735; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2737 = 8'hae == _GEN_14503 ? valid_174_1 : _GEN_2736; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2738 = 8'haf == _GEN_14503 ? valid_175_1 : _GEN_2737; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2739 = 8'hb0 == _GEN_14503 ? valid_176_1 : _GEN_2738; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2740 = 8'hb1 == _GEN_14503 ? valid_177_1 : _GEN_2739; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2741 = 8'hb2 == _GEN_14503 ? valid_178_1 : _GEN_2740; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2742 = 8'hb3 == _GEN_14503 ? valid_179_1 : _GEN_2741; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2743 = 8'hb4 == _GEN_14503 ? valid_180_1 : _GEN_2742; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2744 = 8'hb5 == _GEN_14503 ? valid_181_1 : _GEN_2743; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2745 = 8'hb6 == _GEN_14503 ? valid_182_1 : _GEN_2744; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2746 = 8'hb7 == _GEN_14503 ? valid_183_1 : _GEN_2745; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2747 = 8'hb8 == _GEN_14503 ? valid_184_1 : _GEN_2746; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2748 = 8'hb9 == _GEN_14503 ? valid_185_1 : _GEN_2747; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2749 = 8'hba == _GEN_14503 ? valid_186_1 : _GEN_2748; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2750 = 8'hbb == _GEN_14503 ? valid_187_1 : _GEN_2749; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2751 = 8'hbc == _GEN_14503 ? valid_188_1 : _GEN_2750; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2752 = 8'hbd == _GEN_14503 ? valid_189_1 : _GEN_2751; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2753 = 8'hbe == _GEN_14503 ? valid_190_1 : _GEN_2752; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2754 = 8'hbf == _GEN_14503 ? valid_191_1 : _GEN_2753; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2755 = 8'hc0 == _GEN_14503 ? valid_192_1 : _GEN_2754; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2756 = 8'hc1 == _GEN_14503 ? valid_193_1 : _GEN_2755; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2757 = 8'hc2 == _GEN_14503 ? valid_194_1 : _GEN_2756; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2758 = 8'hc3 == _GEN_14503 ? valid_195_1 : _GEN_2757; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2759 = 8'hc4 == _GEN_14503 ? valid_196_1 : _GEN_2758; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2760 = 8'hc5 == _GEN_14503 ? valid_197_1 : _GEN_2759; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2761 = 8'hc6 == _GEN_14503 ? valid_198_1 : _GEN_2760; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2762 = 8'hc7 == _GEN_14503 ? valid_199_1 : _GEN_2761; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2763 = 8'hc8 == _GEN_14503 ? valid_200_1 : _GEN_2762; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2764 = 8'hc9 == _GEN_14503 ? valid_201_1 : _GEN_2763; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2765 = 8'hca == _GEN_14503 ? valid_202_1 : _GEN_2764; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2766 = 8'hcb == _GEN_14503 ? valid_203_1 : _GEN_2765; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2767 = 8'hcc == _GEN_14503 ? valid_204_1 : _GEN_2766; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2768 = 8'hcd == _GEN_14503 ? valid_205_1 : _GEN_2767; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2769 = 8'hce == _GEN_14503 ? valid_206_1 : _GEN_2768; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2770 = 8'hcf == _GEN_14503 ? valid_207_1 : _GEN_2769; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2771 = 8'hd0 == _GEN_14503 ? valid_208_1 : _GEN_2770; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2772 = 8'hd1 == _GEN_14503 ? valid_209_1 : _GEN_2771; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2773 = 8'hd2 == _GEN_14503 ? valid_210_1 : _GEN_2772; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2774 = 8'hd3 == _GEN_14503 ? valid_211_1 : _GEN_2773; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2775 = 8'hd4 == _GEN_14503 ? valid_212_1 : _GEN_2774; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2776 = 8'hd5 == _GEN_14503 ? valid_213_1 : _GEN_2775; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2777 = 8'hd6 == _GEN_14503 ? valid_214_1 : _GEN_2776; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2778 = 8'hd7 == _GEN_14503 ? valid_215_1 : _GEN_2777; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2779 = 8'hd8 == _GEN_14503 ? valid_216_1 : _GEN_2778; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2780 = 8'hd9 == _GEN_14503 ? valid_217_1 : _GEN_2779; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2781 = 8'hda == _GEN_14503 ? valid_218_1 : _GEN_2780; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2782 = 8'hdb == _GEN_14503 ? valid_219_1 : _GEN_2781; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2783 = 8'hdc == _GEN_14503 ? valid_220_1 : _GEN_2782; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2784 = 8'hdd == _GEN_14503 ? valid_221_1 : _GEN_2783; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2785 = 8'hde == _GEN_14503 ? valid_222_1 : _GEN_2784; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2786 = 8'hdf == _GEN_14503 ? valid_223_1 : _GEN_2785; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2787 = 8'he0 == _GEN_14503 ? valid_224_1 : _GEN_2786; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2788 = 8'he1 == _GEN_14503 ? valid_225_1 : _GEN_2787; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2789 = 8'he2 == _GEN_14503 ? valid_226_1 : _GEN_2788; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2790 = 8'he3 == _GEN_14503 ? valid_227_1 : _GEN_2789; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2791 = 8'he4 == _GEN_14503 ? valid_228_1 : _GEN_2790; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2792 = 8'he5 == _GEN_14503 ? valid_229_1 : _GEN_2791; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2793 = 8'he6 == _GEN_14503 ? valid_230_1 : _GEN_2792; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2794 = 8'he7 == _GEN_14503 ? valid_231_1 : _GEN_2793; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2795 = 8'he8 == _GEN_14503 ? valid_232_1 : _GEN_2794; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2796 = 8'he9 == _GEN_14503 ? valid_233_1 : _GEN_2795; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2797 = 8'hea == _GEN_14503 ? valid_234_1 : _GEN_2796; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2798 = 8'heb == _GEN_14503 ? valid_235_1 : _GEN_2797; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2799 = 8'hec == _GEN_14503 ? valid_236_1 : _GEN_2798; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2800 = 8'hed == _GEN_14503 ? valid_237_1 : _GEN_2799; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2801 = 8'hee == _GEN_14503 ? valid_238_1 : _GEN_2800; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2802 = 8'hef == _GEN_14503 ? valid_239_1 : _GEN_2801; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2803 = 8'hf0 == _GEN_14503 ? valid_240_1 : _GEN_2802; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2804 = 8'hf1 == _GEN_14503 ? valid_241_1 : _GEN_2803; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2805 = 8'hf2 == _GEN_14503 ? valid_242_1 : _GEN_2804; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2806 = 8'hf3 == _GEN_14503 ? valid_243_1 : _GEN_2805; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2807 = 8'hf4 == _GEN_14503 ? valid_244_1 : _GEN_2806; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2808 = 8'hf5 == _GEN_14503 ? valid_245_1 : _GEN_2807; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2809 = 8'hf6 == _GEN_14503 ? valid_246_1 : _GEN_2808; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2810 = 8'hf7 == _GEN_14503 ? valid_247_1 : _GEN_2809; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2811 = 8'hf8 == _GEN_14503 ? valid_248_1 : _GEN_2810; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2812 = 8'hf9 == _GEN_14503 ? valid_249_1 : _GEN_2811; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2813 = 8'hfa == _GEN_14503 ? valid_250_1 : _GEN_2812; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2814 = 8'hfb == _GEN_14503 ? valid_251_1 : _GEN_2813; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2815 = 8'hfc == _GEN_14503 ? valid_252_1 : _GEN_2814; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2816 = 8'hfd == _GEN_14503 ? valid_253_1 : _GEN_2815; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2817 = 8'hfe == _GEN_14503 ? valid_254_1 : _GEN_2816; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2818 = 8'hff == _GEN_14503 ? valid_255_1 : _GEN_2817; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2819 = 9'h100 == _GEN_14631 ? valid_256_1 : _GEN_2818; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2820 = 9'h101 == _GEN_14631 ? valid_257_1 : _GEN_2819; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2821 = 9'h102 == _GEN_14631 ? valid_258_1 : _GEN_2820; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2822 = 9'h103 == _GEN_14631 ? valid_259_1 : _GEN_2821; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2823 = 9'h104 == _GEN_14631 ? valid_260_1 : _GEN_2822; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2824 = 9'h105 == _GEN_14631 ? valid_261_1 : _GEN_2823; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2825 = 9'h106 == _GEN_14631 ? valid_262_1 : _GEN_2824; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2826 = 9'h107 == _GEN_14631 ? valid_263_1 : _GEN_2825; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2827 = 9'h108 == _GEN_14631 ? valid_264_1 : _GEN_2826; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2828 = 9'h109 == _GEN_14631 ? valid_265_1 : _GEN_2827; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2829 = 9'h10a == _GEN_14631 ? valid_266_1 : _GEN_2828; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2830 = 9'h10b == _GEN_14631 ? valid_267_1 : _GEN_2829; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2831 = 9'h10c == _GEN_14631 ? valid_268_1 : _GEN_2830; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2832 = 9'h10d == _GEN_14631 ? valid_269_1 : _GEN_2831; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2833 = 9'h10e == _GEN_14631 ? valid_270_1 : _GEN_2832; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2834 = 9'h10f == _GEN_14631 ? valid_271_1 : _GEN_2833; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2835 = 9'h110 == _GEN_14631 ? valid_272_1 : _GEN_2834; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2836 = 9'h111 == _GEN_14631 ? valid_273_1 : _GEN_2835; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2837 = 9'h112 == _GEN_14631 ? valid_274_1 : _GEN_2836; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2838 = 9'h113 == _GEN_14631 ? valid_275_1 : _GEN_2837; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2839 = 9'h114 == _GEN_14631 ? valid_276_1 : _GEN_2838; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2840 = 9'h115 == _GEN_14631 ? valid_277_1 : _GEN_2839; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2841 = 9'h116 == _GEN_14631 ? valid_278_1 : _GEN_2840; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2842 = 9'h117 == _GEN_14631 ? valid_279_1 : _GEN_2841; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2843 = 9'h118 == _GEN_14631 ? valid_280_1 : _GEN_2842; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2844 = 9'h119 == _GEN_14631 ? valid_281_1 : _GEN_2843; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2845 = 9'h11a == _GEN_14631 ? valid_282_1 : _GEN_2844; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2846 = 9'h11b == _GEN_14631 ? valid_283_1 : _GEN_2845; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2847 = 9'h11c == _GEN_14631 ? valid_284_1 : _GEN_2846; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2848 = 9'h11d == _GEN_14631 ? valid_285_1 : _GEN_2847; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2849 = 9'h11e == _GEN_14631 ? valid_286_1 : _GEN_2848; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2850 = 9'h11f == _GEN_14631 ? valid_287_1 : _GEN_2849; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2851 = 9'h120 == _GEN_14631 ? valid_288_1 : _GEN_2850; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2852 = 9'h121 == _GEN_14631 ? valid_289_1 : _GEN_2851; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2853 = 9'h122 == _GEN_14631 ? valid_290_1 : _GEN_2852; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2854 = 9'h123 == _GEN_14631 ? valid_291_1 : _GEN_2853; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2855 = 9'h124 == _GEN_14631 ? valid_292_1 : _GEN_2854; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2856 = 9'h125 == _GEN_14631 ? valid_293_1 : _GEN_2855; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2857 = 9'h126 == _GEN_14631 ? valid_294_1 : _GEN_2856; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2858 = 9'h127 == _GEN_14631 ? valid_295_1 : _GEN_2857; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2859 = 9'h128 == _GEN_14631 ? valid_296_1 : _GEN_2858; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2860 = 9'h129 == _GEN_14631 ? valid_297_1 : _GEN_2859; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2861 = 9'h12a == _GEN_14631 ? valid_298_1 : _GEN_2860; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2862 = 9'h12b == _GEN_14631 ? valid_299_1 : _GEN_2861; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2863 = 9'h12c == _GEN_14631 ? valid_300_1 : _GEN_2862; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2864 = 9'h12d == _GEN_14631 ? valid_301_1 : _GEN_2863; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2865 = 9'h12e == _GEN_14631 ? valid_302_1 : _GEN_2864; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2866 = 9'h12f == _GEN_14631 ? valid_303_1 : _GEN_2865; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2867 = 9'h130 == _GEN_14631 ? valid_304_1 : _GEN_2866; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2868 = 9'h131 == _GEN_14631 ? valid_305_1 : _GEN_2867; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2869 = 9'h132 == _GEN_14631 ? valid_306_1 : _GEN_2868; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2870 = 9'h133 == _GEN_14631 ? valid_307_1 : _GEN_2869; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2871 = 9'h134 == _GEN_14631 ? valid_308_1 : _GEN_2870; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2872 = 9'h135 == _GEN_14631 ? valid_309_1 : _GEN_2871; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2873 = 9'h136 == _GEN_14631 ? valid_310_1 : _GEN_2872; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2874 = 9'h137 == _GEN_14631 ? valid_311_1 : _GEN_2873; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2875 = 9'h138 == _GEN_14631 ? valid_312_1 : _GEN_2874; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2876 = 9'h139 == _GEN_14631 ? valid_313_1 : _GEN_2875; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2877 = 9'h13a == _GEN_14631 ? valid_314_1 : _GEN_2876; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2878 = 9'h13b == _GEN_14631 ? valid_315_1 : _GEN_2877; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2879 = 9'h13c == _GEN_14631 ? valid_316_1 : _GEN_2878; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2880 = 9'h13d == _GEN_14631 ? valid_317_1 : _GEN_2879; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2881 = 9'h13e == _GEN_14631 ? valid_318_1 : _GEN_2880; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2882 = 9'h13f == _GEN_14631 ? valid_319_1 : _GEN_2881; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2883 = 9'h140 == _GEN_14631 ? valid_320_1 : _GEN_2882; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2884 = 9'h141 == _GEN_14631 ? valid_321_1 : _GEN_2883; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2885 = 9'h142 == _GEN_14631 ? valid_322_1 : _GEN_2884; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2886 = 9'h143 == _GEN_14631 ? valid_323_1 : _GEN_2885; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2887 = 9'h144 == _GEN_14631 ? valid_324_1 : _GEN_2886; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2888 = 9'h145 == _GEN_14631 ? valid_325_1 : _GEN_2887; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2889 = 9'h146 == _GEN_14631 ? valid_326_1 : _GEN_2888; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2890 = 9'h147 == _GEN_14631 ? valid_327_1 : _GEN_2889; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2891 = 9'h148 == _GEN_14631 ? valid_328_1 : _GEN_2890; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2892 = 9'h149 == _GEN_14631 ? valid_329_1 : _GEN_2891; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2893 = 9'h14a == _GEN_14631 ? valid_330_1 : _GEN_2892; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2894 = 9'h14b == _GEN_14631 ? valid_331_1 : _GEN_2893; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2895 = 9'h14c == _GEN_14631 ? valid_332_1 : _GEN_2894; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2896 = 9'h14d == _GEN_14631 ? valid_333_1 : _GEN_2895; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2897 = 9'h14e == _GEN_14631 ? valid_334_1 : _GEN_2896; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2898 = 9'h14f == _GEN_14631 ? valid_335_1 : _GEN_2897; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2899 = 9'h150 == _GEN_14631 ? valid_336_1 : _GEN_2898; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2900 = 9'h151 == _GEN_14631 ? valid_337_1 : _GEN_2899; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2901 = 9'h152 == _GEN_14631 ? valid_338_1 : _GEN_2900; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2902 = 9'h153 == _GEN_14631 ? valid_339_1 : _GEN_2901; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2903 = 9'h154 == _GEN_14631 ? valid_340_1 : _GEN_2902; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2904 = 9'h155 == _GEN_14631 ? valid_341_1 : _GEN_2903; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2905 = 9'h156 == _GEN_14631 ? valid_342_1 : _GEN_2904; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2906 = 9'h157 == _GEN_14631 ? valid_343_1 : _GEN_2905; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2907 = 9'h158 == _GEN_14631 ? valid_344_1 : _GEN_2906; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2908 = 9'h159 == _GEN_14631 ? valid_345_1 : _GEN_2907; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2909 = 9'h15a == _GEN_14631 ? valid_346_1 : _GEN_2908; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2910 = 9'h15b == _GEN_14631 ? valid_347_1 : _GEN_2909; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2911 = 9'h15c == _GEN_14631 ? valid_348_1 : _GEN_2910; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2912 = 9'h15d == _GEN_14631 ? valid_349_1 : _GEN_2911; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2913 = 9'h15e == _GEN_14631 ? valid_350_1 : _GEN_2912; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2914 = 9'h15f == _GEN_14631 ? valid_351_1 : _GEN_2913; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2915 = 9'h160 == _GEN_14631 ? valid_352_1 : _GEN_2914; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2916 = 9'h161 == _GEN_14631 ? valid_353_1 : _GEN_2915; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2917 = 9'h162 == _GEN_14631 ? valid_354_1 : _GEN_2916; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2918 = 9'h163 == _GEN_14631 ? valid_355_1 : _GEN_2917; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2919 = 9'h164 == _GEN_14631 ? valid_356_1 : _GEN_2918; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2920 = 9'h165 == _GEN_14631 ? valid_357_1 : _GEN_2919; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2921 = 9'h166 == _GEN_14631 ? valid_358_1 : _GEN_2920; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2922 = 9'h167 == _GEN_14631 ? valid_359_1 : _GEN_2921; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2923 = 9'h168 == _GEN_14631 ? valid_360_1 : _GEN_2922; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2924 = 9'h169 == _GEN_14631 ? valid_361_1 : _GEN_2923; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2925 = 9'h16a == _GEN_14631 ? valid_362_1 : _GEN_2924; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2926 = 9'h16b == _GEN_14631 ? valid_363_1 : _GEN_2925; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2927 = 9'h16c == _GEN_14631 ? valid_364_1 : _GEN_2926; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2928 = 9'h16d == _GEN_14631 ? valid_365_1 : _GEN_2927; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2929 = 9'h16e == _GEN_14631 ? valid_366_1 : _GEN_2928; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2930 = 9'h16f == _GEN_14631 ? valid_367_1 : _GEN_2929; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2931 = 9'h170 == _GEN_14631 ? valid_368_1 : _GEN_2930; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2932 = 9'h171 == _GEN_14631 ? valid_369_1 : _GEN_2931; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2933 = 9'h172 == _GEN_14631 ? valid_370_1 : _GEN_2932; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2934 = 9'h173 == _GEN_14631 ? valid_371_1 : _GEN_2933; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2935 = 9'h174 == _GEN_14631 ? valid_372_1 : _GEN_2934; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2936 = 9'h175 == _GEN_14631 ? valid_373_1 : _GEN_2935; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2937 = 9'h176 == _GEN_14631 ? valid_374_1 : _GEN_2936; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2938 = 9'h177 == _GEN_14631 ? valid_375_1 : _GEN_2937; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2939 = 9'h178 == _GEN_14631 ? valid_376_1 : _GEN_2938; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2940 = 9'h179 == _GEN_14631 ? valid_377_1 : _GEN_2939; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2941 = 9'h17a == _GEN_14631 ? valid_378_1 : _GEN_2940; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2942 = 9'h17b == _GEN_14631 ? valid_379_1 : _GEN_2941; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2943 = 9'h17c == _GEN_14631 ? valid_380_1 : _GEN_2942; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2944 = 9'h17d == _GEN_14631 ? valid_381_1 : _GEN_2943; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2945 = 9'h17e == _GEN_14631 ? valid_382_1 : _GEN_2944; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2946 = 9'h17f == _GEN_14631 ? valid_383_1 : _GEN_2945; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2947 = 9'h180 == _GEN_14631 ? valid_384_1 : _GEN_2946; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2948 = 9'h181 == _GEN_14631 ? valid_385_1 : _GEN_2947; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2949 = 9'h182 == _GEN_14631 ? valid_386_1 : _GEN_2948; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2950 = 9'h183 == _GEN_14631 ? valid_387_1 : _GEN_2949; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2951 = 9'h184 == _GEN_14631 ? valid_388_1 : _GEN_2950; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2952 = 9'h185 == _GEN_14631 ? valid_389_1 : _GEN_2951; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2953 = 9'h186 == _GEN_14631 ? valid_390_1 : _GEN_2952; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2954 = 9'h187 == _GEN_14631 ? valid_391_1 : _GEN_2953; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2955 = 9'h188 == _GEN_14631 ? valid_392_1 : _GEN_2954; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2956 = 9'h189 == _GEN_14631 ? valid_393_1 : _GEN_2955; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2957 = 9'h18a == _GEN_14631 ? valid_394_1 : _GEN_2956; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2958 = 9'h18b == _GEN_14631 ? valid_395_1 : _GEN_2957; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2959 = 9'h18c == _GEN_14631 ? valid_396_1 : _GEN_2958; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2960 = 9'h18d == _GEN_14631 ? valid_397_1 : _GEN_2959; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2961 = 9'h18e == _GEN_14631 ? valid_398_1 : _GEN_2960; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2962 = 9'h18f == _GEN_14631 ? valid_399_1 : _GEN_2961; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2963 = 9'h190 == _GEN_14631 ? valid_400_1 : _GEN_2962; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2964 = 9'h191 == _GEN_14631 ? valid_401_1 : _GEN_2963; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2965 = 9'h192 == _GEN_14631 ? valid_402_1 : _GEN_2964; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2966 = 9'h193 == _GEN_14631 ? valid_403_1 : _GEN_2965; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2967 = 9'h194 == _GEN_14631 ? valid_404_1 : _GEN_2966; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2968 = 9'h195 == _GEN_14631 ? valid_405_1 : _GEN_2967; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2969 = 9'h196 == _GEN_14631 ? valid_406_1 : _GEN_2968; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2970 = 9'h197 == _GEN_14631 ? valid_407_1 : _GEN_2969; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2971 = 9'h198 == _GEN_14631 ? valid_408_1 : _GEN_2970; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2972 = 9'h199 == _GEN_14631 ? valid_409_1 : _GEN_2971; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2973 = 9'h19a == _GEN_14631 ? valid_410_1 : _GEN_2972; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2974 = 9'h19b == _GEN_14631 ? valid_411_1 : _GEN_2973; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2975 = 9'h19c == _GEN_14631 ? valid_412_1 : _GEN_2974; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2976 = 9'h19d == _GEN_14631 ? valid_413_1 : _GEN_2975; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2977 = 9'h19e == _GEN_14631 ? valid_414_1 : _GEN_2976; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2978 = 9'h19f == _GEN_14631 ? valid_415_1 : _GEN_2977; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2979 = 9'h1a0 == _GEN_14631 ? valid_416_1 : _GEN_2978; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2980 = 9'h1a1 == _GEN_14631 ? valid_417_1 : _GEN_2979; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2981 = 9'h1a2 == _GEN_14631 ? valid_418_1 : _GEN_2980; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2982 = 9'h1a3 == _GEN_14631 ? valid_419_1 : _GEN_2981; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2983 = 9'h1a4 == _GEN_14631 ? valid_420_1 : _GEN_2982; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2984 = 9'h1a5 == _GEN_14631 ? valid_421_1 : _GEN_2983; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2985 = 9'h1a6 == _GEN_14631 ? valid_422_1 : _GEN_2984; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2986 = 9'h1a7 == _GEN_14631 ? valid_423_1 : _GEN_2985; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2987 = 9'h1a8 == _GEN_14631 ? valid_424_1 : _GEN_2986; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2988 = 9'h1a9 == _GEN_14631 ? valid_425_1 : _GEN_2987; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2989 = 9'h1aa == _GEN_14631 ? valid_426_1 : _GEN_2988; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2990 = 9'h1ab == _GEN_14631 ? valid_427_1 : _GEN_2989; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2991 = 9'h1ac == _GEN_14631 ? valid_428_1 : _GEN_2990; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2992 = 9'h1ad == _GEN_14631 ? valid_429_1 : _GEN_2991; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2993 = 9'h1ae == _GEN_14631 ? valid_430_1 : _GEN_2992; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2994 = 9'h1af == _GEN_14631 ? valid_431_1 : _GEN_2993; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2995 = 9'h1b0 == _GEN_14631 ? valid_432_1 : _GEN_2994; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2996 = 9'h1b1 == _GEN_14631 ? valid_433_1 : _GEN_2995; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2997 = 9'h1b2 == _GEN_14631 ? valid_434_1 : _GEN_2996; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2998 = 9'h1b3 == _GEN_14631 ? valid_435_1 : _GEN_2997; // @[ICache.scala 101:{81,81}]
  wire  _GEN_2999 = 9'h1b4 == _GEN_14631 ? valid_436_1 : _GEN_2998; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3000 = 9'h1b5 == _GEN_14631 ? valid_437_1 : _GEN_2999; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3001 = 9'h1b6 == _GEN_14631 ? valid_438_1 : _GEN_3000; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3002 = 9'h1b7 == _GEN_14631 ? valid_439_1 : _GEN_3001; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3003 = 9'h1b8 == _GEN_14631 ? valid_440_1 : _GEN_3002; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3004 = 9'h1b9 == _GEN_14631 ? valid_441_1 : _GEN_3003; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3005 = 9'h1ba == _GEN_14631 ? valid_442_1 : _GEN_3004; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3006 = 9'h1bb == _GEN_14631 ? valid_443_1 : _GEN_3005; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3007 = 9'h1bc == _GEN_14631 ? valid_444_1 : _GEN_3006; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3008 = 9'h1bd == _GEN_14631 ? valid_445_1 : _GEN_3007; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3009 = 9'h1be == _GEN_14631 ? valid_446_1 : _GEN_3008; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3010 = 9'h1bf == _GEN_14631 ? valid_447_1 : _GEN_3009; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3011 = 9'h1c0 == _GEN_14631 ? valid_448_1 : _GEN_3010; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3012 = 9'h1c1 == _GEN_14631 ? valid_449_1 : _GEN_3011; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3013 = 9'h1c2 == _GEN_14631 ? valid_450_1 : _GEN_3012; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3014 = 9'h1c3 == _GEN_14631 ? valid_451_1 : _GEN_3013; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3015 = 9'h1c4 == _GEN_14631 ? valid_452_1 : _GEN_3014; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3016 = 9'h1c5 == _GEN_14631 ? valid_453_1 : _GEN_3015; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3017 = 9'h1c6 == _GEN_14631 ? valid_454_1 : _GEN_3016; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3018 = 9'h1c7 == _GEN_14631 ? valid_455_1 : _GEN_3017; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3019 = 9'h1c8 == _GEN_14631 ? valid_456_1 : _GEN_3018; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3020 = 9'h1c9 == _GEN_14631 ? valid_457_1 : _GEN_3019; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3021 = 9'h1ca == _GEN_14631 ? valid_458_1 : _GEN_3020; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3022 = 9'h1cb == _GEN_14631 ? valid_459_1 : _GEN_3021; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3023 = 9'h1cc == _GEN_14631 ? valid_460_1 : _GEN_3022; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3024 = 9'h1cd == _GEN_14631 ? valid_461_1 : _GEN_3023; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3025 = 9'h1ce == _GEN_14631 ? valid_462_1 : _GEN_3024; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3026 = 9'h1cf == _GEN_14631 ? valid_463_1 : _GEN_3025; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3027 = 9'h1d0 == _GEN_14631 ? valid_464_1 : _GEN_3026; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3028 = 9'h1d1 == _GEN_14631 ? valid_465_1 : _GEN_3027; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3029 = 9'h1d2 == _GEN_14631 ? valid_466_1 : _GEN_3028; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3030 = 9'h1d3 == _GEN_14631 ? valid_467_1 : _GEN_3029; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3031 = 9'h1d4 == _GEN_14631 ? valid_468_1 : _GEN_3030; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3032 = 9'h1d5 == _GEN_14631 ? valid_469_1 : _GEN_3031; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3033 = 9'h1d6 == _GEN_14631 ? valid_470_1 : _GEN_3032; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3034 = 9'h1d7 == _GEN_14631 ? valid_471_1 : _GEN_3033; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3035 = 9'h1d8 == _GEN_14631 ? valid_472_1 : _GEN_3034; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3036 = 9'h1d9 == _GEN_14631 ? valid_473_1 : _GEN_3035; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3037 = 9'h1da == _GEN_14631 ? valid_474_1 : _GEN_3036; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3038 = 9'h1db == _GEN_14631 ? valid_475_1 : _GEN_3037; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3039 = 9'h1dc == _GEN_14631 ? valid_476_1 : _GEN_3038; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3040 = 9'h1dd == _GEN_14631 ? valid_477_1 : _GEN_3039; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3041 = 9'h1de == _GEN_14631 ? valid_478_1 : _GEN_3040; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3042 = 9'h1df == _GEN_14631 ? valid_479_1 : _GEN_3041; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3043 = 9'h1e0 == _GEN_14631 ? valid_480_1 : _GEN_3042; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3044 = 9'h1e1 == _GEN_14631 ? valid_481_1 : _GEN_3043; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3045 = 9'h1e2 == _GEN_14631 ? valid_482_1 : _GEN_3044; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3046 = 9'h1e3 == _GEN_14631 ? valid_483_1 : _GEN_3045; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3047 = 9'h1e4 == _GEN_14631 ? valid_484_1 : _GEN_3046; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3048 = 9'h1e5 == _GEN_14631 ? valid_485_1 : _GEN_3047; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3049 = 9'h1e6 == _GEN_14631 ? valid_486_1 : _GEN_3048; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3050 = 9'h1e7 == _GEN_14631 ? valid_487_1 : _GEN_3049; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3051 = 9'h1e8 == _GEN_14631 ? valid_488_1 : _GEN_3050; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3052 = 9'h1e9 == _GEN_14631 ? valid_489_1 : _GEN_3051; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3053 = 9'h1ea == _GEN_14631 ? valid_490_1 : _GEN_3052; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3054 = 9'h1eb == _GEN_14631 ? valid_491_1 : _GEN_3053; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3055 = 9'h1ec == _GEN_14631 ? valid_492_1 : _GEN_3054; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3056 = 9'h1ed == _GEN_14631 ? valid_493_1 : _GEN_3055; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3057 = 9'h1ee == _GEN_14631 ? valid_494_1 : _GEN_3056; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3058 = 9'h1ef == _GEN_14631 ? valid_495_1 : _GEN_3057; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3059 = 9'h1f0 == _GEN_14631 ? valid_496_1 : _GEN_3058; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3060 = 9'h1f1 == _GEN_14631 ? valid_497_1 : _GEN_3059; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3061 = 9'h1f2 == _GEN_14631 ? valid_498_1 : _GEN_3060; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3062 = 9'h1f3 == _GEN_14631 ? valid_499_1 : _GEN_3061; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3063 = 9'h1f4 == _GEN_14631 ? valid_500_1 : _GEN_3062; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3064 = 9'h1f5 == _GEN_14631 ? valid_501_1 : _GEN_3063; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3065 = 9'h1f6 == _GEN_14631 ? valid_502_1 : _GEN_3064; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3066 = 9'h1f7 == _GEN_14631 ? valid_503_1 : _GEN_3065; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3067 = 9'h1f8 == _GEN_14631 ? valid_504_1 : _GEN_3066; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3068 = 9'h1f9 == _GEN_14631 ? valid_505_1 : _GEN_3067; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3069 = 9'h1fa == _GEN_14631 ? valid_506_1 : _GEN_3068; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3070 = 9'h1fb == _GEN_14631 ? valid_507_1 : _GEN_3069; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3071 = 9'h1fc == _GEN_14631 ? valid_508_1 : _GEN_3070; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3072 = 9'h1fd == _GEN_14631 ? valid_509_1 : _GEN_3071; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3073 = 9'h1fe == _GEN_14631 ? valid_510_1 : _GEN_3072; // @[ICache.scala 101:{81,81}]
  wire  _GEN_3074 = 9'h1ff == _GEN_14631 ? valid_511_1 : _GEN_3073; // @[ICache.scala 101:{81,81}]
  wire  tag_compare_valid_1 = tag_1 == inst_tag & _GEN_3074; // @[ICache.scala 101:81]
  wire  cache_hit = tag_compare_valid_0 | tag_compare_valid_1; // @[ICache.scala 102:55]
  wire  cache_hit_available = cache_hit & translation_ok & ~uncached; // @[ICache.scala 103:57]
  wire  inst_valid_1 = cache_hit_available & ~io_cpu_addr_0[2]; // @[ICache.scala 107:40]
  wire [31:0] data_0_1 = bank_1_io_rdata; // @[ICache.scala 54:18 125:19]
  wire [31:0] data_1_1 = bank_3_io_rdata; // @[ICache.scala 54:18 125:19]
  wire [31:0] inst_1 = tag_compare_valid_1 ? data_1_1 : data_0_1; // @[ICache.scala 111:{49,49}]
  wire [31:0] data_0_0 = bank_io_rdata; // @[ICache.scala 54:18 125:19]
  wire [31:0] data_1_0 = bank_2_io_rdata; // @[ICache.scala 54:18 125:19]
  wire [31:0] _GEN_3078 = tag_compare_valid_1 ? data_1_0 : data_0_0; // @[ICache.scala 111:{49,49}]
  wire [31:0] inst_0 = io_cpu_addr_0[2] ? inst_1 : _GEN_3078; // @[ICache.scala 111:49]
  reg [31:0] saved_0_inst; // @[ICache.scala 113:22]
  reg  saved_0_valid; // @[ICache.scala 113:22]
  reg [31:0] saved_1_inst; // @[ICache.scala 113:22]
  reg  saved_1_valid; // @[ICache.scala 113:22]
  reg [4:0] axi_cnt_value; // @[Counter.scala 61:40]
  wire  _io_cpu_inst_valid_0_T_4 = _should_next_addr_T ? cache_hit_available : saved_0_valid; // @[ICache.scala 142:32]
  wire  _io_cpu_inst_valid_1_T_4 = _should_next_addr_T ? inst_valid_1 : saved_1_valid; // @[ICache.scala 142:32]
  reg [31:0] ar_addr; // @[ICache.scala 149:24]
  reg [7:0] ar_len; // @[ICache.scala 149:24]
  reg [2:0] ar_size; // @[ICache.scala 149:24]
  reg  arvalid; // @[ICache.scala 150:24]
  reg  rready; // @[ICache.scala 155:23]
  reg  tlb1_invalid; // @[ICache.scala 159:29]
  wire  _io_cpu_tlb2_vpn_T_2 = ~translation_ok; // @[ICache.scala 162:76]
  wire  _io_cpu_tlb2_vpn_T_3 = _should_next_addr_T & io_cpu_req & ~translation_ok; // @[ICache.scala 162:73]
  reg [19:0] io_cpu_tlb2_vpn_r; // @[Reg.scala 19:16]
  wire [31:0] _ar_addr_T_1 = {inst_pa[31:6],6'h0}; // @[Cat.scala 33:92]
  wire  _GEN_3081 = 6'h1 == vset ? lru_1 : lru_0; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3082 = 6'h2 == vset ? lru_2 : _GEN_3081; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3083 = 6'h3 == vset ? lru_3 : _GEN_3082; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3084 = 6'h4 == vset ? lru_4 : _GEN_3083; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3085 = 6'h5 == vset ? lru_5 : _GEN_3084; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3086 = 6'h6 == vset ? lru_6 : _GEN_3085; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3087 = 6'h7 == vset ? lru_7 : _GEN_3086; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3088 = 6'h8 == vset ? lru_8 : _GEN_3087; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3089 = 6'h9 == vset ? lru_9 : _GEN_3088; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3090 = 6'ha == vset ? lru_10 : _GEN_3089; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3091 = 6'hb == vset ? lru_11 : _GEN_3090; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3092 = 6'hc == vset ? lru_12 : _GEN_3091; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3093 = 6'hd == vset ? lru_13 : _GEN_3092; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3094 = 6'he == vset ? lru_14 : _GEN_3093; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3095 = 6'hf == vset ? lru_15 : _GEN_3094; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3096 = 6'h10 == vset ? lru_16 : _GEN_3095; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3097 = 6'h11 == vset ? lru_17 : _GEN_3096; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3098 = 6'h12 == vset ? lru_18 : _GEN_3097; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3099 = 6'h13 == vset ? lru_19 : _GEN_3098; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3100 = 6'h14 == vset ? lru_20 : _GEN_3099; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3101 = 6'h15 == vset ? lru_21 : _GEN_3100; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3102 = 6'h16 == vset ? lru_22 : _GEN_3101; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3103 = 6'h17 == vset ? lru_23 : _GEN_3102; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3104 = 6'h18 == vset ? lru_24 : _GEN_3103; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3105 = 6'h19 == vset ? lru_25 : _GEN_3104; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3106 = 6'h1a == vset ? lru_26 : _GEN_3105; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3107 = 6'h1b == vset ? lru_27 : _GEN_3106; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3108 = 6'h1c == vset ? lru_28 : _GEN_3107; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3109 = 6'h1d == vset ? lru_29 : _GEN_3108; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3110 = 6'h1e == vset ? lru_30 : _GEN_3109; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3111 = 6'h1f == vset ? lru_31 : _GEN_3110; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3112 = 6'h20 == vset ? lru_32 : _GEN_3111; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3113 = 6'h21 == vset ? lru_33 : _GEN_3112; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3114 = 6'h22 == vset ? lru_34 : _GEN_3113; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3115 = 6'h23 == vset ? lru_35 : _GEN_3114; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3116 = 6'h24 == vset ? lru_36 : _GEN_3115; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3117 = 6'h25 == vset ? lru_37 : _GEN_3116; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3118 = 6'h26 == vset ? lru_38 : _GEN_3117; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3119 = 6'h27 == vset ? lru_39 : _GEN_3118; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3120 = 6'h28 == vset ? lru_40 : _GEN_3119; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3121 = 6'h29 == vset ? lru_41 : _GEN_3120; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3122 = 6'h2a == vset ? lru_42 : _GEN_3121; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3123 = 6'h2b == vset ? lru_43 : _GEN_3122; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3124 = 6'h2c == vset ? lru_44 : _GEN_3123; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3125 = 6'h2d == vset ? lru_45 : _GEN_3124; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3126 = 6'h2e == vset ? lru_46 : _GEN_3125; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3127 = 6'h2f == vset ? lru_47 : _GEN_3126; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3128 = 6'h30 == vset ? lru_48 : _GEN_3127; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3129 = 6'h31 == vset ? lru_49 : _GEN_3128; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3130 = 6'h32 == vset ? lru_50 : _GEN_3129; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3131 = 6'h33 == vset ? lru_51 : _GEN_3130; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3132 = 6'h34 == vset ? lru_52 : _GEN_3131; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3133 = 6'h35 == vset ? lru_53 : _GEN_3132; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3134 = 6'h36 == vset ? lru_54 : _GEN_3133; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3135 = 6'h37 == vset ? lru_55 : _GEN_3134; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3136 = 6'h38 == vset ? lru_56 : _GEN_3135; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3137 = 6'h39 == vset ? lru_57 : _GEN_3136; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3138 = 6'h3a == vset ? lru_58 : _GEN_3137; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3139 = 6'h3b == vset ? lru_59 : _GEN_3138; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3140 = 6'h3c == vset ? lru_60 : _GEN_3139; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3141 = 6'h3d == vset ? lru_61 : _GEN_3140; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3142 = 6'h3e == vset ? lru_62 : _GEN_3141; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3143 = 6'h3f == vset ? lru_63 : _GEN_3142; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3144 = 7'h40 == _GEN_14439 ? lru_64 : _GEN_3143; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3145 = 7'h41 == _GEN_14439 ? lru_65 : _GEN_3144; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3146 = 7'h42 == _GEN_14439 ? lru_66 : _GEN_3145; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3147 = 7'h43 == _GEN_14439 ? lru_67 : _GEN_3146; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3148 = 7'h44 == _GEN_14439 ? lru_68 : _GEN_3147; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3149 = 7'h45 == _GEN_14439 ? lru_69 : _GEN_3148; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3150 = 7'h46 == _GEN_14439 ? lru_70 : _GEN_3149; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3151 = 7'h47 == _GEN_14439 ? lru_71 : _GEN_3150; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3152 = 7'h48 == _GEN_14439 ? lru_72 : _GEN_3151; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3153 = 7'h49 == _GEN_14439 ? lru_73 : _GEN_3152; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3154 = 7'h4a == _GEN_14439 ? lru_74 : _GEN_3153; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3155 = 7'h4b == _GEN_14439 ? lru_75 : _GEN_3154; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3156 = 7'h4c == _GEN_14439 ? lru_76 : _GEN_3155; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3157 = 7'h4d == _GEN_14439 ? lru_77 : _GEN_3156; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3158 = 7'h4e == _GEN_14439 ? lru_78 : _GEN_3157; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3159 = 7'h4f == _GEN_14439 ? lru_79 : _GEN_3158; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3160 = 7'h50 == _GEN_14439 ? lru_80 : _GEN_3159; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3161 = 7'h51 == _GEN_14439 ? lru_81 : _GEN_3160; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3162 = 7'h52 == _GEN_14439 ? lru_82 : _GEN_3161; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3163 = 7'h53 == _GEN_14439 ? lru_83 : _GEN_3162; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3164 = 7'h54 == _GEN_14439 ? lru_84 : _GEN_3163; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3165 = 7'h55 == _GEN_14439 ? lru_85 : _GEN_3164; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3166 = 7'h56 == _GEN_14439 ? lru_86 : _GEN_3165; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3167 = 7'h57 == _GEN_14439 ? lru_87 : _GEN_3166; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3168 = 7'h58 == _GEN_14439 ? lru_88 : _GEN_3167; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3169 = 7'h59 == _GEN_14439 ? lru_89 : _GEN_3168; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3170 = 7'h5a == _GEN_14439 ? lru_90 : _GEN_3169; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3171 = 7'h5b == _GEN_14439 ? lru_91 : _GEN_3170; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3172 = 7'h5c == _GEN_14439 ? lru_92 : _GEN_3171; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3173 = 7'h5d == _GEN_14439 ? lru_93 : _GEN_3172; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3174 = 7'h5e == _GEN_14439 ? lru_94 : _GEN_3173; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3175 = 7'h5f == _GEN_14439 ? lru_95 : _GEN_3174; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3176 = 7'h60 == _GEN_14439 ? lru_96 : _GEN_3175; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3177 = 7'h61 == _GEN_14439 ? lru_97 : _GEN_3176; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3178 = 7'h62 == _GEN_14439 ? lru_98 : _GEN_3177; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3179 = 7'h63 == _GEN_14439 ? lru_99 : _GEN_3178; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3180 = 7'h64 == _GEN_14439 ? lru_100 : _GEN_3179; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3181 = 7'h65 == _GEN_14439 ? lru_101 : _GEN_3180; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3182 = 7'h66 == _GEN_14439 ? lru_102 : _GEN_3181; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3183 = 7'h67 == _GEN_14439 ? lru_103 : _GEN_3182; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3184 = 7'h68 == _GEN_14439 ? lru_104 : _GEN_3183; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3185 = 7'h69 == _GEN_14439 ? lru_105 : _GEN_3184; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3186 = 7'h6a == _GEN_14439 ? lru_106 : _GEN_3185; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3187 = 7'h6b == _GEN_14439 ? lru_107 : _GEN_3186; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3188 = 7'h6c == _GEN_14439 ? lru_108 : _GEN_3187; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3189 = 7'h6d == _GEN_14439 ? lru_109 : _GEN_3188; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3190 = 7'h6e == _GEN_14439 ? lru_110 : _GEN_3189; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3191 = 7'h6f == _GEN_14439 ? lru_111 : _GEN_3190; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3192 = 7'h70 == _GEN_14439 ? lru_112 : _GEN_3191; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3193 = 7'h71 == _GEN_14439 ? lru_113 : _GEN_3192; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3194 = 7'h72 == _GEN_14439 ? lru_114 : _GEN_3193; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3195 = 7'h73 == _GEN_14439 ? lru_115 : _GEN_3194; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3196 = 7'h74 == _GEN_14439 ? lru_116 : _GEN_3195; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3197 = 7'h75 == _GEN_14439 ? lru_117 : _GEN_3196; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3198 = 7'h76 == _GEN_14439 ? lru_118 : _GEN_3197; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3199 = 7'h77 == _GEN_14439 ? lru_119 : _GEN_3198; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3200 = 7'h78 == _GEN_14439 ? lru_120 : _GEN_3199; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3201 = 7'h79 == _GEN_14439 ? lru_121 : _GEN_3200; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3202 = 7'h7a == _GEN_14439 ? lru_122 : _GEN_3201; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3203 = 7'h7b == _GEN_14439 ? lru_123 : _GEN_3202; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3204 = 7'h7c == _GEN_14439 ? lru_124 : _GEN_3203; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3205 = 7'h7d == _GEN_14439 ? lru_125 : _GEN_3204; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3206 = 7'h7e == _GEN_14439 ? lru_126 : _GEN_3205; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3207 = 7'h7f == _GEN_14439 ? lru_127 : _GEN_3206; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3208 = 8'h80 == _GEN_14503 ? lru_128 : _GEN_3207; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3209 = 8'h81 == _GEN_14503 ? lru_129 : _GEN_3208; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3210 = 8'h82 == _GEN_14503 ? lru_130 : _GEN_3209; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3211 = 8'h83 == _GEN_14503 ? lru_131 : _GEN_3210; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3212 = 8'h84 == _GEN_14503 ? lru_132 : _GEN_3211; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3213 = 8'h85 == _GEN_14503 ? lru_133 : _GEN_3212; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3214 = 8'h86 == _GEN_14503 ? lru_134 : _GEN_3213; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3215 = 8'h87 == _GEN_14503 ? lru_135 : _GEN_3214; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3216 = 8'h88 == _GEN_14503 ? lru_136 : _GEN_3215; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3217 = 8'h89 == _GEN_14503 ? lru_137 : _GEN_3216; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3218 = 8'h8a == _GEN_14503 ? lru_138 : _GEN_3217; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3219 = 8'h8b == _GEN_14503 ? lru_139 : _GEN_3218; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3220 = 8'h8c == _GEN_14503 ? lru_140 : _GEN_3219; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3221 = 8'h8d == _GEN_14503 ? lru_141 : _GEN_3220; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3222 = 8'h8e == _GEN_14503 ? lru_142 : _GEN_3221; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3223 = 8'h8f == _GEN_14503 ? lru_143 : _GEN_3222; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3224 = 8'h90 == _GEN_14503 ? lru_144 : _GEN_3223; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3225 = 8'h91 == _GEN_14503 ? lru_145 : _GEN_3224; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3226 = 8'h92 == _GEN_14503 ? lru_146 : _GEN_3225; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3227 = 8'h93 == _GEN_14503 ? lru_147 : _GEN_3226; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3228 = 8'h94 == _GEN_14503 ? lru_148 : _GEN_3227; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3229 = 8'h95 == _GEN_14503 ? lru_149 : _GEN_3228; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3230 = 8'h96 == _GEN_14503 ? lru_150 : _GEN_3229; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3231 = 8'h97 == _GEN_14503 ? lru_151 : _GEN_3230; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3232 = 8'h98 == _GEN_14503 ? lru_152 : _GEN_3231; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3233 = 8'h99 == _GEN_14503 ? lru_153 : _GEN_3232; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3234 = 8'h9a == _GEN_14503 ? lru_154 : _GEN_3233; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3235 = 8'h9b == _GEN_14503 ? lru_155 : _GEN_3234; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3236 = 8'h9c == _GEN_14503 ? lru_156 : _GEN_3235; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3237 = 8'h9d == _GEN_14503 ? lru_157 : _GEN_3236; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3238 = 8'h9e == _GEN_14503 ? lru_158 : _GEN_3237; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3239 = 8'h9f == _GEN_14503 ? lru_159 : _GEN_3238; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3240 = 8'ha0 == _GEN_14503 ? lru_160 : _GEN_3239; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3241 = 8'ha1 == _GEN_14503 ? lru_161 : _GEN_3240; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3242 = 8'ha2 == _GEN_14503 ? lru_162 : _GEN_3241; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3243 = 8'ha3 == _GEN_14503 ? lru_163 : _GEN_3242; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3244 = 8'ha4 == _GEN_14503 ? lru_164 : _GEN_3243; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3245 = 8'ha5 == _GEN_14503 ? lru_165 : _GEN_3244; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3246 = 8'ha6 == _GEN_14503 ? lru_166 : _GEN_3245; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3247 = 8'ha7 == _GEN_14503 ? lru_167 : _GEN_3246; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3248 = 8'ha8 == _GEN_14503 ? lru_168 : _GEN_3247; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3249 = 8'ha9 == _GEN_14503 ? lru_169 : _GEN_3248; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3250 = 8'haa == _GEN_14503 ? lru_170 : _GEN_3249; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3251 = 8'hab == _GEN_14503 ? lru_171 : _GEN_3250; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3252 = 8'hac == _GEN_14503 ? lru_172 : _GEN_3251; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3253 = 8'had == _GEN_14503 ? lru_173 : _GEN_3252; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3254 = 8'hae == _GEN_14503 ? lru_174 : _GEN_3253; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3255 = 8'haf == _GEN_14503 ? lru_175 : _GEN_3254; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3256 = 8'hb0 == _GEN_14503 ? lru_176 : _GEN_3255; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3257 = 8'hb1 == _GEN_14503 ? lru_177 : _GEN_3256; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3258 = 8'hb2 == _GEN_14503 ? lru_178 : _GEN_3257; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3259 = 8'hb3 == _GEN_14503 ? lru_179 : _GEN_3258; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3260 = 8'hb4 == _GEN_14503 ? lru_180 : _GEN_3259; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3261 = 8'hb5 == _GEN_14503 ? lru_181 : _GEN_3260; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3262 = 8'hb6 == _GEN_14503 ? lru_182 : _GEN_3261; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3263 = 8'hb7 == _GEN_14503 ? lru_183 : _GEN_3262; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3264 = 8'hb8 == _GEN_14503 ? lru_184 : _GEN_3263; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3265 = 8'hb9 == _GEN_14503 ? lru_185 : _GEN_3264; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3266 = 8'hba == _GEN_14503 ? lru_186 : _GEN_3265; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3267 = 8'hbb == _GEN_14503 ? lru_187 : _GEN_3266; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3268 = 8'hbc == _GEN_14503 ? lru_188 : _GEN_3267; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3269 = 8'hbd == _GEN_14503 ? lru_189 : _GEN_3268; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3270 = 8'hbe == _GEN_14503 ? lru_190 : _GEN_3269; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3271 = 8'hbf == _GEN_14503 ? lru_191 : _GEN_3270; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3272 = 8'hc0 == _GEN_14503 ? lru_192 : _GEN_3271; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3273 = 8'hc1 == _GEN_14503 ? lru_193 : _GEN_3272; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3274 = 8'hc2 == _GEN_14503 ? lru_194 : _GEN_3273; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3275 = 8'hc3 == _GEN_14503 ? lru_195 : _GEN_3274; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3276 = 8'hc4 == _GEN_14503 ? lru_196 : _GEN_3275; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3277 = 8'hc5 == _GEN_14503 ? lru_197 : _GEN_3276; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3278 = 8'hc6 == _GEN_14503 ? lru_198 : _GEN_3277; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3279 = 8'hc7 == _GEN_14503 ? lru_199 : _GEN_3278; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3280 = 8'hc8 == _GEN_14503 ? lru_200 : _GEN_3279; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3281 = 8'hc9 == _GEN_14503 ? lru_201 : _GEN_3280; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3282 = 8'hca == _GEN_14503 ? lru_202 : _GEN_3281; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3283 = 8'hcb == _GEN_14503 ? lru_203 : _GEN_3282; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3284 = 8'hcc == _GEN_14503 ? lru_204 : _GEN_3283; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3285 = 8'hcd == _GEN_14503 ? lru_205 : _GEN_3284; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3286 = 8'hce == _GEN_14503 ? lru_206 : _GEN_3285; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3287 = 8'hcf == _GEN_14503 ? lru_207 : _GEN_3286; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3288 = 8'hd0 == _GEN_14503 ? lru_208 : _GEN_3287; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3289 = 8'hd1 == _GEN_14503 ? lru_209 : _GEN_3288; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3290 = 8'hd2 == _GEN_14503 ? lru_210 : _GEN_3289; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3291 = 8'hd3 == _GEN_14503 ? lru_211 : _GEN_3290; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3292 = 8'hd4 == _GEN_14503 ? lru_212 : _GEN_3291; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3293 = 8'hd5 == _GEN_14503 ? lru_213 : _GEN_3292; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3294 = 8'hd6 == _GEN_14503 ? lru_214 : _GEN_3293; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3295 = 8'hd7 == _GEN_14503 ? lru_215 : _GEN_3294; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3296 = 8'hd8 == _GEN_14503 ? lru_216 : _GEN_3295; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3297 = 8'hd9 == _GEN_14503 ? lru_217 : _GEN_3296; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3298 = 8'hda == _GEN_14503 ? lru_218 : _GEN_3297; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3299 = 8'hdb == _GEN_14503 ? lru_219 : _GEN_3298; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3300 = 8'hdc == _GEN_14503 ? lru_220 : _GEN_3299; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3301 = 8'hdd == _GEN_14503 ? lru_221 : _GEN_3300; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3302 = 8'hde == _GEN_14503 ? lru_222 : _GEN_3301; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3303 = 8'hdf == _GEN_14503 ? lru_223 : _GEN_3302; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3304 = 8'he0 == _GEN_14503 ? lru_224 : _GEN_3303; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3305 = 8'he1 == _GEN_14503 ? lru_225 : _GEN_3304; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3306 = 8'he2 == _GEN_14503 ? lru_226 : _GEN_3305; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3307 = 8'he3 == _GEN_14503 ? lru_227 : _GEN_3306; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3308 = 8'he4 == _GEN_14503 ? lru_228 : _GEN_3307; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3309 = 8'he5 == _GEN_14503 ? lru_229 : _GEN_3308; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3310 = 8'he6 == _GEN_14503 ? lru_230 : _GEN_3309; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3311 = 8'he7 == _GEN_14503 ? lru_231 : _GEN_3310; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3312 = 8'he8 == _GEN_14503 ? lru_232 : _GEN_3311; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3313 = 8'he9 == _GEN_14503 ? lru_233 : _GEN_3312; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3314 = 8'hea == _GEN_14503 ? lru_234 : _GEN_3313; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3315 = 8'heb == _GEN_14503 ? lru_235 : _GEN_3314; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3316 = 8'hec == _GEN_14503 ? lru_236 : _GEN_3315; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3317 = 8'hed == _GEN_14503 ? lru_237 : _GEN_3316; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3318 = 8'hee == _GEN_14503 ? lru_238 : _GEN_3317; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3319 = 8'hef == _GEN_14503 ? lru_239 : _GEN_3318; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3320 = 8'hf0 == _GEN_14503 ? lru_240 : _GEN_3319; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3321 = 8'hf1 == _GEN_14503 ? lru_241 : _GEN_3320; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3322 = 8'hf2 == _GEN_14503 ? lru_242 : _GEN_3321; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3323 = 8'hf3 == _GEN_14503 ? lru_243 : _GEN_3322; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3324 = 8'hf4 == _GEN_14503 ? lru_244 : _GEN_3323; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3325 = 8'hf5 == _GEN_14503 ? lru_245 : _GEN_3324; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3326 = 8'hf6 == _GEN_14503 ? lru_246 : _GEN_3325; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3327 = 8'hf7 == _GEN_14503 ? lru_247 : _GEN_3326; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3328 = 8'hf8 == _GEN_14503 ? lru_248 : _GEN_3327; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3329 = 8'hf9 == _GEN_14503 ? lru_249 : _GEN_3328; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3330 = 8'hfa == _GEN_14503 ? lru_250 : _GEN_3329; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3331 = 8'hfb == _GEN_14503 ? lru_251 : _GEN_3330; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3332 = 8'hfc == _GEN_14503 ? lru_252 : _GEN_3331; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3333 = 8'hfd == _GEN_14503 ? lru_253 : _GEN_3332; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3334 = 8'hfe == _GEN_14503 ? lru_254 : _GEN_3333; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3335 = 8'hff == _GEN_14503 ? lru_255 : _GEN_3334; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3336 = 9'h100 == _GEN_14631 ? lru_256 : _GEN_3335; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3337 = 9'h101 == _GEN_14631 ? lru_257 : _GEN_3336; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3338 = 9'h102 == _GEN_14631 ? lru_258 : _GEN_3337; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3339 = 9'h103 == _GEN_14631 ? lru_259 : _GEN_3338; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3340 = 9'h104 == _GEN_14631 ? lru_260 : _GEN_3339; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3341 = 9'h105 == _GEN_14631 ? lru_261 : _GEN_3340; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3342 = 9'h106 == _GEN_14631 ? lru_262 : _GEN_3341; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3343 = 9'h107 == _GEN_14631 ? lru_263 : _GEN_3342; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3344 = 9'h108 == _GEN_14631 ? lru_264 : _GEN_3343; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3345 = 9'h109 == _GEN_14631 ? lru_265 : _GEN_3344; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3346 = 9'h10a == _GEN_14631 ? lru_266 : _GEN_3345; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3347 = 9'h10b == _GEN_14631 ? lru_267 : _GEN_3346; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3348 = 9'h10c == _GEN_14631 ? lru_268 : _GEN_3347; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3349 = 9'h10d == _GEN_14631 ? lru_269 : _GEN_3348; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3350 = 9'h10e == _GEN_14631 ? lru_270 : _GEN_3349; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3351 = 9'h10f == _GEN_14631 ? lru_271 : _GEN_3350; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3352 = 9'h110 == _GEN_14631 ? lru_272 : _GEN_3351; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3353 = 9'h111 == _GEN_14631 ? lru_273 : _GEN_3352; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3354 = 9'h112 == _GEN_14631 ? lru_274 : _GEN_3353; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3355 = 9'h113 == _GEN_14631 ? lru_275 : _GEN_3354; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3356 = 9'h114 == _GEN_14631 ? lru_276 : _GEN_3355; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3357 = 9'h115 == _GEN_14631 ? lru_277 : _GEN_3356; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3358 = 9'h116 == _GEN_14631 ? lru_278 : _GEN_3357; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3359 = 9'h117 == _GEN_14631 ? lru_279 : _GEN_3358; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3360 = 9'h118 == _GEN_14631 ? lru_280 : _GEN_3359; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3361 = 9'h119 == _GEN_14631 ? lru_281 : _GEN_3360; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3362 = 9'h11a == _GEN_14631 ? lru_282 : _GEN_3361; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3363 = 9'h11b == _GEN_14631 ? lru_283 : _GEN_3362; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3364 = 9'h11c == _GEN_14631 ? lru_284 : _GEN_3363; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3365 = 9'h11d == _GEN_14631 ? lru_285 : _GEN_3364; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3366 = 9'h11e == _GEN_14631 ? lru_286 : _GEN_3365; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3367 = 9'h11f == _GEN_14631 ? lru_287 : _GEN_3366; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3368 = 9'h120 == _GEN_14631 ? lru_288 : _GEN_3367; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3369 = 9'h121 == _GEN_14631 ? lru_289 : _GEN_3368; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3370 = 9'h122 == _GEN_14631 ? lru_290 : _GEN_3369; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3371 = 9'h123 == _GEN_14631 ? lru_291 : _GEN_3370; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3372 = 9'h124 == _GEN_14631 ? lru_292 : _GEN_3371; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3373 = 9'h125 == _GEN_14631 ? lru_293 : _GEN_3372; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3374 = 9'h126 == _GEN_14631 ? lru_294 : _GEN_3373; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3375 = 9'h127 == _GEN_14631 ? lru_295 : _GEN_3374; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3376 = 9'h128 == _GEN_14631 ? lru_296 : _GEN_3375; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3377 = 9'h129 == _GEN_14631 ? lru_297 : _GEN_3376; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3378 = 9'h12a == _GEN_14631 ? lru_298 : _GEN_3377; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3379 = 9'h12b == _GEN_14631 ? lru_299 : _GEN_3378; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3380 = 9'h12c == _GEN_14631 ? lru_300 : _GEN_3379; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3381 = 9'h12d == _GEN_14631 ? lru_301 : _GEN_3380; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3382 = 9'h12e == _GEN_14631 ? lru_302 : _GEN_3381; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3383 = 9'h12f == _GEN_14631 ? lru_303 : _GEN_3382; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3384 = 9'h130 == _GEN_14631 ? lru_304 : _GEN_3383; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3385 = 9'h131 == _GEN_14631 ? lru_305 : _GEN_3384; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3386 = 9'h132 == _GEN_14631 ? lru_306 : _GEN_3385; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3387 = 9'h133 == _GEN_14631 ? lru_307 : _GEN_3386; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3388 = 9'h134 == _GEN_14631 ? lru_308 : _GEN_3387; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3389 = 9'h135 == _GEN_14631 ? lru_309 : _GEN_3388; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3390 = 9'h136 == _GEN_14631 ? lru_310 : _GEN_3389; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3391 = 9'h137 == _GEN_14631 ? lru_311 : _GEN_3390; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3392 = 9'h138 == _GEN_14631 ? lru_312 : _GEN_3391; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3393 = 9'h139 == _GEN_14631 ? lru_313 : _GEN_3392; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3394 = 9'h13a == _GEN_14631 ? lru_314 : _GEN_3393; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3395 = 9'h13b == _GEN_14631 ? lru_315 : _GEN_3394; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3396 = 9'h13c == _GEN_14631 ? lru_316 : _GEN_3395; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3397 = 9'h13d == _GEN_14631 ? lru_317 : _GEN_3396; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3398 = 9'h13e == _GEN_14631 ? lru_318 : _GEN_3397; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3399 = 9'h13f == _GEN_14631 ? lru_319 : _GEN_3398; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3400 = 9'h140 == _GEN_14631 ? lru_320 : _GEN_3399; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3401 = 9'h141 == _GEN_14631 ? lru_321 : _GEN_3400; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3402 = 9'h142 == _GEN_14631 ? lru_322 : _GEN_3401; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3403 = 9'h143 == _GEN_14631 ? lru_323 : _GEN_3402; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3404 = 9'h144 == _GEN_14631 ? lru_324 : _GEN_3403; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3405 = 9'h145 == _GEN_14631 ? lru_325 : _GEN_3404; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3406 = 9'h146 == _GEN_14631 ? lru_326 : _GEN_3405; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3407 = 9'h147 == _GEN_14631 ? lru_327 : _GEN_3406; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3408 = 9'h148 == _GEN_14631 ? lru_328 : _GEN_3407; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3409 = 9'h149 == _GEN_14631 ? lru_329 : _GEN_3408; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3410 = 9'h14a == _GEN_14631 ? lru_330 : _GEN_3409; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3411 = 9'h14b == _GEN_14631 ? lru_331 : _GEN_3410; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3412 = 9'h14c == _GEN_14631 ? lru_332 : _GEN_3411; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3413 = 9'h14d == _GEN_14631 ? lru_333 : _GEN_3412; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3414 = 9'h14e == _GEN_14631 ? lru_334 : _GEN_3413; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3415 = 9'h14f == _GEN_14631 ? lru_335 : _GEN_3414; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3416 = 9'h150 == _GEN_14631 ? lru_336 : _GEN_3415; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3417 = 9'h151 == _GEN_14631 ? lru_337 : _GEN_3416; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3418 = 9'h152 == _GEN_14631 ? lru_338 : _GEN_3417; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3419 = 9'h153 == _GEN_14631 ? lru_339 : _GEN_3418; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3420 = 9'h154 == _GEN_14631 ? lru_340 : _GEN_3419; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3421 = 9'h155 == _GEN_14631 ? lru_341 : _GEN_3420; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3422 = 9'h156 == _GEN_14631 ? lru_342 : _GEN_3421; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3423 = 9'h157 == _GEN_14631 ? lru_343 : _GEN_3422; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3424 = 9'h158 == _GEN_14631 ? lru_344 : _GEN_3423; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3425 = 9'h159 == _GEN_14631 ? lru_345 : _GEN_3424; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3426 = 9'h15a == _GEN_14631 ? lru_346 : _GEN_3425; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3427 = 9'h15b == _GEN_14631 ? lru_347 : _GEN_3426; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3428 = 9'h15c == _GEN_14631 ? lru_348 : _GEN_3427; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3429 = 9'h15d == _GEN_14631 ? lru_349 : _GEN_3428; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3430 = 9'h15e == _GEN_14631 ? lru_350 : _GEN_3429; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3431 = 9'h15f == _GEN_14631 ? lru_351 : _GEN_3430; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3432 = 9'h160 == _GEN_14631 ? lru_352 : _GEN_3431; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3433 = 9'h161 == _GEN_14631 ? lru_353 : _GEN_3432; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3434 = 9'h162 == _GEN_14631 ? lru_354 : _GEN_3433; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3435 = 9'h163 == _GEN_14631 ? lru_355 : _GEN_3434; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3436 = 9'h164 == _GEN_14631 ? lru_356 : _GEN_3435; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3437 = 9'h165 == _GEN_14631 ? lru_357 : _GEN_3436; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3438 = 9'h166 == _GEN_14631 ? lru_358 : _GEN_3437; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3439 = 9'h167 == _GEN_14631 ? lru_359 : _GEN_3438; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3440 = 9'h168 == _GEN_14631 ? lru_360 : _GEN_3439; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3441 = 9'h169 == _GEN_14631 ? lru_361 : _GEN_3440; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3442 = 9'h16a == _GEN_14631 ? lru_362 : _GEN_3441; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3443 = 9'h16b == _GEN_14631 ? lru_363 : _GEN_3442; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3444 = 9'h16c == _GEN_14631 ? lru_364 : _GEN_3443; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3445 = 9'h16d == _GEN_14631 ? lru_365 : _GEN_3444; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3446 = 9'h16e == _GEN_14631 ? lru_366 : _GEN_3445; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3447 = 9'h16f == _GEN_14631 ? lru_367 : _GEN_3446; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3448 = 9'h170 == _GEN_14631 ? lru_368 : _GEN_3447; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3449 = 9'h171 == _GEN_14631 ? lru_369 : _GEN_3448; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3450 = 9'h172 == _GEN_14631 ? lru_370 : _GEN_3449; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3451 = 9'h173 == _GEN_14631 ? lru_371 : _GEN_3450; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3452 = 9'h174 == _GEN_14631 ? lru_372 : _GEN_3451; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3453 = 9'h175 == _GEN_14631 ? lru_373 : _GEN_3452; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3454 = 9'h176 == _GEN_14631 ? lru_374 : _GEN_3453; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3455 = 9'h177 == _GEN_14631 ? lru_375 : _GEN_3454; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3456 = 9'h178 == _GEN_14631 ? lru_376 : _GEN_3455; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3457 = 9'h179 == _GEN_14631 ? lru_377 : _GEN_3456; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3458 = 9'h17a == _GEN_14631 ? lru_378 : _GEN_3457; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3459 = 9'h17b == _GEN_14631 ? lru_379 : _GEN_3458; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3460 = 9'h17c == _GEN_14631 ? lru_380 : _GEN_3459; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3461 = 9'h17d == _GEN_14631 ? lru_381 : _GEN_3460; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3462 = 9'h17e == _GEN_14631 ? lru_382 : _GEN_3461; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3463 = 9'h17f == _GEN_14631 ? lru_383 : _GEN_3462; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3464 = 9'h180 == _GEN_14631 ? lru_384 : _GEN_3463; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3465 = 9'h181 == _GEN_14631 ? lru_385 : _GEN_3464; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3466 = 9'h182 == _GEN_14631 ? lru_386 : _GEN_3465; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3467 = 9'h183 == _GEN_14631 ? lru_387 : _GEN_3466; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3468 = 9'h184 == _GEN_14631 ? lru_388 : _GEN_3467; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3469 = 9'h185 == _GEN_14631 ? lru_389 : _GEN_3468; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3470 = 9'h186 == _GEN_14631 ? lru_390 : _GEN_3469; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3471 = 9'h187 == _GEN_14631 ? lru_391 : _GEN_3470; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3472 = 9'h188 == _GEN_14631 ? lru_392 : _GEN_3471; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3473 = 9'h189 == _GEN_14631 ? lru_393 : _GEN_3472; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3474 = 9'h18a == _GEN_14631 ? lru_394 : _GEN_3473; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3475 = 9'h18b == _GEN_14631 ? lru_395 : _GEN_3474; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3476 = 9'h18c == _GEN_14631 ? lru_396 : _GEN_3475; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3477 = 9'h18d == _GEN_14631 ? lru_397 : _GEN_3476; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3478 = 9'h18e == _GEN_14631 ? lru_398 : _GEN_3477; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3479 = 9'h18f == _GEN_14631 ? lru_399 : _GEN_3478; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3480 = 9'h190 == _GEN_14631 ? lru_400 : _GEN_3479; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3481 = 9'h191 == _GEN_14631 ? lru_401 : _GEN_3480; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3482 = 9'h192 == _GEN_14631 ? lru_402 : _GEN_3481; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3483 = 9'h193 == _GEN_14631 ? lru_403 : _GEN_3482; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3484 = 9'h194 == _GEN_14631 ? lru_404 : _GEN_3483; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3485 = 9'h195 == _GEN_14631 ? lru_405 : _GEN_3484; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3486 = 9'h196 == _GEN_14631 ? lru_406 : _GEN_3485; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3487 = 9'h197 == _GEN_14631 ? lru_407 : _GEN_3486; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3488 = 9'h198 == _GEN_14631 ? lru_408 : _GEN_3487; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3489 = 9'h199 == _GEN_14631 ? lru_409 : _GEN_3488; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3490 = 9'h19a == _GEN_14631 ? lru_410 : _GEN_3489; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3491 = 9'h19b == _GEN_14631 ? lru_411 : _GEN_3490; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3492 = 9'h19c == _GEN_14631 ? lru_412 : _GEN_3491; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3493 = 9'h19d == _GEN_14631 ? lru_413 : _GEN_3492; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3494 = 9'h19e == _GEN_14631 ? lru_414 : _GEN_3493; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3495 = 9'h19f == _GEN_14631 ? lru_415 : _GEN_3494; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3496 = 9'h1a0 == _GEN_14631 ? lru_416 : _GEN_3495; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3497 = 9'h1a1 == _GEN_14631 ? lru_417 : _GEN_3496; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3498 = 9'h1a2 == _GEN_14631 ? lru_418 : _GEN_3497; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3499 = 9'h1a3 == _GEN_14631 ? lru_419 : _GEN_3498; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3500 = 9'h1a4 == _GEN_14631 ? lru_420 : _GEN_3499; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3501 = 9'h1a5 == _GEN_14631 ? lru_421 : _GEN_3500; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3502 = 9'h1a6 == _GEN_14631 ? lru_422 : _GEN_3501; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3503 = 9'h1a7 == _GEN_14631 ? lru_423 : _GEN_3502; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3504 = 9'h1a8 == _GEN_14631 ? lru_424 : _GEN_3503; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3505 = 9'h1a9 == _GEN_14631 ? lru_425 : _GEN_3504; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3506 = 9'h1aa == _GEN_14631 ? lru_426 : _GEN_3505; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3507 = 9'h1ab == _GEN_14631 ? lru_427 : _GEN_3506; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3508 = 9'h1ac == _GEN_14631 ? lru_428 : _GEN_3507; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3509 = 9'h1ad == _GEN_14631 ? lru_429 : _GEN_3508; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3510 = 9'h1ae == _GEN_14631 ? lru_430 : _GEN_3509; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3511 = 9'h1af == _GEN_14631 ? lru_431 : _GEN_3510; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3512 = 9'h1b0 == _GEN_14631 ? lru_432 : _GEN_3511; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3513 = 9'h1b1 == _GEN_14631 ? lru_433 : _GEN_3512; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3514 = 9'h1b2 == _GEN_14631 ? lru_434 : _GEN_3513; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3515 = 9'h1b3 == _GEN_14631 ? lru_435 : _GEN_3514; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3516 = 9'h1b4 == _GEN_14631 ? lru_436 : _GEN_3515; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3517 = 9'h1b5 == _GEN_14631 ? lru_437 : _GEN_3516; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3518 = 9'h1b6 == _GEN_14631 ? lru_438 : _GEN_3517; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3519 = 9'h1b7 == _GEN_14631 ? lru_439 : _GEN_3518; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3520 = 9'h1b8 == _GEN_14631 ? lru_440 : _GEN_3519; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3521 = 9'h1b9 == _GEN_14631 ? lru_441 : _GEN_3520; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3522 = 9'h1ba == _GEN_14631 ? lru_442 : _GEN_3521; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3523 = 9'h1bb == _GEN_14631 ? lru_443 : _GEN_3522; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3524 = 9'h1bc == _GEN_14631 ? lru_444 : _GEN_3523; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3525 = 9'h1bd == _GEN_14631 ? lru_445 : _GEN_3524; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3526 = 9'h1be == _GEN_14631 ? lru_446 : _GEN_3525; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3527 = 9'h1bf == _GEN_14631 ? lru_447 : _GEN_3526; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3528 = 9'h1c0 == _GEN_14631 ? lru_448 : _GEN_3527; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3529 = 9'h1c1 == _GEN_14631 ? lru_449 : _GEN_3528; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3530 = 9'h1c2 == _GEN_14631 ? lru_450 : _GEN_3529; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3531 = 9'h1c3 == _GEN_14631 ? lru_451 : _GEN_3530; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3532 = 9'h1c4 == _GEN_14631 ? lru_452 : _GEN_3531; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3533 = 9'h1c5 == _GEN_14631 ? lru_453 : _GEN_3532; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3534 = 9'h1c6 == _GEN_14631 ? lru_454 : _GEN_3533; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3535 = 9'h1c7 == _GEN_14631 ? lru_455 : _GEN_3534; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3536 = 9'h1c8 == _GEN_14631 ? lru_456 : _GEN_3535; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3537 = 9'h1c9 == _GEN_14631 ? lru_457 : _GEN_3536; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3538 = 9'h1ca == _GEN_14631 ? lru_458 : _GEN_3537; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3539 = 9'h1cb == _GEN_14631 ? lru_459 : _GEN_3538; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3540 = 9'h1cc == _GEN_14631 ? lru_460 : _GEN_3539; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3541 = 9'h1cd == _GEN_14631 ? lru_461 : _GEN_3540; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3542 = 9'h1ce == _GEN_14631 ? lru_462 : _GEN_3541; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3543 = 9'h1cf == _GEN_14631 ? lru_463 : _GEN_3542; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3544 = 9'h1d0 == _GEN_14631 ? lru_464 : _GEN_3543; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3545 = 9'h1d1 == _GEN_14631 ? lru_465 : _GEN_3544; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3546 = 9'h1d2 == _GEN_14631 ? lru_466 : _GEN_3545; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3547 = 9'h1d3 == _GEN_14631 ? lru_467 : _GEN_3546; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3548 = 9'h1d4 == _GEN_14631 ? lru_468 : _GEN_3547; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3549 = 9'h1d5 == _GEN_14631 ? lru_469 : _GEN_3548; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3550 = 9'h1d6 == _GEN_14631 ? lru_470 : _GEN_3549; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3551 = 9'h1d7 == _GEN_14631 ? lru_471 : _GEN_3550; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3552 = 9'h1d8 == _GEN_14631 ? lru_472 : _GEN_3551; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3553 = 9'h1d9 == _GEN_14631 ? lru_473 : _GEN_3552; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3554 = 9'h1da == _GEN_14631 ? lru_474 : _GEN_3553; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3555 = 9'h1db == _GEN_14631 ? lru_475 : _GEN_3554; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3556 = 9'h1dc == _GEN_14631 ? lru_476 : _GEN_3555; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3557 = 9'h1dd == _GEN_14631 ? lru_477 : _GEN_3556; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3558 = 9'h1de == _GEN_14631 ? lru_478 : _GEN_3557; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3559 = 9'h1df == _GEN_14631 ? lru_479 : _GEN_3558; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3560 = 9'h1e0 == _GEN_14631 ? lru_480 : _GEN_3559; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3561 = 9'h1e1 == _GEN_14631 ? lru_481 : _GEN_3560; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3562 = 9'h1e2 == _GEN_14631 ? lru_482 : _GEN_3561; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3563 = 9'h1e3 == _GEN_14631 ? lru_483 : _GEN_3562; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3564 = 9'h1e4 == _GEN_14631 ? lru_484 : _GEN_3563; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3565 = 9'h1e5 == _GEN_14631 ? lru_485 : _GEN_3564; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3566 = 9'h1e6 == _GEN_14631 ? lru_486 : _GEN_3565; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3567 = 9'h1e7 == _GEN_14631 ? lru_487 : _GEN_3566; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3568 = 9'h1e8 == _GEN_14631 ? lru_488 : _GEN_3567; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3569 = 9'h1e9 == _GEN_14631 ? lru_489 : _GEN_3568; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3570 = 9'h1ea == _GEN_14631 ? lru_490 : _GEN_3569; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3571 = 9'h1eb == _GEN_14631 ? lru_491 : _GEN_3570; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3572 = 9'h1ec == _GEN_14631 ? lru_492 : _GEN_3571; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3573 = 9'h1ed == _GEN_14631 ? lru_493 : _GEN_3572; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3574 = 9'h1ee == _GEN_14631 ? lru_494 : _GEN_3573; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3575 = 9'h1ef == _GEN_14631 ? lru_495 : _GEN_3574; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3576 = 9'h1f0 == _GEN_14631 ? lru_496 : _GEN_3575; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3577 = 9'h1f1 == _GEN_14631 ? lru_497 : _GEN_3576; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3578 = 9'h1f2 == _GEN_14631 ? lru_498 : _GEN_3577; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3579 = 9'h1f3 == _GEN_14631 ? lru_499 : _GEN_3578; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3580 = 9'h1f4 == _GEN_14631 ? lru_500 : _GEN_3579; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3581 = 9'h1f5 == _GEN_14631 ? lru_501 : _GEN_3580; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3582 = 9'h1f6 == _GEN_14631 ? lru_502 : _GEN_3581; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3583 = 9'h1f7 == _GEN_14631 ? lru_503 : _GEN_3582; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3584 = 9'h1f8 == _GEN_14631 ? lru_504 : _GEN_3583; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3585 = 9'h1f9 == _GEN_14631 ? lru_505 : _GEN_3584; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3586 = 9'h1fa == _GEN_14631 ? lru_506 : _GEN_3585; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3587 = 9'h1fb == _GEN_14631 ? lru_507 : _GEN_3586; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3588 = 9'h1fc == _GEN_14631 ? lru_508 : _GEN_3587; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3589 = 9'h1fd == _GEN_14631 ? lru_509 : _GEN_3588; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3590 = 9'h1fe == _GEN_14631 ? lru_510 : _GEN_3589; // @[ICache.scala 183:{36,36}]
  wire  _GEN_3591 = 9'h1ff == _GEN_14631 ? lru_511 : _GEN_3590; // @[ICache.scala 183:{36,36}]
  wire [3:0] _GEN_3592 = ~_GEN_3591 ? 4'hf : data_wstrb_0_0; // @[ICache.scala 183:{36,36} 61:27]
  wire [3:0] _GEN_3593 = _GEN_3591 ? 4'hf : data_wstrb_1_0; // @[ICache.scala 183:{36,36} 61:27]
  wire [3:0] _GEN_3594 = ~_GEN_3591 ? 4'h0 : data_wstrb_0_1; // @[ICache.scala 184:{36,36} 61:27]
  wire [3:0] _GEN_3595 = _GEN_3591 ? 4'h0 : data_wstrb_1_1; // @[ICache.scala 184:{36,36} 61:27]
  wire  _GEN_15783 = ~_GEN_3591; // @[ICache.scala 185:{36,36} 64:26]
  wire  _GEN_3596 = ~_GEN_3591 | tag_wstrb_0; // @[ICache.scala 185:{36,36} 64:26]
  wire  _GEN_3597 = _GEN_3591 | tag_wstrb_1; // @[ICache.scala 185:{36,36} 64:26]
  wire  _GEN_3598 = 6'h0 == vset & _GEN_15783 | _GEN_1027; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3599 = 6'h0 == vset & _GEN_3591 | _GEN_1539; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3600 = 6'h1 == vset & _GEN_15783 | _GEN_1028; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3601 = 6'h1 == vset & _GEN_3591 | _GEN_1540; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3602 = 6'h2 == vset & _GEN_15783 | _GEN_1029; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3603 = 6'h2 == vset & _GEN_3591 | _GEN_1541; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3604 = 6'h3 == vset & _GEN_15783 | _GEN_1030; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3605 = 6'h3 == vset & _GEN_3591 | _GEN_1542; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3606 = 6'h4 == vset & _GEN_15783 | _GEN_1031; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3607 = 6'h4 == vset & _GEN_3591 | _GEN_1543; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3608 = 6'h5 == vset & _GEN_15783 | _GEN_1032; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3609 = 6'h5 == vset & _GEN_3591 | _GEN_1544; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3610 = 6'h6 == vset & _GEN_15783 | _GEN_1033; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3611 = 6'h6 == vset & _GEN_3591 | _GEN_1545; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3612 = 6'h7 == vset & _GEN_15783 | _GEN_1034; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3613 = 6'h7 == vset & _GEN_3591 | _GEN_1546; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3614 = 6'h8 == vset & _GEN_15783 | _GEN_1035; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3615 = 6'h8 == vset & _GEN_3591 | _GEN_1547; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3616 = 6'h9 == vset & _GEN_15783 | _GEN_1036; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3617 = 6'h9 == vset & _GEN_3591 | _GEN_1548; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3618 = 6'ha == vset & _GEN_15783 | _GEN_1037; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3619 = 6'ha == vset & _GEN_3591 | _GEN_1549; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3620 = 6'hb == vset & _GEN_15783 | _GEN_1038; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3621 = 6'hb == vset & _GEN_3591 | _GEN_1550; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3622 = 6'hc == vset & _GEN_15783 | _GEN_1039; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3623 = 6'hc == vset & _GEN_3591 | _GEN_1551; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3624 = 6'hd == vset & _GEN_15783 | _GEN_1040; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3625 = 6'hd == vset & _GEN_3591 | _GEN_1552; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3626 = 6'he == vset & _GEN_15783 | _GEN_1041; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3627 = 6'he == vset & _GEN_3591 | _GEN_1553; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3628 = 6'hf == vset & _GEN_15783 | _GEN_1042; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3629 = 6'hf == vset & _GEN_3591 | _GEN_1554; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3630 = 6'h10 == vset & _GEN_15783 | _GEN_1043; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3631 = 6'h10 == vset & _GEN_3591 | _GEN_1555; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3632 = 6'h11 == vset & _GEN_15783 | _GEN_1044; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3633 = 6'h11 == vset & _GEN_3591 | _GEN_1556; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3634 = 6'h12 == vset & _GEN_15783 | _GEN_1045; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3635 = 6'h12 == vset & _GEN_3591 | _GEN_1557; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3636 = 6'h13 == vset & _GEN_15783 | _GEN_1046; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3637 = 6'h13 == vset & _GEN_3591 | _GEN_1558; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3638 = 6'h14 == vset & _GEN_15783 | _GEN_1047; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3639 = 6'h14 == vset & _GEN_3591 | _GEN_1559; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3640 = 6'h15 == vset & _GEN_15783 | _GEN_1048; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3641 = 6'h15 == vset & _GEN_3591 | _GEN_1560; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3642 = 6'h16 == vset & _GEN_15783 | _GEN_1049; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3643 = 6'h16 == vset & _GEN_3591 | _GEN_1561; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3644 = 6'h17 == vset & _GEN_15783 | _GEN_1050; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3645 = 6'h17 == vset & _GEN_3591 | _GEN_1562; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3646 = 6'h18 == vset & _GEN_15783 | _GEN_1051; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3647 = 6'h18 == vset & _GEN_3591 | _GEN_1563; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3648 = 6'h19 == vset & _GEN_15783 | _GEN_1052; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3649 = 6'h19 == vset & _GEN_3591 | _GEN_1564; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3650 = 6'h1a == vset & _GEN_15783 | _GEN_1053; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3651 = 6'h1a == vset & _GEN_3591 | _GEN_1565; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3652 = 6'h1b == vset & _GEN_15783 | _GEN_1054; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3653 = 6'h1b == vset & _GEN_3591 | _GEN_1566; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3654 = 6'h1c == vset & _GEN_15783 | _GEN_1055; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3655 = 6'h1c == vset & _GEN_3591 | _GEN_1567; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3656 = 6'h1d == vset & _GEN_15783 | _GEN_1056; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3657 = 6'h1d == vset & _GEN_3591 | _GEN_1568; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3658 = 6'h1e == vset & _GEN_15783 | _GEN_1057; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3659 = 6'h1e == vset & _GEN_3591 | _GEN_1569; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3660 = 6'h1f == vset & _GEN_15783 | _GEN_1058; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3661 = 6'h1f == vset & _GEN_3591 | _GEN_1570; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3662 = 6'h20 == vset & _GEN_15783 | _GEN_1059; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3663 = 6'h20 == vset & _GEN_3591 | _GEN_1571; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3664 = 6'h21 == vset & _GEN_15783 | _GEN_1060; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3665 = 6'h21 == vset & _GEN_3591 | _GEN_1572; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3666 = 6'h22 == vset & _GEN_15783 | _GEN_1061; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3667 = 6'h22 == vset & _GEN_3591 | _GEN_1573; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3668 = 6'h23 == vset & _GEN_15783 | _GEN_1062; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3669 = 6'h23 == vset & _GEN_3591 | _GEN_1574; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3670 = 6'h24 == vset & _GEN_15783 | _GEN_1063; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3671 = 6'h24 == vset & _GEN_3591 | _GEN_1575; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3672 = 6'h25 == vset & _GEN_15783 | _GEN_1064; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3673 = 6'h25 == vset & _GEN_3591 | _GEN_1576; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3674 = 6'h26 == vset & _GEN_15783 | _GEN_1065; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3675 = 6'h26 == vset & _GEN_3591 | _GEN_1577; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3676 = 6'h27 == vset & _GEN_15783 | _GEN_1066; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3677 = 6'h27 == vset & _GEN_3591 | _GEN_1578; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3678 = 6'h28 == vset & _GEN_15783 | _GEN_1067; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3679 = 6'h28 == vset & _GEN_3591 | _GEN_1579; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3680 = 6'h29 == vset & _GEN_15783 | _GEN_1068; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3681 = 6'h29 == vset & _GEN_3591 | _GEN_1580; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3682 = 6'h2a == vset & _GEN_15783 | _GEN_1069; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3683 = 6'h2a == vset & _GEN_3591 | _GEN_1581; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3684 = 6'h2b == vset & _GEN_15783 | _GEN_1070; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3685 = 6'h2b == vset & _GEN_3591 | _GEN_1582; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3686 = 6'h2c == vset & _GEN_15783 | _GEN_1071; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3687 = 6'h2c == vset & _GEN_3591 | _GEN_1583; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3688 = 6'h2d == vset & _GEN_15783 | _GEN_1072; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3689 = 6'h2d == vset & _GEN_3591 | _GEN_1584; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3690 = 6'h2e == vset & _GEN_15783 | _GEN_1073; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3691 = 6'h2e == vset & _GEN_3591 | _GEN_1585; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3692 = 6'h2f == vset & _GEN_15783 | _GEN_1074; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3693 = 6'h2f == vset & _GEN_3591 | _GEN_1586; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3694 = 6'h30 == vset & _GEN_15783 | _GEN_1075; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3695 = 6'h30 == vset & _GEN_3591 | _GEN_1587; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3696 = 6'h31 == vset & _GEN_15783 | _GEN_1076; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3697 = 6'h31 == vset & _GEN_3591 | _GEN_1588; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3698 = 6'h32 == vset & _GEN_15783 | _GEN_1077; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3699 = 6'h32 == vset & _GEN_3591 | _GEN_1589; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3700 = 6'h33 == vset & _GEN_15783 | _GEN_1078; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3701 = 6'h33 == vset & _GEN_3591 | _GEN_1590; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3702 = 6'h34 == vset & _GEN_15783 | _GEN_1079; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3703 = 6'h34 == vset & _GEN_3591 | _GEN_1591; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3704 = 6'h35 == vset & _GEN_15783 | _GEN_1080; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3705 = 6'h35 == vset & _GEN_3591 | _GEN_1592; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3706 = 6'h36 == vset & _GEN_15783 | _GEN_1081; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3707 = 6'h36 == vset & _GEN_3591 | _GEN_1593; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3708 = 6'h37 == vset & _GEN_15783 | _GEN_1082; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3709 = 6'h37 == vset & _GEN_3591 | _GEN_1594; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3710 = 6'h38 == vset & _GEN_15783 | _GEN_1083; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3711 = 6'h38 == vset & _GEN_3591 | _GEN_1595; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3712 = 6'h39 == vset & _GEN_15783 | _GEN_1084; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3713 = 6'h39 == vset & _GEN_3591 | _GEN_1596; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3714 = 6'h3a == vset & _GEN_15783 | _GEN_1085; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3715 = 6'h3a == vset & _GEN_3591 | _GEN_1597; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3716 = 6'h3b == vset & _GEN_15783 | _GEN_1086; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3717 = 6'h3b == vset & _GEN_3591 | _GEN_1598; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3718 = 6'h3c == vset & _GEN_15783 | _GEN_1087; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3719 = 6'h3c == vset & _GEN_3591 | _GEN_1599; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3720 = 6'h3d == vset & _GEN_15783 | _GEN_1088; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3721 = 6'h3d == vset & _GEN_3591 | _GEN_1600; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3722 = 6'h3e == vset & _GEN_15783 | _GEN_1089; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3723 = 6'h3e == vset & _GEN_3591 | _GEN_1601; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3724 = 6'h3f == vset & _GEN_15783 | _GEN_1090; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3725 = 6'h3f == vset & _GEN_3591 | _GEN_1602; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3726 = 7'h40 == _GEN_14439 & _GEN_15783 | _GEN_1091; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3727 = 7'h40 == _GEN_14439 & _GEN_3591 | _GEN_1603; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3728 = 7'h41 == _GEN_14439 & _GEN_15783 | _GEN_1092; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3729 = 7'h41 == _GEN_14439 & _GEN_3591 | _GEN_1604; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3730 = 7'h42 == _GEN_14439 & _GEN_15783 | _GEN_1093; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3731 = 7'h42 == _GEN_14439 & _GEN_3591 | _GEN_1605; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3732 = 7'h43 == _GEN_14439 & _GEN_15783 | _GEN_1094; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3733 = 7'h43 == _GEN_14439 & _GEN_3591 | _GEN_1606; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3734 = 7'h44 == _GEN_14439 & _GEN_15783 | _GEN_1095; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3735 = 7'h44 == _GEN_14439 & _GEN_3591 | _GEN_1607; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3736 = 7'h45 == _GEN_14439 & _GEN_15783 | _GEN_1096; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3737 = 7'h45 == _GEN_14439 & _GEN_3591 | _GEN_1608; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3738 = 7'h46 == _GEN_14439 & _GEN_15783 | _GEN_1097; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3739 = 7'h46 == _GEN_14439 & _GEN_3591 | _GEN_1609; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3740 = 7'h47 == _GEN_14439 & _GEN_15783 | _GEN_1098; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3741 = 7'h47 == _GEN_14439 & _GEN_3591 | _GEN_1610; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3742 = 7'h48 == _GEN_14439 & _GEN_15783 | _GEN_1099; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3743 = 7'h48 == _GEN_14439 & _GEN_3591 | _GEN_1611; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3744 = 7'h49 == _GEN_14439 & _GEN_15783 | _GEN_1100; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3745 = 7'h49 == _GEN_14439 & _GEN_3591 | _GEN_1612; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3746 = 7'h4a == _GEN_14439 & _GEN_15783 | _GEN_1101; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3747 = 7'h4a == _GEN_14439 & _GEN_3591 | _GEN_1613; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3748 = 7'h4b == _GEN_14439 & _GEN_15783 | _GEN_1102; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3749 = 7'h4b == _GEN_14439 & _GEN_3591 | _GEN_1614; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3750 = 7'h4c == _GEN_14439 & _GEN_15783 | _GEN_1103; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3751 = 7'h4c == _GEN_14439 & _GEN_3591 | _GEN_1615; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3752 = 7'h4d == _GEN_14439 & _GEN_15783 | _GEN_1104; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3753 = 7'h4d == _GEN_14439 & _GEN_3591 | _GEN_1616; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3754 = 7'h4e == _GEN_14439 & _GEN_15783 | _GEN_1105; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3755 = 7'h4e == _GEN_14439 & _GEN_3591 | _GEN_1617; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3756 = 7'h4f == _GEN_14439 & _GEN_15783 | _GEN_1106; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3757 = 7'h4f == _GEN_14439 & _GEN_3591 | _GEN_1618; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3758 = 7'h50 == _GEN_14439 & _GEN_15783 | _GEN_1107; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3759 = 7'h50 == _GEN_14439 & _GEN_3591 | _GEN_1619; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3760 = 7'h51 == _GEN_14439 & _GEN_15783 | _GEN_1108; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3761 = 7'h51 == _GEN_14439 & _GEN_3591 | _GEN_1620; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3762 = 7'h52 == _GEN_14439 & _GEN_15783 | _GEN_1109; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3763 = 7'h52 == _GEN_14439 & _GEN_3591 | _GEN_1621; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3764 = 7'h53 == _GEN_14439 & _GEN_15783 | _GEN_1110; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3765 = 7'h53 == _GEN_14439 & _GEN_3591 | _GEN_1622; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3766 = 7'h54 == _GEN_14439 & _GEN_15783 | _GEN_1111; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3767 = 7'h54 == _GEN_14439 & _GEN_3591 | _GEN_1623; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3768 = 7'h55 == _GEN_14439 & _GEN_15783 | _GEN_1112; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3769 = 7'h55 == _GEN_14439 & _GEN_3591 | _GEN_1624; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3770 = 7'h56 == _GEN_14439 & _GEN_15783 | _GEN_1113; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3771 = 7'h56 == _GEN_14439 & _GEN_3591 | _GEN_1625; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3772 = 7'h57 == _GEN_14439 & _GEN_15783 | _GEN_1114; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3773 = 7'h57 == _GEN_14439 & _GEN_3591 | _GEN_1626; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3774 = 7'h58 == _GEN_14439 & _GEN_15783 | _GEN_1115; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3775 = 7'h58 == _GEN_14439 & _GEN_3591 | _GEN_1627; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3776 = 7'h59 == _GEN_14439 & _GEN_15783 | _GEN_1116; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3777 = 7'h59 == _GEN_14439 & _GEN_3591 | _GEN_1628; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3778 = 7'h5a == _GEN_14439 & _GEN_15783 | _GEN_1117; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3779 = 7'h5a == _GEN_14439 & _GEN_3591 | _GEN_1629; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3780 = 7'h5b == _GEN_14439 & _GEN_15783 | _GEN_1118; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3781 = 7'h5b == _GEN_14439 & _GEN_3591 | _GEN_1630; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3782 = 7'h5c == _GEN_14439 & _GEN_15783 | _GEN_1119; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3783 = 7'h5c == _GEN_14439 & _GEN_3591 | _GEN_1631; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3784 = 7'h5d == _GEN_14439 & _GEN_15783 | _GEN_1120; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3785 = 7'h5d == _GEN_14439 & _GEN_3591 | _GEN_1632; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3786 = 7'h5e == _GEN_14439 & _GEN_15783 | _GEN_1121; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3787 = 7'h5e == _GEN_14439 & _GEN_3591 | _GEN_1633; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3788 = 7'h5f == _GEN_14439 & _GEN_15783 | _GEN_1122; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3789 = 7'h5f == _GEN_14439 & _GEN_3591 | _GEN_1634; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3790 = 7'h60 == _GEN_14439 & _GEN_15783 | _GEN_1123; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3791 = 7'h60 == _GEN_14439 & _GEN_3591 | _GEN_1635; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3792 = 7'h61 == _GEN_14439 & _GEN_15783 | _GEN_1124; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3793 = 7'h61 == _GEN_14439 & _GEN_3591 | _GEN_1636; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3794 = 7'h62 == _GEN_14439 & _GEN_15783 | _GEN_1125; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3795 = 7'h62 == _GEN_14439 & _GEN_3591 | _GEN_1637; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3796 = 7'h63 == _GEN_14439 & _GEN_15783 | _GEN_1126; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3797 = 7'h63 == _GEN_14439 & _GEN_3591 | _GEN_1638; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3798 = 7'h64 == _GEN_14439 & _GEN_15783 | _GEN_1127; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3799 = 7'h64 == _GEN_14439 & _GEN_3591 | _GEN_1639; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3800 = 7'h65 == _GEN_14439 & _GEN_15783 | _GEN_1128; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3801 = 7'h65 == _GEN_14439 & _GEN_3591 | _GEN_1640; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3802 = 7'h66 == _GEN_14439 & _GEN_15783 | _GEN_1129; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3803 = 7'h66 == _GEN_14439 & _GEN_3591 | _GEN_1641; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3804 = 7'h67 == _GEN_14439 & _GEN_15783 | _GEN_1130; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3805 = 7'h67 == _GEN_14439 & _GEN_3591 | _GEN_1642; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3806 = 7'h68 == _GEN_14439 & _GEN_15783 | _GEN_1131; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3807 = 7'h68 == _GEN_14439 & _GEN_3591 | _GEN_1643; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3808 = 7'h69 == _GEN_14439 & _GEN_15783 | _GEN_1132; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3809 = 7'h69 == _GEN_14439 & _GEN_3591 | _GEN_1644; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3810 = 7'h6a == _GEN_14439 & _GEN_15783 | _GEN_1133; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3811 = 7'h6a == _GEN_14439 & _GEN_3591 | _GEN_1645; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3812 = 7'h6b == _GEN_14439 & _GEN_15783 | _GEN_1134; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3813 = 7'h6b == _GEN_14439 & _GEN_3591 | _GEN_1646; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3814 = 7'h6c == _GEN_14439 & _GEN_15783 | _GEN_1135; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3815 = 7'h6c == _GEN_14439 & _GEN_3591 | _GEN_1647; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3816 = 7'h6d == _GEN_14439 & _GEN_15783 | _GEN_1136; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3817 = 7'h6d == _GEN_14439 & _GEN_3591 | _GEN_1648; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3818 = 7'h6e == _GEN_14439 & _GEN_15783 | _GEN_1137; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3819 = 7'h6e == _GEN_14439 & _GEN_3591 | _GEN_1649; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3820 = 7'h6f == _GEN_14439 & _GEN_15783 | _GEN_1138; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3821 = 7'h6f == _GEN_14439 & _GEN_3591 | _GEN_1650; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3822 = 7'h70 == _GEN_14439 & _GEN_15783 | _GEN_1139; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3823 = 7'h70 == _GEN_14439 & _GEN_3591 | _GEN_1651; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3824 = 7'h71 == _GEN_14439 & _GEN_15783 | _GEN_1140; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3825 = 7'h71 == _GEN_14439 & _GEN_3591 | _GEN_1652; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3826 = 7'h72 == _GEN_14439 & _GEN_15783 | _GEN_1141; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3827 = 7'h72 == _GEN_14439 & _GEN_3591 | _GEN_1653; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3828 = 7'h73 == _GEN_14439 & _GEN_15783 | _GEN_1142; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3829 = 7'h73 == _GEN_14439 & _GEN_3591 | _GEN_1654; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3830 = 7'h74 == _GEN_14439 & _GEN_15783 | _GEN_1143; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3831 = 7'h74 == _GEN_14439 & _GEN_3591 | _GEN_1655; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3832 = 7'h75 == _GEN_14439 & _GEN_15783 | _GEN_1144; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3833 = 7'h75 == _GEN_14439 & _GEN_3591 | _GEN_1656; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3834 = 7'h76 == _GEN_14439 & _GEN_15783 | _GEN_1145; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3835 = 7'h76 == _GEN_14439 & _GEN_3591 | _GEN_1657; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3836 = 7'h77 == _GEN_14439 & _GEN_15783 | _GEN_1146; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3837 = 7'h77 == _GEN_14439 & _GEN_3591 | _GEN_1658; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3838 = 7'h78 == _GEN_14439 & _GEN_15783 | _GEN_1147; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3839 = 7'h78 == _GEN_14439 & _GEN_3591 | _GEN_1659; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3840 = 7'h79 == _GEN_14439 & _GEN_15783 | _GEN_1148; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3841 = 7'h79 == _GEN_14439 & _GEN_3591 | _GEN_1660; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3842 = 7'h7a == _GEN_14439 & _GEN_15783 | _GEN_1149; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3843 = 7'h7a == _GEN_14439 & _GEN_3591 | _GEN_1661; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3844 = 7'h7b == _GEN_14439 & _GEN_15783 | _GEN_1150; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3845 = 7'h7b == _GEN_14439 & _GEN_3591 | _GEN_1662; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3846 = 7'h7c == _GEN_14439 & _GEN_15783 | _GEN_1151; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3847 = 7'h7c == _GEN_14439 & _GEN_3591 | _GEN_1663; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3848 = 7'h7d == _GEN_14439 & _GEN_15783 | _GEN_1152; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3849 = 7'h7d == _GEN_14439 & _GEN_3591 | _GEN_1664; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3850 = 7'h7e == _GEN_14439 & _GEN_15783 | _GEN_1153; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3851 = 7'h7e == _GEN_14439 & _GEN_3591 | _GEN_1665; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3852 = 7'h7f == _GEN_14439 & _GEN_15783 | _GEN_1154; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3853 = 7'h7f == _GEN_14439 & _GEN_3591 | _GEN_1666; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3854 = 8'h80 == _GEN_14503 & _GEN_15783 | _GEN_1155; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3855 = 8'h80 == _GEN_14503 & _GEN_3591 | _GEN_1667; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3856 = 8'h81 == _GEN_14503 & _GEN_15783 | _GEN_1156; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3857 = 8'h81 == _GEN_14503 & _GEN_3591 | _GEN_1668; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3858 = 8'h82 == _GEN_14503 & _GEN_15783 | _GEN_1157; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3859 = 8'h82 == _GEN_14503 & _GEN_3591 | _GEN_1669; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3860 = 8'h83 == _GEN_14503 & _GEN_15783 | _GEN_1158; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3861 = 8'h83 == _GEN_14503 & _GEN_3591 | _GEN_1670; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3862 = 8'h84 == _GEN_14503 & _GEN_15783 | _GEN_1159; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3863 = 8'h84 == _GEN_14503 & _GEN_3591 | _GEN_1671; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3864 = 8'h85 == _GEN_14503 & _GEN_15783 | _GEN_1160; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3865 = 8'h85 == _GEN_14503 & _GEN_3591 | _GEN_1672; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3866 = 8'h86 == _GEN_14503 & _GEN_15783 | _GEN_1161; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3867 = 8'h86 == _GEN_14503 & _GEN_3591 | _GEN_1673; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3868 = 8'h87 == _GEN_14503 & _GEN_15783 | _GEN_1162; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3869 = 8'h87 == _GEN_14503 & _GEN_3591 | _GEN_1674; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3870 = 8'h88 == _GEN_14503 & _GEN_15783 | _GEN_1163; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3871 = 8'h88 == _GEN_14503 & _GEN_3591 | _GEN_1675; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3872 = 8'h89 == _GEN_14503 & _GEN_15783 | _GEN_1164; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3873 = 8'h89 == _GEN_14503 & _GEN_3591 | _GEN_1676; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3874 = 8'h8a == _GEN_14503 & _GEN_15783 | _GEN_1165; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3875 = 8'h8a == _GEN_14503 & _GEN_3591 | _GEN_1677; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3876 = 8'h8b == _GEN_14503 & _GEN_15783 | _GEN_1166; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3877 = 8'h8b == _GEN_14503 & _GEN_3591 | _GEN_1678; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3878 = 8'h8c == _GEN_14503 & _GEN_15783 | _GEN_1167; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3879 = 8'h8c == _GEN_14503 & _GEN_3591 | _GEN_1679; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3880 = 8'h8d == _GEN_14503 & _GEN_15783 | _GEN_1168; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3881 = 8'h8d == _GEN_14503 & _GEN_3591 | _GEN_1680; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3882 = 8'h8e == _GEN_14503 & _GEN_15783 | _GEN_1169; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3883 = 8'h8e == _GEN_14503 & _GEN_3591 | _GEN_1681; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3884 = 8'h8f == _GEN_14503 & _GEN_15783 | _GEN_1170; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3885 = 8'h8f == _GEN_14503 & _GEN_3591 | _GEN_1682; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3886 = 8'h90 == _GEN_14503 & _GEN_15783 | _GEN_1171; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3887 = 8'h90 == _GEN_14503 & _GEN_3591 | _GEN_1683; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3888 = 8'h91 == _GEN_14503 & _GEN_15783 | _GEN_1172; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3889 = 8'h91 == _GEN_14503 & _GEN_3591 | _GEN_1684; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3890 = 8'h92 == _GEN_14503 & _GEN_15783 | _GEN_1173; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3891 = 8'h92 == _GEN_14503 & _GEN_3591 | _GEN_1685; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3892 = 8'h93 == _GEN_14503 & _GEN_15783 | _GEN_1174; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3893 = 8'h93 == _GEN_14503 & _GEN_3591 | _GEN_1686; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3894 = 8'h94 == _GEN_14503 & _GEN_15783 | _GEN_1175; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3895 = 8'h94 == _GEN_14503 & _GEN_3591 | _GEN_1687; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3896 = 8'h95 == _GEN_14503 & _GEN_15783 | _GEN_1176; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3897 = 8'h95 == _GEN_14503 & _GEN_3591 | _GEN_1688; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3898 = 8'h96 == _GEN_14503 & _GEN_15783 | _GEN_1177; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3899 = 8'h96 == _GEN_14503 & _GEN_3591 | _GEN_1689; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3900 = 8'h97 == _GEN_14503 & _GEN_15783 | _GEN_1178; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3901 = 8'h97 == _GEN_14503 & _GEN_3591 | _GEN_1690; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3902 = 8'h98 == _GEN_14503 & _GEN_15783 | _GEN_1179; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3903 = 8'h98 == _GEN_14503 & _GEN_3591 | _GEN_1691; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3904 = 8'h99 == _GEN_14503 & _GEN_15783 | _GEN_1180; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3905 = 8'h99 == _GEN_14503 & _GEN_3591 | _GEN_1692; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3906 = 8'h9a == _GEN_14503 & _GEN_15783 | _GEN_1181; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3907 = 8'h9a == _GEN_14503 & _GEN_3591 | _GEN_1693; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3908 = 8'h9b == _GEN_14503 & _GEN_15783 | _GEN_1182; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3909 = 8'h9b == _GEN_14503 & _GEN_3591 | _GEN_1694; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3910 = 8'h9c == _GEN_14503 & _GEN_15783 | _GEN_1183; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3911 = 8'h9c == _GEN_14503 & _GEN_3591 | _GEN_1695; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3912 = 8'h9d == _GEN_14503 & _GEN_15783 | _GEN_1184; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3913 = 8'h9d == _GEN_14503 & _GEN_3591 | _GEN_1696; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3914 = 8'h9e == _GEN_14503 & _GEN_15783 | _GEN_1185; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3915 = 8'h9e == _GEN_14503 & _GEN_3591 | _GEN_1697; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3916 = 8'h9f == _GEN_14503 & _GEN_15783 | _GEN_1186; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3917 = 8'h9f == _GEN_14503 & _GEN_3591 | _GEN_1698; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3918 = 8'ha0 == _GEN_14503 & _GEN_15783 | _GEN_1187; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3919 = 8'ha0 == _GEN_14503 & _GEN_3591 | _GEN_1699; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3920 = 8'ha1 == _GEN_14503 & _GEN_15783 | _GEN_1188; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3921 = 8'ha1 == _GEN_14503 & _GEN_3591 | _GEN_1700; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3922 = 8'ha2 == _GEN_14503 & _GEN_15783 | _GEN_1189; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3923 = 8'ha2 == _GEN_14503 & _GEN_3591 | _GEN_1701; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3924 = 8'ha3 == _GEN_14503 & _GEN_15783 | _GEN_1190; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3925 = 8'ha3 == _GEN_14503 & _GEN_3591 | _GEN_1702; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3926 = 8'ha4 == _GEN_14503 & _GEN_15783 | _GEN_1191; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3927 = 8'ha4 == _GEN_14503 & _GEN_3591 | _GEN_1703; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3928 = 8'ha5 == _GEN_14503 & _GEN_15783 | _GEN_1192; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3929 = 8'ha5 == _GEN_14503 & _GEN_3591 | _GEN_1704; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3930 = 8'ha6 == _GEN_14503 & _GEN_15783 | _GEN_1193; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3931 = 8'ha6 == _GEN_14503 & _GEN_3591 | _GEN_1705; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3932 = 8'ha7 == _GEN_14503 & _GEN_15783 | _GEN_1194; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3933 = 8'ha7 == _GEN_14503 & _GEN_3591 | _GEN_1706; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3934 = 8'ha8 == _GEN_14503 & _GEN_15783 | _GEN_1195; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3935 = 8'ha8 == _GEN_14503 & _GEN_3591 | _GEN_1707; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3936 = 8'ha9 == _GEN_14503 & _GEN_15783 | _GEN_1196; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3937 = 8'ha9 == _GEN_14503 & _GEN_3591 | _GEN_1708; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3938 = 8'haa == _GEN_14503 & _GEN_15783 | _GEN_1197; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3939 = 8'haa == _GEN_14503 & _GEN_3591 | _GEN_1709; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3940 = 8'hab == _GEN_14503 & _GEN_15783 | _GEN_1198; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3941 = 8'hab == _GEN_14503 & _GEN_3591 | _GEN_1710; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3942 = 8'hac == _GEN_14503 & _GEN_15783 | _GEN_1199; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3943 = 8'hac == _GEN_14503 & _GEN_3591 | _GEN_1711; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3944 = 8'had == _GEN_14503 & _GEN_15783 | _GEN_1200; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3945 = 8'had == _GEN_14503 & _GEN_3591 | _GEN_1712; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3946 = 8'hae == _GEN_14503 & _GEN_15783 | _GEN_1201; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3947 = 8'hae == _GEN_14503 & _GEN_3591 | _GEN_1713; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3948 = 8'haf == _GEN_14503 & _GEN_15783 | _GEN_1202; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3949 = 8'haf == _GEN_14503 & _GEN_3591 | _GEN_1714; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3950 = 8'hb0 == _GEN_14503 & _GEN_15783 | _GEN_1203; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3951 = 8'hb0 == _GEN_14503 & _GEN_3591 | _GEN_1715; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3952 = 8'hb1 == _GEN_14503 & _GEN_15783 | _GEN_1204; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3953 = 8'hb1 == _GEN_14503 & _GEN_3591 | _GEN_1716; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3954 = 8'hb2 == _GEN_14503 & _GEN_15783 | _GEN_1205; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3955 = 8'hb2 == _GEN_14503 & _GEN_3591 | _GEN_1717; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3956 = 8'hb3 == _GEN_14503 & _GEN_15783 | _GEN_1206; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3957 = 8'hb3 == _GEN_14503 & _GEN_3591 | _GEN_1718; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3958 = 8'hb4 == _GEN_14503 & _GEN_15783 | _GEN_1207; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3959 = 8'hb4 == _GEN_14503 & _GEN_3591 | _GEN_1719; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3960 = 8'hb5 == _GEN_14503 & _GEN_15783 | _GEN_1208; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3961 = 8'hb5 == _GEN_14503 & _GEN_3591 | _GEN_1720; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3962 = 8'hb6 == _GEN_14503 & _GEN_15783 | _GEN_1209; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3963 = 8'hb6 == _GEN_14503 & _GEN_3591 | _GEN_1721; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3964 = 8'hb7 == _GEN_14503 & _GEN_15783 | _GEN_1210; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3965 = 8'hb7 == _GEN_14503 & _GEN_3591 | _GEN_1722; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3966 = 8'hb8 == _GEN_14503 & _GEN_15783 | _GEN_1211; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3967 = 8'hb8 == _GEN_14503 & _GEN_3591 | _GEN_1723; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3968 = 8'hb9 == _GEN_14503 & _GEN_15783 | _GEN_1212; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3969 = 8'hb9 == _GEN_14503 & _GEN_3591 | _GEN_1724; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3970 = 8'hba == _GEN_14503 & _GEN_15783 | _GEN_1213; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3971 = 8'hba == _GEN_14503 & _GEN_3591 | _GEN_1725; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3972 = 8'hbb == _GEN_14503 & _GEN_15783 | _GEN_1214; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3973 = 8'hbb == _GEN_14503 & _GEN_3591 | _GEN_1726; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3974 = 8'hbc == _GEN_14503 & _GEN_15783 | _GEN_1215; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3975 = 8'hbc == _GEN_14503 & _GEN_3591 | _GEN_1727; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3976 = 8'hbd == _GEN_14503 & _GEN_15783 | _GEN_1216; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3977 = 8'hbd == _GEN_14503 & _GEN_3591 | _GEN_1728; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3978 = 8'hbe == _GEN_14503 & _GEN_15783 | _GEN_1217; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3979 = 8'hbe == _GEN_14503 & _GEN_3591 | _GEN_1729; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3980 = 8'hbf == _GEN_14503 & _GEN_15783 | _GEN_1218; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3981 = 8'hbf == _GEN_14503 & _GEN_3591 | _GEN_1730; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3982 = 8'hc0 == _GEN_14503 & _GEN_15783 | _GEN_1219; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3983 = 8'hc0 == _GEN_14503 & _GEN_3591 | _GEN_1731; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3984 = 8'hc1 == _GEN_14503 & _GEN_15783 | _GEN_1220; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3985 = 8'hc1 == _GEN_14503 & _GEN_3591 | _GEN_1732; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3986 = 8'hc2 == _GEN_14503 & _GEN_15783 | _GEN_1221; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3987 = 8'hc2 == _GEN_14503 & _GEN_3591 | _GEN_1733; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3988 = 8'hc3 == _GEN_14503 & _GEN_15783 | _GEN_1222; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3989 = 8'hc3 == _GEN_14503 & _GEN_3591 | _GEN_1734; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3990 = 8'hc4 == _GEN_14503 & _GEN_15783 | _GEN_1223; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3991 = 8'hc4 == _GEN_14503 & _GEN_3591 | _GEN_1735; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3992 = 8'hc5 == _GEN_14503 & _GEN_15783 | _GEN_1224; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3993 = 8'hc5 == _GEN_14503 & _GEN_3591 | _GEN_1736; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3994 = 8'hc6 == _GEN_14503 & _GEN_15783 | _GEN_1225; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3995 = 8'hc6 == _GEN_14503 & _GEN_3591 | _GEN_1737; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3996 = 8'hc7 == _GEN_14503 & _GEN_15783 | _GEN_1226; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3997 = 8'hc7 == _GEN_14503 & _GEN_3591 | _GEN_1738; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3998 = 8'hc8 == _GEN_14503 & _GEN_15783 | _GEN_1227; // @[ICache.scala 187:{36,36}]
  wire  _GEN_3999 = 8'hc8 == _GEN_14503 & _GEN_3591 | _GEN_1739; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4000 = 8'hc9 == _GEN_14503 & _GEN_15783 | _GEN_1228; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4001 = 8'hc9 == _GEN_14503 & _GEN_3591 | _GEN_1740; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4002 = 8'hca == _GEN_14503 & _GEN_15783 | _GEN_1229; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4003 = 8'hca == _GEN_14503 & _GEN_3591 | _GEN_1741; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4004 = 8'hcb == _GEN_14503 & _GEN_15783 | _GEN_1230; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4005 = 8'hcb == _GEN_14503 & _GEN_3591 | _GEN_1742; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4006 = 8'hcc == _GEN_14503 & _GEN_15783 | _GEN_1231; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4007 = 8'hcc == _GEN_14503 & _GEN_3591 | _GEN_1743; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4008 = 8'hcd == _GEN_14503 & _GEN_15783 | _GEN_1232; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4009 = 8'hcd == _GEN_14503 & _GEN_3591 | _GEN_1744; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4010 = 8'hce == _GEN_14503 & _GEN_15783 | _GEN_1233; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4011 = 8'hce == _GEN_14503 & _GEN_3591 | _GEN_1745; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4012 = 8'hcf == _GEN_14503 & _GEN_15783 | _GEN_1234; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4013 = 8'hcf == _GEN_14503 & _GEN_3591 | _GEN_1746; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4014 = 8'hd0 == _GEN_14503 & _GEN_15783 | _GEN_1235; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4015 = 8'hd0 == _GEN_14503 & _GEN_3591 | _GEN_1747; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4016 = 8'hd1 == _GEN_14503 & _GEN_15783 | _GEN_1236; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4017 = 8'hd1 == _GEN_14503 & _GEN_3591 | _GEN_1748; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4018 = 8'hd2 == _GEN_14503 & _GEN_15783 | _GEN_1237; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4019 = 8'hd2 == _GEN_14503 & _GEN_3591 | _GEN_1749; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4020 = 8'hd3 == _GEN_14503 & _GEN_15783 | _GEN_1238; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4021 = 8'hd3 == _GEN_14503 & _GEN_3591 | _GEN_1750; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4022 = 8'hd4 == _GEN_14503 & _GEN_15783 | _GEN_1239; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4023 = 8'hd4 == _GEN_14503 & _GEN_3591 | _GEN_1751; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4024 = 8'hd5 == _GEN_14503 & _GEN_15783 | _GEN_1240; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4025 = 8'hd5 == _GEN_14503 & _GEN_3591 | _GEN_1752; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4026 = 8'hd6 == _GEN_14503 & _GEN_15783 | _GEN_1241; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4027 = 8'hd6 == _GEN_14503 & _GEN_3591 | _GEN_1753; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4028 = 8'hd7 == _GEN_14503 & _GEN_15783 | _GEN_1242; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4029 = 8'hd7 == _GEN_14503 & _GEN_3591 | _GEN_1754; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4030 = 8'hd8 == _GEN_14503 & _GEN_15783 | _GEN_1243; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4031 = 8'hd8 == _GEN_14503 & _GEN_3591 | _GEN_1755; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4032 = 8'hd9 == _GEN_14503 & _GEN_15783 | _GEN_1244; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4033 = 8'hd9 == _GEN_14503 & _GEN_3591 | _GEN_1756; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4034 = 8'hda == _GEN_14503 & _GEN_15783 | _GEN_1245; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4035 = 8'hda == _GEN_14503 & _GEN_3591 | _GEN_1757; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4036 = 8'hdb == _GEN_14503 & _GEN_15783 | _GEN_1246; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4037 = 8'hdb == _GEN_14503 & _GEN_3591 | _GEN_1758; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4038 = 8'hdc == _GEN_14503 & _GEN_15783 | _GEN_1247; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4039 = 8'hdc == _GEN_14503 & _GEN_3591 | _GEN_1759; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4040 = 8'hdd == _GEN_14503 & _GEN_15783 | _GEN_1248; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4041 = 8'hdd == _GEN_14503 & _GEN_3591 | _GEN_1760; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4042 = 8'hde == _GEN_14503 & _GEN_15783 | _GEN_1249; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4043 = 8'hde == _GEN_14503 & _GEN_3591 | _GEN_1761; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4044 = 8'hdf == _GEN_14503 & _GEN_15783 | _GEN_1250; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4045 = 8'hdf == _GEN_14503 & _GEN_3591 | _GEN_1762; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4046 = 8'he0 == _GEN_14503 & _GEN_15783 | _GEN_1251; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4047 = 8'he0 == _GEN_14503 & _GEN_3591 | _GEN_1763; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4048 = 8'he1 == _GEN_14503 & _GEN_15783 | _GEN_1252; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4049 = 8'he1 == _GEN_14503 & _GEN_3591 | _GEN_1764; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4050 = 8'he2 == _GEN_14503 & _GEN_15783 | _GEN_1253; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4051 = 8'he2 == _GEN_14503 & _GEN_3591 | _GEN_1765; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4052 = 8'he3 == _GEN_14503 & _GEN_15783 | _GEN_1254; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4053 = 8'he3 == _GEN_14503 & _GEN_3591 | _GEN_1766; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4054 = 8'he4 == _GEN_14503 & _GEN_15783 | _GEN_1255; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4055 = 8'he4 == _GEN_14503 & _GEN_3591 | _GEN_1767; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4056 = 8'he5 == _GEN_14503 & _GEN_15783 | _GEN_1256; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4057 = 8'he5 == _GEN_14503 & _GEN_3591 | _GEN_1768; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4058 = 8'he6 == _GEN_14503 & _GEN_15783 | _GEN_1257; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4059 = 8'he6 == _GEN_14503 & _GEN_3591 | _GEN_1769; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4060 = 8'he7 == _GEN_14503 & _GEN_15783 | _GEN_1258; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4061 = 8'he7 == _GEN_14503 & _GEN_3591 | _GEN_1770; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4062 = 8'he8 == _GEN_14503 & _GEN_15783 | _GEN_1259; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4063 = 8'he8 == _GEN_14503 & _GEN_3591 | _GEN_1771; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4064 = 8'he9 == _GEN_14503 & _GEN_15783 | _GEN_1260; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4065 = 8'he9 == _GEN_14503 & _GEN_3591 | _GEN_1772; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4066 = 8'hea == _GEN_14503 & _GEN_15783 | _GEN_1261; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4067 = 8'hea == _GEN_14503 & _GEN_3591 | _GEN_1773; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4068 = 8'heb == _GEN_14503 & _GEN_15783 | _GEN_1262; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4069 = 8'heb == _GEN_14503 & _GEN_3591 | _GEN_1774; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4070 = 8'hec == _GEN_14503 & _GEN_15783 | _GEN_1263; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4071 = 8'hec == _GEN_14503 & _GEN_3591 | _GEN_1775; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4072 = 8'hed == _GEN_14503 & _GEN_15783 | _GEN_1264; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4073 = 8'hed == _GEN_14503 & _GEN_3591 | _GEN_1776; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4074 = 8'hee == _GEN_14503 & _GEN_15783 | _GEN_1265; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4075 = 8'hee == _GEN_14503 & _GEN_3591 | _GEN_1777; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4076 = 8'hef == _GEN_14503 & _GEN_15783 | _GEN_1266; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4077 = 8'hef == _GEN_14503 & _GEN_3591 | _GEN_1778; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4078 = 8'hf0 == _GEN_14503 & _GEN_15783 | _GEN_1267; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4079 = 8'hf0 == _GEN_14503 & _GEN_3591 | _GEN_1779; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4080 = 8'hf1 == _GEN_14503 & _GEN_15783 | _GEN_1268; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4081 = 8'hf1 == _GEN_14503 & _GEN_3591 | _GEN_1780; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4082 = 8'hf2 == _GEN_14503 & _GEN_15783 | _GEN_1269; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4083 = 8'hf2 == _GEN_14503 & _GEN_3591 | _GEN_1781; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4084 = 8'hf3 == _GEN_14503 & _GEN_15783 | _GEN_1270; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4085 = 8'hf3 == _GEN_14503 & _GEN_3591 | _GEN_1782; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4086 = 8'hf4 == _GEN_14503 & _GEN_15783 | _GEN_1271; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4087 = 8'hf4 == _GEN_14503 & _GEN_3591 | _GEN_1783; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4088 = 8'hf5 == _GEN_14503 & _GEN_15783 | _GEN_1272; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4089 = 8'hf5 == _GEN_14503 & _GEN_3591 | _GEN_1784; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4090 = 8'hf6 == _GEN_14503 & _GEN_15783 | _GEN_1273; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4091 = 8'hf6 == _GEN_14503 & _GEN_3591 | _GEN_1785; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4092 = 8'hf7 == _GEN_14503 & _GEN_15783 | _GEN_1274; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4093 = 8'hf7 == _GEN_14503 & _GEN_3591 | _GEN_1786; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4094 = 8'hf8 == _GEN_14503 & _GEN_15783 | _GEN_1275; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4095 = 8'hf8 == _GEN_14503 & _GEN_3591 | _GEN_1787; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4096 = 8'hf9 == _GEN_14503 & _GEN_15783 | _GEN_1276; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4097 = 8'hf9 == _GEN_14503 & _GEN_3591 | _GEN_1788; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4098 = 8'hfa == _GEN_14503 & _GEN_15783 | _GEN_1277; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4099 = 8'hfa == _GEN_14503 & _GEN_3591 | _GEN_1789; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4100 = 8'hfb == _GEN_14503 & _GEN_15783 | _GEN_1278; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4101 = 8'hfb == _GEN_14503 & _GEN_3591 | _GEN_1790; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4102 = 8'hfc == _GEN_14503 & _GEN_15783 | _GEN_1279; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4103 = 8'hfc == _GEN_14503 & _GEN_3591 | _GEN_1791; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4104 = 8'hfd == _GEN_14503 & _GEN_15783 | _GEN_1280; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4105 = 8'hfd == _GEN_14503 & _GEN_3591 | _GEN_1792; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4106 = 8'hfe == _GEN_14503 & _GEN_15783 | _GEN_1281; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4107 = 8'hfe == _GEN_14503 & _GEN_3591 | _GEN_1793; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4108 = 8'hff == _GEN_14503 & _GEN_15783 | _GEN_1282; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4109 = 8'hff == _GEN_14503 & _GEN_3591 | _GEN_1794; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4110 = 9'h100 == _GEN_14631 & _GEN_15783 | _GEN_1283; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4111 = 9'h100 == _GEN_14631 & _GEN_3591 | _GEN_1795; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4112 = 9'h101 == _GEN_14631 & _GEN_15783 | _GEN_1284; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4113 = 9'h101 == _GEN_14631 & _GEN_3591 | _GEN_1796; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4114 = 9'h102 == _GEN_14631 & _GEN_15783 | _GEN_1285; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4115 = 9'h102 == _GEN_14631 & _GEN_3591 | _GEN_1797; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4116 = 9'h103 == _GEN_14631 & _GEN_15783 | _GEN_1286; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4117 = 9'h103 == _GEN_14631 & _GEN_3591 | _GEN_1798; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4118 = 9'h104 == _GEN_14631 & _GEN_15783 | _GEN_1287; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4119 = 9'h104 == _GEN_14631 & _GEN_3591 | _GEN_1799; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4120 = 9'h105 == _GEN_14631 & _GEN_15783 | _GEN_1288; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4121 = 9'h105 == _GEN_14631 & _GEN_3591 | _GEN_1800; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4122 = 9'h106 == _GEN_14631 & _GEN_15783 | _GEN_1289; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4123 = 9'h106 == _GEN_14631 & _GEN_3591 | _GEN_1801; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4124 = 9'h107 == _GEN_14631 & _GEN_15783 | _GEN_1290; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4125 = 9'h107 == _GEN_14631 & _GEN_3591 | _GEN_1802; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4126 = 9'h108 == _GEN_14631 & _GEN_15783 | _GEN_1291; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4127 = 9'h108 == _GEN_14631 & _GEN_3591 | _GEN_1803; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4128 = 9'h109 == _GEN_14631 & _GEN_15783 | _GEN_1292; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4129 = 9'h109 == _GEN_14631 & _GEN_3591 | _GEN_1804; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4130 = 9'h10a == _GEN_14631 & _GEN_15783 | _GEN_1293; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4131 = 9'h10a == _GEN_14631 & _GEN_3591 | _GEN_1805; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4132 = 9'h10b == _GEN_14631 & _GEN_15783 | _GEN_1294; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4133 = 9'h10b == _GEN_14631 & _GEN_3591 | _GEN_1806; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4134 = 9'h10c == _GEN_14631 & _GEN_15783 | _GEN_1295; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4135 = 9'h10c == _GEN_14631 & _GEN_3591 | _GEN_1807; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4136 = 9'h10d == _GEN_14631 & _GEN_15783 | _GEN_1296; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4137 = 9'h10d == _GEN_14631 & _GEN_3591 | _GEN_1808; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4138 = 9'h10e == _GEN_14631 & _GEN_15783 | _GEN_1297; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4139 = 9'h10e == _GEN_14631 & _GEN_3591 | _GEN_1809; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4140 = 9'h10f == _GEN_14631 & _GEN_15783 | _GEN_1298; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4141 = 9'h10f == _GEN_14631 & _GEN_3591 | _GEN_1810; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4142 = 9'h110 == _GEN_14631 & _GEN_15783 | _GEN_1299; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4143 = 9'h110 == _GEN_14631 & _GEN_3591 | _GEN_1811; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4144 = 9'h111 == _GEN_14631 & _GEN_15783 | _GEN_1300; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4145 = 9'h111 == _GEN_14631 & _GEN_3591 | _GEN_1812; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4146 = 9'h112 == _GEN_14631 & _GEN_15783 | _GEN_1301; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4147 = 9'h112 == _GEN_14631 & _GEN_3591 | _GEN_1813; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4148 = 9'h113 == _GEN_14631 & _GEN_15783 | _GEN_1302; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4149 = 9'h113 == _GEN_14631 & _GEN_3591 | _GEN_1814; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4150 = 9'h114 == _GEN_14631 & _GEN_15783 | _GEN_1303; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4151 = 9'h114 == _GEN_14631 & _GEN_3591 | _GEN_1815; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4152 = 9'h115 == _GEN_14631 & _GEN_15783 | _GEN_1304; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4153 = 9'h115 == _GEN_14631 & _GEN_3591 | _GEN_1816; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4154 = 9'h116 == _GEN_14631 & _GEN_15783 | _GEN_1305; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4155 = 9'h116 == _GEN_14631 & _GEN_3591 | _GEN_1817; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4156 = 9'h117 == _GEN_14631 & _GEN_15783 | _GEN_1306; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4157 = 9'h117 == _GEN_14631 & _GEN_3591 | _GEN_1818; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4158 = 9'h118 == _GEN_14631 & _GEN_15783 | _GEN_1307; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4159 = 9'h118 == _GEN_14631 & _GEN_3591 | _GEN_1819; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4160 = 9'h119 == _GEN_14631 & _GEN_15783 | _GEN_1308; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4161 = 9'h119 == _GEN_14631 & _GEN_3591 | _GEN_1820; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4162 = 9'h11a == _GEN_14631 & _GEN_15783 | _GEN_1309; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4163 = 9'h11a == _GEN_14631 & _GEN_3591 | _GEN_1821; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4164 = 9'h11b == _GEN_14631 & _GEN_15783 | _GEN_1310; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4165 = 9'h11b == _GEN_14631 & _GEN_3591 | _GEN_1822; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4166 = 9'h11c == _GEN_14631 & _GEN_15783 | _GEN_1311; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4167 = 9'h11c == _GEN_14631 & _GEN_3591 | _GEN_1823; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4168 = 9'h11d == _GEN_14631 & _GEN_15783 | _GEN_1312; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4169 = 9'h11d == _GEN_14631 & _GEN_3591 | _GEN_1824; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4170 = 9'h11e == _GEN_14631 & _GEN_15783 | _GEN_1313; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4171 = 9'h11e == _GEN_14631 & _GEN_3591 | _GEN_1825; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4172 = 9'h11f == _GEN_14631 & _GEN_15783 | _GEN_1314; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4173 = 9'h11f == _GEN_14631 & _GEN_3591 | _GEN_1826; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4174 = 9'h120 == _GEN_14631 & _GEN_15783 | _GEN_1315; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4175 = 9'h120 == _GEN_14631 & _GEN_3591 | _GEN_1827; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4176 = 9'h121 == _GEN_14631 & _GEN_15783 | _GEN_1316; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4177 = 9'h121 == _GEN_14631 & _GEN_3591 | _GEN_1828; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4178 = 9'h122 == _GEN_14631 & _GEN_15783 | _GEN_1317; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4179 = 9'h122 == _GEN_14631 & _GEN_3591 | _GEN_1829; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4180 = 9'h123 == _GEN_14631 & _GEN_15783 | _GEN_1318; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4181 = 9'h123 == _GEN_14631 & _GEN_3591 | _GEN_1830; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4182 = 9'h124 == _GEN_14631 & _GEN_15783 | _GEN_1319; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4183 = 9'h124 == _GEN_14631 & _GEN_3591 | _GEN_1831; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4184 = 9'h125 == _GEN_14631 & _GEN_15783 | _GEN_1320; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4185 = 9'h125 == _GEN_14631 & _GEN_3591 | _GEN_1832; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4186 = 9'h126 == _GEN_14631 & _GEN_15783 | _GEN_1321; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4187 = 9'h126 == _GEN_14631 & _GEN_3591 | _GEN_1833; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4188 = 9'h127 == _GEN_14631 & _GEN_15783 | _GEN_1322; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4189 = 9'h127 == _GEN_14631 & _GEN_3591 | _GEN_1834; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4190 = 9'h128 == _GEN_14631 & _GEN_15783 | _GEN_1323; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4191 = 9'h128 == _GEN_14631 & _GEN_3591 | _GEN_1835; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4192 = 9'h129 == _GEN_14631 & _GEN_15783 | _GEN_1324; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4193 = 9'h129 == _GEN_14631 & _GEN_3591 | _GEN_1836; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4194 = 9'h12a == _GEN_14631 & _GEN_15783 | _GEN_1325; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4195 = 9'h12a == _GEN_14631 & _GEN_3591 | _GEN_1837; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4196 = 9'h12b == _GEN_14631 & _GEN_15783 | _GEN_1326; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4197 = 9'h12b == _GEN_14631 & _GEN_3591 | _GEN_1838; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4198 = 9'h12c == _GEN_14631 & _GEN_15783 | _GEN_1327; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4199 = 9'h12c == _GEN_14631 & _GEN_3591 | _GEN_1839; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4200 = 9'h12d == _GEN_14631 & _GEN_15783 | _GEN_1328; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4201 = 9'h12d == _GEN_14631 & _GEN_3591 | _GEN_1840; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4202 = 9'h12e == _GEN_14631 & _GEN_15783 | _GEN_1329; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4203 = 9'h12e == _GEN_14631 & _GEN_3591 | _GEN_1841; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4204 = 9'h12f == _GEN_14631 & _GEN_15783 | _GEN_1330; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4205 = 9'h12f == _GEN_14631 & _GEN_3591 | _GEN_1842; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4206 = 9'h130 == _GEN_14631 & _GEN_15783 | _GEN_1331; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4207 = 9'h130 == _GEN_14631 & _GEN_3591 | _GEN_1843; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4208 = 9'h131 == _GEN_14631 & _GEN_15783 | _GEN_1332; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4209 = 9'h131 == _GEN_14631 & _GEN_3591 | _GEN_1844; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4210 = 9'h132 == _GEN_14631 & _GEN_15783 | _GEN_1333; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4211 = 9'h132 == _GEN_14631 & _GEN_3591 | _GEN_1845; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4212 = 9'h133 == _GEN_14631 & _GEN_15783 | _GEN_1334; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4213 = 9'h133 == _GEN_14631 & _GEN_3591 | _GEN_1846; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4214 = 9'h134 == _GEN_14631 & _GEN_15783 | _GEN_1335; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4215 = 9'h134 == _GEN_14631 & _GEN_3591 | _GEN_1847; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4216 = 9'h135 == _GEN_14631 & _GEN_15783 | _GEN_1336; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4217 = 9'h135 == _GEN_14631 & _GEN_3591 | _GEN_1848; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4218 = 9'h136 == _GEN_14631 & _GEN_15783 | _GEN_1337; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4219 = 9'h136 == _GEN_14631 & _GEN_3591 | _GEN_1849; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4220 = 9'h137 == _GEN_14631 & _GEN_15783 | _GEN_1338; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4221 = 9'h137 == _GEN_14631 & _GEN_3591 | _GEN_1850; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4222 = 9'h138 == _GEN_14631 & _GEN_15783 | _GEN_1339; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4223 = 9'h138 == _GEN_14631 & _GEN_3591 | _GEN_1851; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4224 = 9'h139 == _GEN_14631 & _GEN_15783 | _GEN_1340; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4225 = 9'h139 == _GEN_14631 & _GEN_3591 | _GEN_1852; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4226 = 9'h13a == _GEN_14631 & _GEN_15783 | _GEN_1341; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4227 = 9'h13a == _GEN_14631 & _GEN_3591 | _GEN_1853; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4228 = 9'h13b == _GEN_14631 & _GEN_15783 | _GEN_1342; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4229 = 9'h13b == _GEN_14631 & _GEN_3591 | _GEN_1854; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4230 = 9'h13c == _GEN_14631 & _GEN_15783 | _GEN_1343; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4231 = 9'h13c == _GEN_14631 & _GEN_3591 | _GEN_1855; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4232 = 9'h13d == _GEN_14631 & _GEN_15783 | _GEN_1344; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4233 = 9'h13d == _GEN_14631 & _GEN_3591 | _GEN_1856; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4234 = 9'h13e == _GEN_14631 & _GEN_15783 | _GEN_1345; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4235 = 9'h13e == _GEN_14631 & _GEN_3591 | _GEN_1857; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4236 = 9'h13f == _GEN_14631 & _GEN_15783 | _GEN_1346; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4237 = 9'h13f == _GEN_14631 & _GEN_3591 | _GEN_1858; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4238 = 9'h140 == _GEN_14631 & _GEN_15783 | _GEN_1347; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4239 = 9'h140 == _GEN_14631 & _GEN_3591 | _GEN_1859; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4240 = 9'h141 == _GEN_14631 & _GEN_15783 | _GEN_1348; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4241 = 9'h141 == _GEN_14631 & _GEN_3591 | _GEN_1860; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4242 = 9'h142 == _GEN_14631 & _GEN_15783 | _GEN_1349; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4243 = 9'h142 == _GEN_14631 & _GEN_3591 | _GEN_1861; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4244 = 9'h143 == _GEN_14631 & _GEN_15783 | _GEN_1350; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4245 = 9'h143 == _GEN_14631 & _GEN_3591 | _GEN_1862; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4246 = 9'h144 == _GEN_14631 & _GEN_15783 | _GEN_1351; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4247 = 9'h144 == _GEN_14631 & _GEN_3591 | _GEN_1863; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4248 = 9'h145 == _GEN_14631 & _GEN_15783 | _GEN_1352; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4249 = 9'h145 == _GEN_14631 & _GEN_3591 | _GEN_1864; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4250 = 9'h146 == _GEN_14631 & _GEN_15783 | _GEN_1353; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4251 = 9'h146 == _GEN_14631 & _GEN_3591 | _GEN_1865; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4252 = 9'h147 == _GEN_14631 & _GEN_15783 | _GEN_1354; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4253 = 9'h147 == _GEN_14631 & _GEN_3591 | _GEN_1866; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4254 = 9'h148 == _GEN_14631 & _GEN_15783 | _GEN_1355; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4255 = 9'h148 == _GEN_14631 & _GEN_3591 | _GEN_1867; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4256 = 9'h149 == _GEN_14631 & _GEN_15783 | _GEN_1356; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4257 = 9'h149 == _GEN_14631 & _GEN_3591 | _GEN_1868; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4258 = 9'h14a == _GEN_14631 & _GEN_15783 | _GEN_1357; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4259 = 9'h14a == _GEN_14631 & _GEN_3591 | _GEN_1869; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4260 = 9'h14b == _GEN_14631 & _GEN_15783 | _GEN_1358; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4261 = 9'h14b == _GEN_14631 & _GEN_3591 | _GEN_1870; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4262 = 9'h14c == _GEN_14631 & _GEN_15783 | _GEN_1359; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4263 = 9'h14c == _GEN_14631 & _GEN_3591 | _GEN_1871; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4264 = 9'h14d == _GEN_14631 & _GEN_15783 | _GEN_1360; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4265 = 9'h14d == _GEN_14631 & _GEN_3591 | _GEN_1872; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4266 = 9'h14e == _GEN_14631 & _GEN_15783 | _GEN_1361; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4267 = 9'h14e == _GEN_14631 & _GEN_3591 | _GEN_1873; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4268 = 9'h14f == _GEN_14631 & _GEN_15783 | _GEN_1362; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4269 = 9'h14f == _GEN_14631 & _GEN_3591 | _GEN_1874; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4270 = 9'h150 == _GEN_14631 & _GEN_15783 | _GEN_1363; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4271 = 9'h150 == _GEN_14631 & _GEN_3591 | _GEN_1875; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4272 = 9'h151 == _GEN_14631 & _GEN_15783 | _GEN_1364; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4273 = 9'h151 == _GEN_14631 & _GEN_3591 | _GEN_1876; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4274 = 9'h152 == _GEN_14631 & _GEN_15783 | _GEN_1365; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4275 = 9'h152 == _GEN_14631 & _GEN_3591 | _GEN_1877; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4276 = 9'h153 == _GEN_14631 & _GEN_15783 | _GEN_1366; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4277 = 9'h153 == _GEN_14631 & _GEN_3591 | _GEN_1878; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4278 = 9'h154 == _GEN_14631 & _GEN_15783 | _GEN_1367; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4279 = 9'h154 == _GEN_14631 & _GEN_3591 | _GEN_1879; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4280 = 9'h155 == _GEN_14631 & _GEN_15783 | _GEN_1368; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4281 = 9'h155 == _GEN_14631 & _GEN_3591 | _GEN_1880; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4282 = 9'h156 == _GEN_14631 & _GEN_15783 | _GEN_1369; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4283 = 9'h156 == _GEN_14631 & _GEN_3591 | _GEN_1881; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4284 = 9'h157 == _GEN_14631 & _GEN_15783 | _GEN_1370; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4285 = 9'h157 == _GEN_14631 & _GEN_3591 | _GEN_1882; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4286 = 9'h158 == _GEN_14631 & _GEN_15783 | _GEN_1371; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4287 = 9'h158 == _GEN_14631 & _GEN_3591 | _GEN_1883; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4288 = 9'h159 == _GEN_14631 & _GEN_15783 | _GEN_1372; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4289 = 9'h159 == _GEN_14631 & _GEN_3591 | _GEN_1884; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4290 = 9'h15a == _GEN_14631 & _GEN_15783 | _GEN_1373; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4291 = 9'h15a == _GEN_14631 & _GEN_3591 | _GEN_1885; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4292 = 9'h15b == _GEN_14631 & _GEN_15783 | _GEN_1374; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4293 = 9'h15b == _GEN_14631 & _GEN_3591 | _GEN_1886; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4294 = 9'h15c == _GEN_14631 & _GEN_15783 | _GEN_1375; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4295 = 9'h15c == _GEN_14631 & _GEN_3591 | _GEN_1887; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4296 = 9'h15d == _GEN_14631 & _GEN_15783 | _GEN_1376; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4297 = 9'h15d == _GEN_14631 & _GEN_3591 | _GEN_1888; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4298 = 9'h15e == _GEN_14631 & _GEN_15783 | _GEN_1377; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4299 = 9'h15e == _GEN_14631 & _GEN_3591 | _GEN_1889; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4300 = 9'h15f == _GEN_14631 & _GEN_15783 | _GEN_1378; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4301 = 9'h15f == _GEN_14631 & _GEN_3591 | _GEN_1890; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4302 = 9'h160 == _GEN_14631 & _GEN_15783 | _GEN_1379; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4303 = 9'h160 == _GEN_14631 & _GEN_3591 | _GEN_1891; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4304 = 9'h161 == _GEN_14631 & _GEN_15783 | _GEN_1380; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4305 = 9'h161 == _GEN_14631 & _GEN_3591 | _GEN_1892; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4306 = 9'h162 == _GEN_14631 & _GEN_15783 | _GEN_1381; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4307 = 9'h162 == _GEN_14631 & _GEN_3591 | _GEN_1893; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4308 = 9'h163 == _GEN_14631 & _GEN_15783 | _GEN_1382; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4309 = 9'h163 == _GEN_14631 & _GEN_3591 | _GEN_1894; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4310 = 9'h164 == _GEN_14631 & _GEN_15783 | _GEN_1383; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4311 = 9'h164 == _GEN_14631 & _GEN_3591 | _GEN_1895; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4312 = 9'h165 == _GEN_14631 & _GEN_15783 | _GEN_1384; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4313 = 9'h165 == _GEN_14631 & _GEN_3591 | _GEN_1896; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4314 = 9'h166 == _GEN_14631 & _GEN_15783 | _GEN_1385; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4315 = 9'h166 == _GEN_14631 & _GEN_3591 | _GEN_1897; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4316 = 9'h167 == _GEN_14631 & _GEN_15783 | _GEN_1386; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4317 = 9'h167 == _GEN_14631 & _GEN_3591 | _GEN_1898; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4318 = 9'h168 == _GEN_14631 & _GEN_15783 | _GEN_1387; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4319 = 9'h168 == _GEN_14631 & _GEN_3591 | _GEN_1899; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4320 = 9'h169 == _GEN_14631 & _GEN_15783 | _GEN_1388; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4321 = 9'h169 == _GEN_14631 & _GEN_3591 | _GEN_1900; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4322 = 9'h16a == _GEN_14631 & _GEN_15783 | _GEN_1389; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4323 = 9'h16a == _GEN_14631 & _GEN_3591 | _GEN_1901; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4324 = 9'h16b == _GEN_14631 & _GEN_15783 | _GEN_1390; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4325 = 9'h16b == _GEN_14631 & _GEN_3591 | _GEN_1902; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4326 = 9'h16c == _GEN_14631 & _GEN_15783 | _GEN_1391; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4327 = 9'h16c == _GEN_14631 & _GEN_3591 | _GEN_1903; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4328 = 9'h16d == _GEN_14631 & _GEN_15783 | _GEN_1392; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4329 = 9'h16d == _GEN_14631 & _GEN_3591 | _GEN_1904; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4330 = 9'h16e == _GEN_14631 & _GEN_15783 | _GEN_1393; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4331 = 9'h16e == _GEN_14631 & _GEN_3591 | _GEN_1905; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4332 = 9'h16f == _GEN_14631 & _GEN_15783 | _GEN_1394; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4333 = 9'h16f == _GEN_14631 & _GEN_3591 | _GEN_1906; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4334 = 9'h170 == _GEN_14631 & _GEN_15783 | _GEN_1395; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4335 = 9'h170 == _GEN_14631 & _GEN_3591 | _GEN_1907; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4336 = 9'h171 == _GEN_14631 & _GEN_15783 | _GEN_1396; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4337 = 9'h171 == _GEN_14631 & _GEN_3591 | _GEN_1908; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4338 = 9'h172 == _GEN_14631 & _GEN_15783 | _GEN_1397; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4339 = 9'h172 == _GEN_14631 & _GEN_3591 | _GEN_1909; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4340 = 9'h173 == _GEN_14631 & _GEN_15783 | _GEN_1398; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4341 = 9'h173 == _GEN_14631 & _GEN_3591 | _GEN_1910; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4342 = 9'h174 == _GEN_14631 & _GEN_15783 | _GEN_1399; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4343 = 9'h174 == _GEN_14631 & _GEN_3591 | _GEN_1911; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4344 = 9'h175 == _GEN_14631 & _GEN_15783 | _GEN_1400; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4345 = 9'h175 == _GEN_14631 & _GEN_3591 | _GEN_1912; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4346 = 9'h176 == _GEN_14631 & _GEN_15783 | _GEN_1401; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4347 = 9'h176 == _GEN_14631 & _GEN_3591 | _GEN_1913; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4348 = 9'h177 == _GEN_14631 & _GEN_15783 | _GEN_1402; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4349 = 9'h177 == _GEN_14631 & _GEN_3591 | _GEN_1914; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4350 = 9'h178 == _GEN_14631 & _GEN_15783 | _GEN_1403; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4351 = 9'h178 == _GEN_14631 & _GEN_3591 | _GEN_1915; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4352 = 9'h179 == _GEN_14631 & _GEN_15783 | _GEN_1404; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4353 = 9'h179 == _GEN_14631 & _GEN_3591 | _GEN_1916; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4354 = 9'h17a == _GEN_14631 & _GEN_15783 | _GEN_1405; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4355 = 9'h17a == _GEN_14631 & _GEN_3591 | _GEN_1917; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4356 = 9'h17b == _GEN_14631 & _GEN_15783 | _GEN_1406; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4357 = 9'h17b == _GEN_14631 & _GEN_3591 | _GEN_1918; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4358 = 9'h17c == _GEN_14631 & _GEN_15783 | _GEN_1407; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4359 = 9'h17c == _GEN_14631 & _GEN_3591 | _GEN_1919; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4360 = 9'h17d == _GEN_14631 & _GEN_15783 | _GEN_1408; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4361 = 9'h17d == _GEN_14631 & _GEN_3591 | _GEN_1920; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4362 = 9'h17e == _GEN_14631 & _GEN_15783 | _GEN_1409; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4363 = 9'h17e == _GEN_14631 & _GEN_3591 | _GEN_1921; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4364 = 9'h17f == _GEN_14631 & _GEN_15783 | _GEN_1410; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4365 = 9'h17f == _GEN_14631 & _GEN_3591 | _GEN_1922; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4366 = 9'h180 == _GEN_14631 & _GEN_15783 | _GEN_1411; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4367 = 9'h180 == _GEN_14631 & _GEN_3591 | _GEN_1923; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4368 = 9'h181 == _GEN_14631 & _GEN_15783 | _GEN_1412; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4369 = 9'h181 == _GEN_14631 & _GEN_3591 | _GEN_1924; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4370 = 9'h182 == _GEN_14631 & _GEN_15783 | _GEN_1413; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4371 = 9'h182 == _GEN_14631 & _GEN_3591 | _GEN_1925; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4372 = 9'h183 == _GEN_14631 & _GEN_15783 | _GEN_1414; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4373 = 9'h183 == _GEN_14631 & _GEN_3591 | _GEN_1926; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4374 = 9'h184 == _GEN_14631 & _GEN_15783 | _GEN_1415; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4375 = 9'h184 == _GEN_14631 & _GEN_3591 | _GEN_1927; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4376 = 9'h185 == _GEN_14631 & _GEN_15783 | _GEN_1416; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4377 = 9'h185 == _GEN_14631 & _GEN_3591 | _GEN_1928; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4378 = 9'h186 == _GEN_14631 & _GEN_15783 | _GEN_1417; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4379 = 9'h186 == _GEN_14631 & _GEN_3591 | _GEN_1929; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4380 = 9'h187 == _GEN_14631 & _GEN_15783 | _GEN_1418; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4381 = 9'h187 == _GEN_14631 & _GEN_3591 | _GEN_1930; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4382 = 9'h188 == _GEN_14631 & _GEN_15783 | _GEN_1419; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4383 = 9'h188 == _GEN_14631 & _GEN_3591 | _GEN_1931; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4384 = 9'h189 == _GEN_14631 & _GEN_15783 | _GEN_1420; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4385 = 9'h189 == _GEN_14631 & _GEN_3591 | _GEN_1932; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4386 = 9'h18a == _GEN_14631 & _GEN_15783 | _GEN_1421; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4387 = 9'h18a == _GEN_14631 & _GEN_3591 | _GEN_1933; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4388 = 9'h18b == _GEN_14631 & _GEN_15783 | _GEN_1422; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4389 = 9'h18b == _GEN_14631 & _GEN_3591 | _GEN_1934; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4390 = 9'h18c == _GEN_14631 & _GEN_15783 | _GEN_1423; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4391 = 9'h18c == _GEN_14631 & _GEN_3591 | _GEN_1935; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4392 = 9'h18d == _GEN_14631 & _GEN_15783 | _GEN_1424; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4393 = 9'h18d == _GEN_14631 & _GEN_3591 | _GEN_1936; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4394 = 9'h18e == _GEN_14631 & _GEN_15783 | _GEN_1425; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4395 = 9'h18e == _GEN_14631 & _GEN_3591 | _GEN_1937; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4396 = 9'h18f == _GEN_14631 & _GEN_15783 | _GEN_1426; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4397 = 9'h18f == _GEN_14631 & _GEN_3591 | _GEN_1938; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4398 = 9'h190 == _GEN_14631 & _GEN_15783 | _GEN_1427; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4399 = 9'h190 == _GEN_14631 & _GEN_3591 | _GEN_1939; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4400 = 9'h191 == _GEN_14631 & _GEN_15783 | _GEN_1428; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4401 = 9'h191 == _GEN_14631 & _GEN_3591 | _GEN_1940; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4402 = 9'h192 == _GEN_14631 & _GEN_15783 | _GEN_1429; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4403 = 9'h192 == _GEN_14631 & _GEN_3591 | _GEN_1941; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4404 = 9'h193 == _GEN_14631 & _GEN_15783 | _GEN_1430; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4405 = 9'h193 == _GEN_14631 & _GEN_3591 | _GEN_1942; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4406 = 9'h194 == _GEN_14631 & _GEN_15783 | _GEN_1431; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4407 = 9'h194 == _GEN_14631 & _GEN_3591 | _GEN_1943; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4408 = 9'h195 == _GEN_14631 & _GEN_15783 | _GEN_1432; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4409 = 9'h195 == _GEN_14631 & _GEN_3591 | _GEN_1944; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4410 = 9'h196 == _GEN_14631 & _GEN_15783 | _GEN_1433; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4411 = 9'h196 == _GEN_14631 & _GEN_3591 | _GEN_1945; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4412 = 9'h197 == _GEN_14631 & _GEN_15783 | _GEN_1434; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4413 = 9'h197 == _GEN_14631 & _GEN_3591 | _GEN_1946; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4414 = 9'h198 == _GEN_14631 & _GEN_15783 | _GEN_1435; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4415 = 9'h198 == _GEN_14631 & _GEN_3591 | _GEN_1947; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4416 = 9'h199 == _GEN_14631 & _GEN_15783 | _GEN_1436; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4417 = 9'h199 == _GEN_14631 & _GEN_3591 | _GEN_1948; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4418 = 9'h19a == _GEN_14631 & _GEN_15783 | _GEN_1437; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4419 = 9'h19a == _GEN_14631 & _GEN_3591 | _GEN_1949; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4420 = 9'h19b == _GEN_14631 & _GEN_15783 | _GEN_1438; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4421 = 9'h19b == _GEN_14631 & _GEN_3591 | _GEN_1950; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4422 = 9'h19c == _GEN_14631 & _GEN_15783 | _GEN_1439; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4423 = 9'h19c == _GEN_14631 & _GEN_3591 | _GEN_1951; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4424 = 9'h19d == _GEN_14631 & _GEN_15783 | _GEN_1440; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4425 = 9'h19d == _GEN_14631 & _GEN_3591 | _GEN_1952; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4426 = 9'h19e == _GEN_14631 & _GEN_15783 | _GEN_1441; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4427 = 9'h19e == _GEN_14631 & _GEN_3591 | _GEN_1953; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4428 = 9'h19f == _GEN_14631 & _GEN_15783 | _GEN_1442; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4429 = 9'h19f == _GEN_14631 & _GEN_3591 | _GEN_1954; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4430 = 9'h1a0 == _GEN_14631 & _GEN_15783 | _GEN_1443; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4431 = 9'h1a0 == _GEN_14631 & _GEN_3591 | _GEN_1955; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4432 = 9'h1a1 == _GEN_14631 & _GEN_15783 | _GEN_1444; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4433 = 9'h1a1 == _GEN_14631 & _GEN_3591 | _GEN_1956; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4434 = 9'h1a2 == _GEN_14631 & _GEN_15783 | _GEN_1445; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4435 = 9'h1a2 == _GEN_14631 & _GEN_3591 | _GEN_1957; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4436 = 9'h1a3 == _GEN_14631 & _GEN_15783 | _GEN_1446; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4437 = 9'h1a3 == _GEN_14631 & _GEN_3591 | _GEN_1958; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4438 = 9'h1a4 == _GEN_14631 & _GEN_15783 | _GEN_1447; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4439 = 9'h1a4 == _GEN_14631 & _GEN_3591 | _GEN_1959; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4440 = 9'h1a5 == _GEN_14631 & _GEN_15783 | _GEN_1448; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4441 = 9'h1a5 == _GEN_14631 & _GEN_3591 | _GEN_1960; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4442 = 9'h1a6 == _GEN_14631 & _GEN_15783 | _GEN_1449; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4443 = 9'h1a6 == _GEN_14631 & _GEN_3591 | _GEN_1961; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4444 = 9'h1a7 == _GEN_14631 & _GEN_15783 | _GEN_1450; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4445 = 9'h1a7 == _GEN_14631 & _GEN_3591 | _GEN_1962; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4446 = 9'h1a8 == _GEN_14631 & _GEN_15783 | _GEN_1451; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4447 = 9'h1a8 == _GEN_14631 & _GEN_3591 | _GEN_1963; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4448 = 9'h1a9 == _GEN_14631 & _GEN_15783 | _GEN_1452; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4449 = 9'h1a9 == _GEN_14631 & _GEN_3591 | _GEN_1964; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4450 = 9'h1aa == _GEN_14631 & _GEN_15783 | _GEN_1453; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4451 = 9'h1aa == _GEN_14631 & _GEN_3591 | _GEN_1965; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4452 = 9'h1ab == _GEN_14631 & _GEN_15783 | _GEN_1454; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4453 = 9'h1ab == _GEN_14631 & _GEN_3591 | _GEN_1966; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4454 = 9'h1ac == _GEN_14631 & _GEN_15783 | _GEN_1455; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4455 = 9'h1ac == _GEN_14631 & _GEN_3591 | _GEN_1967; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4456 = 9'h1ad == _GEN_14631 & _GEN_15783 | _GEN_1456; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4457 = 9'h1ad == _GEN_14631 & _GEN_3591 | _GEN_1968; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4458 = 9'h1ae == _GEN_14631 & _GEN_15783 | _GEN_1457; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4459 = 9'h1ae == _GEN_14631 & _GEN_3591 | _GEN_1969; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4460 = 9'h1af == _GEN_14631 & _GEN_15783 | _GEN_1458; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4461 = 9'h1af == _GEN_14631 & _GEN_3591 | _GEN_1970; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4462 = 9'h1b0 == _GEN_14631 & _GEN_15783 | _GEN_1459; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4463 = 9'h1b0 == _GEN_14631 & _GEN_3591 | _GEN_1971; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4464 = 9'h1b1 == _GEN_14631 & _GEN_15783 | _GEN_1460; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4465 = 9'h1b1 == _GEN_14631 & _GEN_3591 | _GEN_1972; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4466 = 9'h1b2 == _GEN_14631 & _GEN_15783 | _GEN_1461; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4467 = 9'h1b2 == _GEN_14631 & _GEN_3591 | _GEN_1973; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4468 = 9'h1b3 == _GEN_14631 & _GEN_15783 | _GEN_1462; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4469 = 9'h1b3 == _GEN_14631 & _GEN_3591 | _GEN_1974; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4470 = 9'h1b4 == _GEN_14631 & _GEN_15783 | _GEN_1463; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4471 = 9'h1b4 == _GEN_14631 & _GEN_3591 | _GEN_1975; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4472 = 9'h1b5 == _GEN_14631 & _GEN_15783 | _GEN_1464; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4473 = 9'h1b5 == _GEN_14631 & _GEN_3591 | _GEN_1976; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4474 = 9'h1b6 == _GEN_14631 & _GEN_15783 | _GEN_1465; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4475 = 9'h1b6 == _GEN_14631 & _GEN_3591 | _GEN_1977; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4476 = 9'h1b7 == _GEN_14631 & _GEN_15783 | _GEN_1466; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4477 = 9'h1b7 == _GEN_14631 & _GEN_3591 | _GEN_1978; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4478 = 9'h1b8 == _GEN_14631 & _GEN_15783 | _GEN_1467; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4479 = 9'h1b8 == _GEN_14631 & _GEN_3591 | _GEN_1979; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4480 = 9'h1b9 == _GEN_14631 & _GEN_15783 | _GEN_1468; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4481 = 9'h1b9 == _GEN_14631 & _GEN_3591 | _GEN_1980; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4482 = 9'h1ba == _GEN_14631 & _GEN_15783 | _GEN_1469; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4483 = 9'h1ba == _GEN_14631 & _GEN_3591 | _GEN_1981; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4484 = 9'h1bb == _GEN_14631 & _GEN_15783 | _GEN_1470; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4485 = 9'h1bb == _GEN_14631 & _GEN_3591 | _GEN_1982; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4486 = 9'h1bc == _GEN_14631 & _GEN_15783 | _GEN_1471; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4487 = 9'h1bc == _GEN_14631 & _GEN_3591 | _GEN_1983; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4488 = 9'h1bd == _GEN_14631 & _GEN_15783 | _GEN_1472; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4489 = 9'h1bd == _GEN_14631 & _GEN_3591 | _GEN_1984; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4490 = 9'h1be == _GEN_14631 & _GEN_15783 | _GEN_1473; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4491 = 9'h1be == _GEN_14631 & _GEN_3591 | _GEN_1985; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4492 = 9'h1bf == _GEN_14631 & _GEN_15783 | _GEN_1474; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4493 = 9'h1bf == _GEN_14631 & _GEN_3591 | _GEN_1986; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4494 = 9'h1c0 == _GEN_14631 & _GEN_15783 | _GEN_1475; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4495 = 9'h1c0 == _GEN_14631 & _GEN_3591 | _GEN_1987; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4496 = 9'h1c1 == _GEN_14631 & _GEN_15783 | _GEN_1476; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4497 = 9'h1c1 == _GEN_14631 & _GEN_3591 | _GEN_1988; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4498 = 9'h1c2 == _GEN_14631 & _GEN_15783 | _GEN_1477; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4499 = 9'h1c2 == _GEN_14631 & _GEN_3591 | _GEN_1989; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4500 = 9'h1c3 == _GEN_14631 & _GEN_15783 | _GEN_1478; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4501 = 9'h1c3 == _GEN_14631 & _GEN_3591 | _GEN_1990; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4502 = 9'h1c4 == _GEN_14631 & _GEN_15783 | _GEN_1479; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4503 = 9'h1c4 == _GEN_14631 & _GEN_3591 | _GEN_1991; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4504 = 9'h1c5 == _GEN_14631 & _GEN_15783 | _GEN_1480; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4505 = 9'h1c5 == _GEN_14631 & _GEN_3591 | _GEN_1992; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4506 = 9'h1c6 == _GEN_14631 & _GEN_15783 | _GEN_1481; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4507 = 9'h1c6 == _GEN_14631 & _GEN_3591 | _GEN_1993; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4508 = 9'h1c7 == _GEN_14631 & _GEN_15783 | _GEN_1482; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4509 = 9'h1c7 == _GEN_14631 & _GEN_3591 | _GEN_1994; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4510 = 9'h1c8 == _GEN_14631 & _GEN_15783 | _GEN_1483; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4511 = 9'h1c8 == _GEN_14631 & _GEN_3591 | _GEN_1995; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4512 = 9'h1c9 == _GEN_14631 & _GEN_15783 | _GEN_1484; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4513 = 9'h1c9 == _GEN_14631 & _GEN_3591 | _GEN_1996; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4514 = 9'h1ca == _GEN_14631 & _GEN_15783 | _GEN_1485; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4515 = 9'h1ca == _GEN_14631 & _GEN_3591 | _GEN_1997; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4516 = 9'h1cb == _GEN_14631 & _GEN_15783 | _GEN_1486; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4517 = 9'h1cb == _GEN_14631 & _GEN_3591 | _GEN_1998; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4518 = 9'h1cc == _GEN_14631 & _GEN_15783 | _GEN_1487; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4519 = 9'h1cc == _GEN_14631 & _GEN_3591 | _GEN_1999; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4520 = 9'h1cd == _GEN_14631 & _GEN_15783 | _GEN_1488; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4521 = 9'h1cd == _GEN_14631 & _GEN_3591 | _GEN_2000; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4522 = 9'h1ce == _GEN_14631 & _GEN_15783 | _GEN_1489; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4523 = 9'h1ce == _GEN_14631 & _GEN_3591 | _GEN_2001; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4524 = 9'h1cf == _GEN_14631 & _GEN_15783 | _GEN_1490; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4525 = 9'h1cf == _GEN_14631 & _GEN_3591 | _GEN_2002; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4526 = 9'h1d0 == _GEN_14631 & _GEN_15783 | _GEN_1491; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4527 = 9'h1d0 == _GEN_14631 & _GEN_3591 | _GEN_2003; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4528 = 9'h1d1 == _GEN_14631 & _GEN_15783 | _GEN_1492; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4529 = 9'h1d1 == _GEN_14631 & _GEN_3591 | _GEN_2004; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4530 = 9'h1d2 == _GEN_14631 & _GEN_15783 | _GEN_1493; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4531 = 9'h1d2 == _GEN_14631 & _GEN_3591 | _GEN_2005; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4532 = 9'h1d3 == _GEN_14631 & _GEN_15783 | _GEN_1494; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4533 = 9'h1d3 == _GEN_14631 & _GEN_3591 | _GEN_2006; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4534 = 9'h1d4 == _GEN_14631 & _GEN_15783 | _GEN_1495; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4535 = 9'h1d4 == _GEN_14631 & _GEN_3591 | _GEN_2007; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4536 = 9'h1d5 == _GEN_14631 & _GEN_15783 | _GEN_1496; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4537 = 9'h1d5 == _GEN_14631 & _GEN_3591 | _GEN_2008; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4538 = 9'h1d6 == _GEN_14631 & _GEN_15783 | _GEN_1497; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4539 = 9'h1d6 == _GEN_14631 & _GEN_3591 | _GEN_2009; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4540 = 9'h1d7 == _GEN_14631 & _GEN_15783 | _GEN_1498; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4541 = 9'h1d7 == _GEN_14631 & _GEN_3591 | _GEN_2010; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4542 = 9'h1d8 == _GEN_14631 & _GEN_15783 | _GEN_1499; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4543 = 9'h1d8 == _GEN_14631 & _GEN_3591 | _GEN_2011; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4544 = 9'h1d9 == _GEN_14631 & _GEN_15783 | _GEN_1500; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4545 = 9'h1d9 == _GEN_14631 & _GEN_3591 | _GEN_2012; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4546 = 9'h1da == _GEN_14631 & _GEN_15783 | _GEN_1501; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4547 = 9'h1da == _GEN_14631 & _GEN_3591 | _GEN_2013; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4548 = 9'h1db == _GEN_14631 & _GEN_15783 | _GEN_1502; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4549 = 9'h1db == _GEN_14631 & _GEN_3591 | _GEN_2014; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4550 = 9'h1dc == _GEN_14631 & _GEN_15783 | _GEN_1503; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4551 = 9'h1dc == _GEN_14631 & _GEN_3591 | _GEN_2015; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4552 = 9'h1dd == _GEN_14631 & _GEN_15783 | _GEN_1504; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4553 = 9'h1dd == _GEN_14631 & _GEN_3591 | _GEN_2016; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4554 = 9'h1de == _GEN_14631 & _GEN_15783 | _GEN_1505; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4555 = 9'h1de == _GEN_14631 & _GEN_3591 | _GEN_2017; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4556 = 9'h1df == _GEN_14631 & _GEN_15783 | _GEN_1506; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4557 = 9'h1df == _GEN_14631 & _GEN_3591 | _GEN_2018; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4558 = 9'h1e0 == _GEN_14631 & _GEN_15783 | _GEN_1507; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4559 = 9'h1e0 == _GEN_14631 & _GEN_3591 | _GEN_2019; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4560 = 9'h1e1 == _GEN_14631 & _GEN_15783 | _GEN_1508; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4561 = 9'h1e1 == _GEN_14631 & _GEN_3591 | _GEN_2020; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4562 = 9'h1e2 == _GEN_14631 & _GEN_15783 | _GEN_1509; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4563 = 9'h1e2 == _GEN_14631 & _GEN_3591 | _GEN_2021; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4564 = 9'h1e3 == _GEN_14631 & _GEN_15783 | _GEN_1510; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4565 = 9'h1e3 == _GEN_14631 & _GEN_3591 | _GEN_2022; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4566 = 9'h1e4 == _GEN_14631 & _GEN_15783 | _GEN_1511; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4567 = 9'h1e4 == _GEN_14631 & _GEN_3591 | _GEN_2023; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4568 = 9'h1e5 == _GEN_14631 & _GEN_15783 | _GEN_1512; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4569 = 9'h1e5 == _GEN_14631 & _GEN_3591 | _GEN_2024; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4570 = 9'h1e6 == _GEN_14631 & _GEN_15783 | _GEN_1513; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4571 = 9'h1e6 == _GEN_14631 & _GEN_3591 | _GEN_2025; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4572 = 9'h1e7 == _GEN_14631 & _GEN_15783 | _GEN_1514; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4573 = 9'h1e7 == _GEN_14631 & _GEN_3591 | _GEN_2026; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4574 = 9'h1e8 == _GEN_14631 & _GEN_15783 | _GEN_1515; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4575 = 9'h1e8 == _GEN_14631 & _GEN_3591 | _GEN_2027; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4576 = 9'h1e9 == _GEN_14631 & _GEN_15783 | _GEN_1516; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4577 = 9'h1e9 == _GEN_14631 & _GEN_3591 | _GEN_2028; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4578 = 9'h1ea == _GEN_14631 & _GEN_15783 | _GEN_1517; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4579 = 9'h1ea == _GEN_14631 & _GEN_3591 | _GEN_2029; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4580 = 9'h1eb == _GEN_14631 & _GEN_15783 | _GEN_1518; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4581 = 9'h1eb == _GEN_14631 & _GEN_3591 | _GEN_2030; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4582 = 9'h1ec == _GEN_14631 & _GEN_15783 | _GEN_1519; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4583 = 9'h1ec == _GEN_14631 & _GEN_3591 | _GEN_2031; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4584 = 9'h1ed == _GEN_14631 & _GEN_15783 | _GEN_1520; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4585 = 9'h1ed == _GEN_14631 & _GEN_3591 | _GEN_2032; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4586 = 9'h1ee == _GEN_14631 & _GEN_15783 | _GEN_1521; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4587 = 9'h1ee == _GEN_14631 & _GEN_3591 | _GEN_2033; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4588 = 9'h1ef == _GEN_14631 & _GEN_15783 | _GEN_1522; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4589 = 9'h1ef == _GEN_14631 & _GEN_3591 | _GEN_2034; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4590 = 9'h1f0 == _GEN_14631 & _GEN_15783 | _GEN_1523; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4591 = 9'h1f0 == _GEN_14631 & _GEN_3591 | _GEN_2035; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4592 = 9'h1f1 == _GEN_14631 & _GEN_15783 | _GEN_1524; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4593 = 9'h1f1 == _GEN_14631 & _GEN_3591 | _GEN_2036; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4594 = 9'h1f2 == _GEN_14631 & _GEN_15783 | _GEN_1525; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4595 = 9'h1f2 == _GEN_14631 & _GEN_3591 | _GEN_2037; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4596 = 9'h1f3 == _GEN_14631 & _GEN_15783 | _GEN_1526; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4597 = 9'h1f3 == _GEN_14631 & _GEN_3591 | _GEN_2038; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4598 = 9'h1f4 == _GEN_14631 & _GEN_15783 | _GEN_1527; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4599 = 9'h1f4 == _GEN_14631 & _GEN_3591 | _GEN_2039; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4600 = 9'h1f5 == _GEN_14631 & _GEN_15783 | _GEN_1528; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4601 = 9'h1f5 == _GEN_14631 & _GEN_3591 | _GEN_2040; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4602 = 9'h1f6 == _GEN_14631 & _GEN_15783 | _GEN_1529; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4603 = 9'h1f6 == _GEN_14631 & _GEN_3591 | _GEN_2041; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4604 = 9'h1f7 == _GEN_14631 & _GEN_15783 | _GEN_1530; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4605 = 9'h1f7 == _GEN_14631 & _GEN_3591 | _GEN_2042; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4606 = 9'h1f8 == _GEN_14631 & _GEN_15783 | _GEN_1531; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4607 = 9'h1f8 == _GEN_14631 & _GEN_3591 | _GEN_2043; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4608 = 9'h1f9 == _GEN_14631 & _GEN_15783 | _GEN_1532; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4609 = 9'h1f9 == _GEN_14631 & _GEN_3591 | _GEN_2044; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4610 = 9'h1fa == _GEN_14631 & _GEN_15783 | _GEN_1533; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4611 = 9'h1fa == _GEN_14631 & _GEN_3591 | _GEN_2045; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4612 = 9'h1fb == _GEN_14631 & _GEN_15783 | _GEN_1534; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4613 = 9'h1fb == _GEN_14631 & _GEN_3591 | _GEN_2046; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4614 = 9'h1fc == _GEN_14631 & _GEN_15783 | _GEN_1535; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4615 = 9'h1fc == _GEN_14631 & _GEN_3591 | _GEN_2047; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4616 = 9'h1fd == _GEN_14631 & _GEN_15783 | _GEN_1536; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4617 = 9'h1fd == _GEN_14631 & _GEN_3591 | _GEN_2048; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4618 = 9'h1fe == _GEN_14631 & _GEN_15783 | _GEN_1537; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4619 = 9'h1fe == _GEN_14631 & _GEN_3591 | _GEN_2049; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4620 = 9'h1ff == _GEN_14631 & _GEN_15783 | _GEN_1538; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4621 = 9'h1ff == _GEN_14631 & _GEN_3591 | _GEN_2050; // @[ICache.scala 187:{36,36}]
  wire  _GEN_4622 = 6'h0 == vset ? ~tag_compare_valid_1 : lru_0; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4623 = 6'h1 == vset ? ~tag_compare_valid_1 : lru_1; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4624 = 6'h2 == vset ? ~tag_compare_valid_1 : lru_2; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4625 = 6'h3 == vset ? ~tag_compare_valid_1 : lru_3; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4626 = 6'h4 == vset ? ~tag_compare_valid_1 : lru_4; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4627 = 6'h5 == vset ? ~tag_compare_valid_1 : lru_5; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4628 = 6'h6 == vset ? ~tag_compare_valid_1 : lru_6; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4629 = 6'h7 == vset ? ~tag_compare_valid_1 : lru_7; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4630 = 6'h8 == vset ? ~tag_compare_valid_1 : lru_8; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4631 = 6'h9 == vset ? ~tag_compare_valid_1 : lru_9; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4632 = 6'ha == vset ? ~tag_compare_valid_1 : lru_10; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4633 = 6'hb == vset ? ~tag_compare_valid_1 : lru_11; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4634 = 6'hc == vset ? ~tag_compare_valid_1 : lru_12; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4635 = 6'hd == vset ? ~tag_compare_valid_1 : lru_13; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4636 = 6'he == vset ? ~tag_compare_valid_1 : lru_14; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4637 = 6'hf == vset ? ~tag_compare_valid_1 : lru_15; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4638 = 6'h10 == vset ? ~tag_compare_valid_1 : lru_16; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4639 = 6'h11 == vset ? ~tag_compare_valid_1 : lru_17; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4640 = 6'h12 == vset ? ~tag_compare_valid_1 : lru_18; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4641 = 6'h13 == vset ? ~tag_compare_valid_1 : lru_19; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4642 = 6'h14 == vset ? ~tag_compare_valid_1 : lru_20; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4643 = 6'h15 == vset ? ~tag_compare_valid_1 : lru_21; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4644 = 6'h16 == vset ? ~tag_compare_valid_1 : lru_22; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4645 = 6'h17 == vset ? ~tag_compare_valid_1 : lru_23; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4646 = 6'h18 == vset ? ~tag_compare_valid_1 : lru_24; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4647 = 6'h19 == vset ? ~tag_compare_valid_1 : lru_25; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4648 = 6'h1a == vset ? ~tag_compare_valid_1 : lru_26; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4649 = 6'h1b == vset ? ~tag_compare_valid_1 : lru_27; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4650 = 6'h1c == vset ? ~tag_compare_valid_1 : lru_28; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4651 = 6'h1d == vset ? ~tag_compare_valid_1 : lru_29; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4652 = 6'h1e == vset ? ~tag_compare_valid_1 : lru_30; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4653 = 6'h1f == vset ? ~tag_compare_valid_1 : lru_31; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4654 = 6'h20 == vset ? ~tag_compare_valid_1 : lru_32; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4655 = 6'h21 == vset ? ~tag_compare_valid_1 : lru_33; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4656 = 6'h22 == vset ? ~tag_compare_valid_1 : lru_34; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4657 = 6'h23 == vset ? ~tag_compare_valid_1 : lru_35; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4658 = 6'h24 == vset ? ~tag_compare_valid_1 : lru_36; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4659 = 6'h25 == vset ? ~tag_compare_valid_1 : lru_37; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4660 = 6'h26 == vset ? ~tag_compare_valid_1 : lru_38; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4661 = 6'h27 == vset ? ~tag_compare_valid_1 : lru_39; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4662 = 6'h28 == vset ? ~tag_compare_valid_1 : lru_40; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4663 = 6'h29 == vset ? ~tag_compare_valid_1 : lru_41; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4664 = 6'h2a == vset ? ~tag_compare_valid_1 : lru_42; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4665 = 6'h2b == vset ? ~tag_compare_valid_1 : lru_43; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4666 = 6'h2c == vset ? ~tag_compare_valid_1 : lru_44; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4667 = 6'h2d == vset ? ~tag_compare_valid_1 : lru_45; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4668 = 6'h2e == vset ? ~tag_compare_valid_1 : lru_46; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4669 = 6'h2f == vset ? ~tag_compare_valid_1 : lru_47; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4670 = 6'h30 == vset ? ~tag_compare_valid_1 : lru_48; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4671 = 6'h31 == vset ? ~tag_compare_valid_1 : lru_49; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4672 = 6'h32 == vset ? ~tag_compare_valid_1 : lru_50; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4673 = 6'h33 == vset ? ~tag_compare_valid_1 : lru_51; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4674 = 6'h34 == vset ? ~tag_compare_valid_1 : lru_52; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4675 = 6'h35 == vset ? ~tag_compare_valid_1 : lru_53; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4676 = 6'h36 == vset ? ~tag_compare_valid_1 : lru_54; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4677 = 6'h37 == vset ? ~tag_compare_valid_1 : lru_55; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4678 = 6'h38 == vset ? ~tag_compare_valid_1 : lru_56; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4679 = 6'h39 == vset ? ~tag_compare_valid_1 : lru_57; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4680 = 6'h3a == vset ? ~tag_compare_valid_1 : lru_58; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4681 = 6'h3b == vset ? ~tag_compare_valid_1 : lru_59; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4682 = 6'h3c == vset ? ~tag_compare_valid_1 : lru_60; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4683 = 6'h3d == vset ? ~tag_compare_valid_1 : lru_61; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4684 = 6'h3e == vset ? ~tag_compare_valid_1 : lru_62; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4685 = 6'h3f == vset ? ~tag_compare_valid_1 : lru_63; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4686 = 7'h40 == _GEN_14439 ? ~tag_compare_valid_1 : lru_64; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4687 = 7'h41 == _GEN_14439 ? ~tag_compare_valid_1 : lru_65; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4688 = 7'h42 == _GEN_14439 ? ~tag_compare_valid_1 : lru_66; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4689 = 7'h43 == _GEN_14439 ? ~tag_compare_valid_1 : lru_67; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4690 = 7'h44 == _GEN_14439 ? ~tag_compare_valid_1 : lru_68; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4691 = 7'h45 == _GEN_14439 ? ~tag_compare_valid_1 : lru_69; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4692 = 7'h46 == _GEN_14439 ? ~tag_compare_valid_1 : lru_70; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4693 = 7'h47 == _GEN_14439 ? ~tag_compare_valid_1 : lru_71; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4694 = 7'h48 == _GEN_14439 ? ~tag_compare_valid_1 : lru_72; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4695 = 7'h49 == _GEN_14439 ? ~tag_compare_valid_1 : lru_73; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4696 = 7'h4a == _GEN_14439 ? ~tag_compare_valid_1 : lru_74; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4697 = 7'h4b == _GEN_14439 ? ~tag_compare_valid_1 : lru_75; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4698 = 7'h4c == _GEN_14439 ? ~tag_compare_valid_1 : lru_76; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4699 = 7'h4d == _GEN_14439 ? ~tag_compare_valid_1 : lru_77; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4700 = 7'h4e == _GEN_14439 ? ~tag_compare_valid_1 : lru_78; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4701 = 7'h4f == _GEN_14439 ? ~tag_compare_valid_1 : lru_79; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4702 = 7'h50 == _GEN_14439 ? ~tag_compare_valid_1 : lru_80; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4703 = 7'h51 == _GEN_14439 ? ~tag_compare_valid_1 : lru_81; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4704 = 7'h52 == _GEN_14439 ? ~tag_compare_valid_1 : lru_82; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4705 = 7'h53 == _GEN_14439 ? ~tag_compare_valid_1 : lru_83; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4706 = 7'h54 == _GEN_14439 ? ~tag_compare_valid_1 : lru_84; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4707 = 7'h55 == _GEN_14439 ? ~tag_compare_valid_1 : lru_85; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4708 = 7'h56 == _GEN_14439 ? ~tag_compare_valid_1 : lru_86; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4709 = 7'h57 == _GEN_14439 ? ~tag_compare_valid_1 : lru_87; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4710 = 7'h58 == _GEN_14439 ? ~tag_compare_valid_1 : lru_88; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4711 = 7'h59 == _GEN_14439 ? ~tag_compare_valid_1 : lru_89; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4712 = 7'h5a == _GEN_14439 ? ~tag_compare_valid_1 : lru_90; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4713 = 7'h5b == _GEN_14439 ? ~tag_compare_valid_1 : lru_91; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4714 = 7'h5c == _GEN_14439 ? ~tag_compare_valid_1 : lru_92; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4715 = 7'h5d == _GEN_14439 ? ~tag_compare_valid_1 : lru_93; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4716 = 7'h5e == _GEN_14439 ? ~tag_compare_valid_1 : lru_94; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4717 = 7'h5f == _GEN_14439 ? ~tag_compare_valid_1 : lru_95; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4718 = 7'h60 == _GEN_14439 ? ~tag_compare_valid_1 : lru_96; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4719 = 7'h61 == _GEN_14439 ? ~tag_compare_valid_1 : lru_97; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4720 = 7'h62 == _GEN_14439 ? ~tag_compare_valid_1 : lru_98; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4721 = 7'h63 == _GEN_14439 ? ~tag_compare_valid_1 : lru_99; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4722 = 7'h64 == _GEN_14439 ? ~tag_compare_valid_1 : lru_100; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4723 = 7'h65 == _GEN_14439 ? ~tag_compare_valid_1 : lru_101; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4724 = 7'h66 == _GEN_14439 ? ~tag_compare_valid_1 : lru_102; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4725 = 7'h67 == _GEN_14439 ? ~tag_compare_valid_1 : lru_103; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4726 = 7'h68 == _GEN_14439 ? ~tag_compare_valid_1 : lru_104; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4727 = 7'h69 == _GEN_14439 ? ~tag_compare_valid_1 : lru_105; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4728 = 7'h6a == _GEN_14439 ? ~tag_compare_valid_1 : lru_106; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4729 = 7'h6b == _GEN_14439 ? ~tag_compare_valid_1 : lru_107; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4730 = 7'h6c == _GEN_14439 ? ~tag_compare_valid_1 : lru_108; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4731 = 7'h6d == _GEN_14439 ? ~tag_compare_valid_1 : lru_109; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4732 = 7'h6e == _GEN_14439 ? ~tag_compare_valid_1 : lru_110; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4733 = 7'h6f == _GEN_14439 ? ~tag_compare_valid_1 : lru_111; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4734 = 7'h70 == _GEN_14439 ? ~tag_compare_valid_1 : lru_112; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4735 = 7'h71 == _GEN_14439 ? ~tag_compare_valid_1 : lru_113; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4736 = 7'h72 == _GEN_14439 ? ~tag_compare_valid_1 : lru_114; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4737 = 7'h73 == _GEN_14439 ? ~tag_compare_valid_1 : lru_115; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4738 = 7'h74 == _GEN_14439 ? ~tag_compare_valid_1 : lru_116; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4739 = 7'h75 == _GEN_14439 ? ~tag_compare_valid_1 : lru_117; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4740 = 7'h76 == _GEN_14439 ? ~tag_compare_valid_1 : lru_118; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4741 = 7'h77 == _GEN_14439 ? ~tag_compare_valid_1 : lru_119; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4742 = 7'h78 == _GEN_14439 ? ~tag_compare_valid_1 : lru_120; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4743 = 7'h79 == _GEN_14439 ? ~tag_compare_valid_1 : lru_121; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4744 = 7'h7a == _GEN_14439 ? ~tag_compare_valid_1 : lru_122; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4745 = 7'h7b == _GEN_14439 ? ~tag_compare_valid_1 : lru_123; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4746 = 7'h7c == _GEN_14439 ? ~tag_compare_valid_1 : lru_124; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4747 = 7'h7d == _GEN_14439 ? ~tag_compare_valid_1 : lru_125; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4748 = 7'h7e == _GEN_14439 ? ~tag_compare_valid_1 : lru_126; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4749 = 7'h7f == _GEN_14439 ? ~tag_compare_valid_1 : lru_127; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4750 = 8'h80 == _GEN_14503 ? ~tag_compare_valid_1 : lru_128; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4751 = 8'h81 == _GEN_14503 ? ~tag_compare_valid_1 : lru_129; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4752 = 8'h82 == _GEN_14503 ? ~tag_compare_valid_1 : lru_130; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4753 = 8'h83 == _GEN_14503 ? ~tag_compare_valid_1 : lru_131; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4754 = 8'h84 == _GEN_14503 ? ~tag_compare_valid_1 : lru_132; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4755 = 8'h85 == _GEN_14503 ? ~tag_compare_valid_1 : lru_133; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4756 = 8'h86 == _GEN_14503 ? ~tag_compare_valid_1 : lru_134; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4757 = 8'h87 == _GEN_14503 ? ~tag_compare_valid_1 : lru_135; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4758 = 8'h88 == _GEN_14503 ? ~tag_compare_valid_1 : lru_136; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4759 = 8'h89 == _GEN_14503 ? ~tag_compare_valid_1 : lru_137; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4760 = 8'h8a == _GEN_14503 ? ~tag_compare_valid_1 : lru_138; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4761 = 8'h8b == _GEN_14503 ? ~tag_compare_valid_1 : lru_139; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4762 = 8'h8c == _GEN_14503 ? ~tag_compare_valid_1 : lru_140; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4763 = 8'h8d == _GEN_14503 ? ~tag_compare_valid_1 : lru_141; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4764 = 8'h8e == _GEN_14503 ? ~tag_compare_valid_1 : lru_142; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4765 = 8'h8f == _GEN_14503 ? ~tag_compare_valid_1 : lru_143; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4766 = 8'h90 == _GEN_14503 ? ~tag_compare_valid_1 : lru_144; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4767 = 8'h91 == _GEN_14503 ? ~tag_compare_valid_1 : lru_145; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4768 = 8'h92 == _GEN_14503 ? ~tag_compare_valid_1 : lru_146; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4769 = 8'h93 == _GEN_14503 ? ~tag_compare_valid_1 : lru_147; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4770 = 8'h94 == _GEN_14503 ? ~tag_compare_valid_1 : lru_148; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4771 = 8'h95 == _GEN_14503 ? ~tag_compare_valid_1 : lru_149; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4772 = 8'h96 == _GEN_14503 ? ~tag_compare_valid_1 : lru_150; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4773 = 8'h97 == _GEN_14503 ? ~tag_compare_valid_1 : lru_151; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4774 = 8'h98 == _GEN_14503 ? ~tag_compare_valid_1 : lru_152; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4775 = 8'h99 == _GEN_14503 ? ~tag_compare_valid_1 : lru_153; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4776 = 8'h9a == _GEN_14503 ? ~tag_compare_valid_1 : lru_154; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4777 = 8'h9b == _GEN_14503 ? ~tag_compare_valid_1 : lru_155; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4778 = 8'h9c == _GEN_14503 ? ~tag_compare_valid_1 : lru_156; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4779 = 8'h9d == _GEN_14503 ? ~tag_compare_valid_1 : lru_157; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4780 = 8'h9e == _GEN_14503 ? ~tag_compare_valid_1 : lru_158; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4781 = 8'h9f == _GEN_14503 ? ~tag_compare_valid_1 : lru_159; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4782 = 8'ha0 == _GEN_14503 ? ~tag_compare_valid_1 : lru_160; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4783 = 8'ha1 == _GEN_14503 ? ~tag_compare_valid_1 : lru_161; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4784 = 8'ha2 == _GEN_14503 ? ~tag_compare_valid_1 : lru_162; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4785 = 8'ha3 == _GEN_14503 ? ~tag_compare_valid_1 : lru_163; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4786 = 8'ha4 == _GEN_14503 ? ~tag_compare_valid_1 : lru_164; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4787 = 8'ha5 == _GEN_14503 ? ~tag_compare_valid_1 : lru_165; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4788 = 8'ha6 == _GEN_14503 ? ~tag_compare_valid_1 : lru_166; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4789 = 8'ha7 == _GEN_14503 ? ~tag_compare_valid_1 : lru_167; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4790 = 8'ha8 == _GEN_14503 ? ~tag_compare_valid_1 : lru_168; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4791 = 8'ha9 == _GEN_14503 ? ~tag_compare_valid_1 : lru_169; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4792 = 8'haa == _GEN_14503 ? ~tag_compare_valid_1 : lru_170; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4793 = 8'hab == _GEN_14503 ? ~tag_compare_valid_1 : lru_171; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4794 = 8'hac == _GEN_14503 ? ~tag_compare_valid_1 : lru_172; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4795 = 8'had == _GEN_14503 ? ~tag_compare_valid_1 : lru_173; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4796 = 8'hae == _GEN_14503 ? ~tag_compare_valid_1 : lru_174; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4797 = 8'haf == _GEN_14503 ? ~tag_compare_valid_1 : lru_175; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4798 = 8'hb0 == _GEN_14503 ? ~tag_compare_valid_1 : lru_176; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4799 = 8'hb1 == _GEN_14503 ? ~tag_compare_valid_1 : lru_177; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4800 = 8'hb2 == _GEN_14503 ? ~tag_compare_valid_1 : lru_178; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4801 = 8'hb3 == _GEN_14503 ? ~tag_compare_valid_1 : lru_179; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4802 = 8'hb4 == _GEN_14503 ? ~tag_compare_valid_1 : lru_180; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4803 = 8'hb5 == _GEN_14503 ? ~tag_compare_valid_1 : lru_181; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4804 = 8'hb6 == _GEN_14503 ? ~tag_compare_valid_1 : lru_182; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4805 = 8'hb7 == _GEN_14503 ? ~tag_compare_valid_1 : lru_183; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4806 = 8'hb8 == _GEN_14503 ? ~tag_compare_valid_1 : lru_184; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4807 = 8'hb9 == _GEN_14503 ? ~tag_compare_valid_1 : lru_185; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4808 = 8'hba == _GEN_14503 ? ~tag_compare_valid_1 : lru_186; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4809 = 8'hbb == _GEN_14503 ? ~tag_compare_valid_1 : lru_187; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4810 = 8'hbc == _GEN_14503 ? ~tag_compare_valid_1 : lru_188; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4811 = 8'hbd == _GEN_14503 ? ~tag_compare_valid_1 : lru_189; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4812 = 8'hbe == _GEN_14503 ? ~tag_compare_valid_1 : lru_190; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4813 = 8'hbf == _GEN_14503 ? ~tag_compare_valid_1 : lru_191; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4814 = 8'hc0 == _GEN_14503 ? ~tag_compare_valid_1 : lru_192; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4815 = 8'hc1 == _GEN_14503 ? ~tag_compare_valid_1 : lru_193; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4816 = 8'hc2 == _GEN_14503 ? ~tag_compare_valid_1 : lru_194; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4817 = 8'hc3 == _GEN_14503 ? ~tag_compare_valid_1 : lru_195; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4818 = 8'hc4 == _GEN_14503 ? ~tag_compare_valid_1 : lru_196; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4819 = 8'hc5 == _GEN_14503 ? ~tag_compare_valid_1 : lru_197; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4820 = 8'hc6 == _GEN_14503 ? ~tag_compare_valid_1 : lru_198; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4821 = 8'hc7 == _GEN_14503 ? ~tag_compare_valid_1 : lru_199; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4822 = 8'hc8 == _GEN_14503 ? ~tag_compare_valid_1 : lru_200; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4823 = 8'hc9 == _GEN_14503 ? ~tag_compare_valid_1 : lru_201; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4824 = 8'hca == _GEN_14503 ? ~tag_compare_valid_1 : lru_202; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4825 = 8'hcb == _GEN_14503 ? ~tag_compare_valid_1 : lru_203; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4826 = 8'hcc == _GEN_14503 ? ~tag_compare_valid_1 : lru_204; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4827 = 8'hcd == _GEN_14503 ? ~tag_compare_valid_1 : lru_205; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4828 = 8'hce == _GEN_14503 ? ~tag_compare_valid_1 : lru_206; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4829 = 8'hcf == _GEN_14503 ? ~tag_compare_valid_1 : lru_207; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4830 = 8'hd0 == _GEN_14503 ? ~tag_compare_valid_1 : lru_208; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4831 = 8'hd1 == _GEN_14503 ? ~tag_compare_valid_1 : lru_209; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4832 = 8'hd2 == _GEN_14503 ? ~tag_compare_valid_1 : lru_210; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4833 = 8'hd3 == _GEN_14503 ? ~tag_compare_valid_1 : lru_211; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4834 = 8'hd4 == _GEN_14503 ? ~tag_compare_valid_1 : lru_212; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4835 = 8'hd5 == _GEN_14503 ? ~tag_compare_valid_1 : lru_213; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4836 = 8'hd6 == _GEN_14503 ? ~tag_compare_valid_1 : lru_214; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4837 = 8'hd7 == _GEN_14503 ? ~tag_compare_valid_1 : lru_215; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4838 = 8'hd8 == _GEN_14503 ? ~tag_compare_valid_1 : lru_216; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4839 = 8'hd9 == _GEN_14503 ? ~tag_compare_valid_1 : lru_217; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4840 = 8'hda == _GEN_14503 ? ~tag_compare_valid_1 : lru_218; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4841 = 8'hdb == _GEN_14503 ? ~tag_compare_valid_1 : lru_219; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4842 = 8'hdc == _GEN_14503 ? ~tag_compare_valid_1 : lru_220; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4843 = 8'hdd == _GEN_14503 ? ~tag_compare_valid_1 : lru_221; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4844 = 8'hde == _GEN_14503 ? ~tag_compare_valid_1 : lru_222; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4845 = 8'hdf == _GEN_14503 ? ~tag_compare_valid_1 : lru_223; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4846 = 8'he0 == _GEN_14503 ? ~tag_compare_valid_1 : lru_224; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4847 = 8'he1 == _GEN_14503 ? ~tag_compare_valid_1 : lru_225; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4848 = 8'he2 == _GEN_14503 ? ~tag_compare_valid_1 : lru_226; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4849 = 8'he3 == _GEN_14503 ? ~tag_compare_valid_1 : lru_227; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4850 = 8'he4 == _GEN_14503 ? ~tag_compare_valid_1 : lru_228; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4851 = 8'he5 == _GEN_14503 ? ~tag_compare_valid_1 : lru_229; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4852 = 8'he6 == _GEN_14503 ? ~tag_compare_valid_1 : lru_230; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4853 = 8'he7 == _GEN_14503 ? ~tag_compare_valid_1 : lru_231; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4854 = 8'he8 == _GEN_14503 ? ~tag_compare_valid_1 : lru_232; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4855 = 8'he9 == _GEN_14503 ? ~tag_compare_valid_1 : lru_233; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4856 = 8'hea == _GEN_14503 ? ~tag_compare_valid_1 : lru_234; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4857 = 8'heb == _GEN_14503 ? ~tag_compare_valid_1 : lru_235; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4858 = 8'hec == _GEN_14503 ? ~tag_compare_valid_1 : lru_236; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4859 = 8'hed == _GEN_14503 ? ~tag_compare_valid_1 : lru_237; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4860 = 8'hee == _GEN_14503 ? ~tag_compare_valid_1 : lru_238; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4861 = 8'hef == _GEN_14503 ? ~tag_compare_valid_1 : lru_239; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4862 = 8'hf0 == _GEN_14503 ? ~tag_compare_valid_1 : lru_240; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4863 = 8'hf1 == _GEN_14503 ? ~tag_compare_valid_1 : lru_241; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4864 = 8'hf2 == _GEN_14503 ? ~tag_compare_valid_1 : lru_242; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4865 = 8'hf3 == _GEN_14503 ? ~tag_compare_valid_1 : lru_243; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4866 = 8'hf4 == _GEN_14503 ? ~tag_compare_valid_1 : lru_244; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4867 = 8'hf5 == _GEN_14503 ? ~tag_compare_valid_1 : lru_245; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4868 = 8'hf6 == _GEN_14503 ? ~tag_compare_valid_1 : lru_246; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4869 = 8'hf7 == _GEN_14503 ? ~tag_compare_valid_1 : lru_247; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4870 = 8'hf8 == _GEN_14503 ? ~tag_compare_valid_1 : lru_248; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4871 = 8'hf9 == _GEN_14503 ? ~tag_compare_valid_1 : lru_249; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4872 = 8'hfa == _GEN_14503 ? ~tag_compare_valid_1 : lru_250; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4873 = 8'hfb == _GEN_14503 ? ~tag_compare_valid_1 : lru_251; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4874 = 8'hfc == _GEN_14503 ? ~tag_compare_valid_1 : lru_252; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4875 = 8'hfd == _GEN_14503 ? ~tag_compare_valid_1 : lru_253; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4876 = 8'hfe == _GEN_14503 ? ~tag_compare_valid_1 : lru_254; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4877 = 8'hff == _GEN_14503 ? ~tag_compare_valid_1 : lru_255; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4878 = 9'h100 == _GEN_14631 ? ~tag_compare_valid_1 : lru_256; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4879 = 9'h101 == _GEN_14631 ? ~tag_compare_valid_1 : lru_257; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4880 = 9'h102 == _GEN_14631 ? ~tag_compare_valid_1 : lru_258; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4881 = 9'h103 == _GEN_14631 ? ~tag_compare_valid_1 : lru_259; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4882 = 9'h104 == _GEN_14631 ? ~tag_compare_valid_1 : lru_260; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4883 = 9'h105 == _GEN_14631 ? ~tag_compare_valid_1 : lru_261; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4884 = 9'h106 == _GEN_14631 ? ~tag_compare_valid_1 : lru_262; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4885 = 9'h107 == _GEN_14631 ? ~tag_compare_valid_1 : lru_263; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4886 = 9'h108 == _GEN_14631 ? ~tag_compare_valid_1 : lru_264; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4887 = 9'h109 == _GEN_14631 ? ~tag_compare_valid_1 : lru_265; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4888 = 9'h10a == _GEN_14631 ? ~tag_compare_valid_1 : lru_266; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4889 = 9'h10b == _GEN_14631 ? ~tag_compare_valid_1 : lru_267; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4890 = 9'h10c == _GEN_14631 ? ~tag_compare_valid_1 : lru_268; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4891 = 9'h10d == _GEN_14631 ? ~tag_compare_valid_1 : lru_269; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4892 = 9'h10e == _GEN_14631 ? ~tag_compare_valid_1 : lru_270; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4893 = 9'h10f == _GEN_14631 ? ~tag_compare_valid_1 : lru_271; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4894 = 9'h110 == _GEN_14631 ? ~tag_compare_valid_1 : lru_272; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4895 = 9'h111 == _GEN_14631 ? ~tag_compare_valid_1 : lru_273; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4896 = 9'h112 == _GEN_14631 ? ~tag_compare_valid_1 : lru_274; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4897 = 9'h113 == _GEN_14631 ? ~tag_compare_valid_1 : lru_275; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4898 = 9'h114 == _GEN_14631 ? ~tag_compare_valid_1 : lru_276; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4899 = 9'h115 == _GEN_14631 ? ~tag_compare_valid_1 : lru_277; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4900 = 9'h116 == _GEN_14631 ? ~tag_compare_valid_1 : lru_278; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4901 = 9'h117 == _GEN_14631 ? ~tag_compare_valid_1 : lru_279; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4902 = 9'h118 == _GEN_14631 ? ~tag_compare_valid_1 : lru_280; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4903 = 9'h119 == _GEN_14631 ? ~tag_compare_valid_1 : lru_281; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4904 = 9'h11a == _GEN_14631 ? ~tag_compare_valid_1 : lru_282; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4905 = 9'h11b == _GEN_14631 ? ~tag_compare_valid_1 : lru_283; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4906 = 9'h11c == _GEN_14631 ? ~tag_compare_valid_1 : lru_284; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4907 = 9'h11d == _GEN_14631 ? ~tag_compare_valid_1 : lru_285; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4908 = 9'h11e == _GEN_14631 ? ~tag_compare_valid_1 : lru_286; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4909 = 9'h11f == _GEN_14631 ? ~tag_compare_valid_1 : lru_287; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4910 = 9'h120 == _GEN_14631 ? ~tag_compare_valid_1 : lru_288; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4911 = 9'h121 == _GEN_14631 ? ~tag_compare_valid_1 : lru_289; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4912 = 9'h122 == _GEN_14631 ? ~tag_compare_valid_1 : lru_290; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4913 = 9'h123 == _GEN_14631 ? ~tag_compare_valid_1 : lru_291; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4914 = 9'h124 == _GEN_14631 ? ~tag_compare_valid_1 : lru_292; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4915 = 9'h125 == _GEN_14631 ? ~tag_compare_valid_1 : lru_293; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4916 = 9'h126 == _GEN_14631 ? ~tag_compare_valid_1 : lru_294; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4917 = 9'h127 == _GEN_14631 ? ~tag_compare_valid_1 : lru_295; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4918 = 9'h128 == _GEN_14631 ? ~tag_compare_valid_1 : lru_296; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4919 = 9'h129 == _GEN_14631 ? ~tag_compare_valid_1 : lru_297; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4920 = 9'h12a == _GEN_14631 ? ~tag_compare_valid_1 : lru_298; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4921 = 9'h12b == _GEN_14631 ? ~tag_compare_valid_1 : lru_299; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4922 = 9'h12c == _GEN_14631 ? ~tag_compare_valid_1 : lru_300; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4923 = 9'h12d == _GEN_14631 ? ~tag_compare_valid_1 : lru_301; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4924 = 9'h12e == _GEN_14631 ? ~tag_compare_valid_1 : lru_302; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4925 = 9'h12f == _GEN_14631 ? ~tag_compare_valid_1 : lru_303; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4926 = 9'h130 == _GEN_14631 ? ~tag_compare_valid_1 : lru_304; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4927 = 9'h131 == _GEN_14631 ? ~tag_compare_valid_1 : lru_305; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4928 = 9'h132 == _GEN_14631 ? ~tag_compare_valid_1 : lru_306; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4929 = 9'h133 == _GEN_14631 ? ~tag_compare_valid_1 : lru_307; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4930 = 9'h134 == _GEN_14631 ? ~tag_compare_valid_1 : lru_308; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4931 = 9'h135 == _GEN_14631 ? ~tag_compare_valid_1 : lru_309; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4932 = 9'h136 == _GEN_14631 ? ~tag_compare_valid_1 : lru_310; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4933 = 9'h137 == _GEN_14631 ? ~tag_compare_valid_1 : lru_311; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4934 = 9'h138 == _GEN_14631 ? ~tag_compare_valid_1 : lru_312; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4935 = 9'h139 == _GEN_14631 ? ~tag_compare_valid_1 : lru_313; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4936 = 9'h13a == _GEN_14631 ? ~tag_compare_valid_1 : lru_314; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4937 = 9'h13b == _GEN_14631 ? ~tag_compare_valid_1 : lru_315; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4938 = 9'h13c == _GEN_14631 ? ~tag_compare_valid_1 : lru_316; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4939 = 9'h13d == _GEN_14631 ? ~tag_compare_valid_1 : lru_317; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4940 = 9'h13e == _GEN_14631 ? ~tag_compare_valid_1 : lru_318; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4941 = 9'h13f == _GEN_14631 ? ~tag_compare_valid_1 : lru_319; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4942 = 9'h140 == _GEN_14631 ? ~tag_compare_valid_1 : lru_320; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4943 = 9'h141 == _GEN_14631 ? ~tag_compare_valid_1 : lru_321; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4944 = 9'h142 == _GEN_14631 ? ~tag_compare_valid_1 : lru_322; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4945 = 9'h143 == _GEN_14631 ? ~tag_compare_valid_1 : lru_323; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4946 = 9'h144 == _GEN_14631 ? ~tag_compare_valid_1 : lru_324; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4947 = 9'h145 == _GEN_14631 ? ~tag_compare_valid_1 : lru_325; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4948 = 9'h146 == _GEN_14631 ? ~tag_compare_valid_1 : lru_326; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4949 = 9'h147 == _GEN_14631 ? ~tag_compare_valid_1 : lru_327; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4950 = 9'h148 == _GEN_14631 ? ~tag_compare_valid_1 : lru_328; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4951 = 9'h149 == _GEN_14631 ? ~tag_compare_valid_1 : lru_329; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4952 = 9'h14a == _GEN_14631 ? ~tag_compare_valid_1 : lru_330; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4953 = 9'h14b == _GEN_14631 ? ~tag_compare_valid_1 : lru_331; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4954 = 9'h14c == _GEN_14631 ? ~tag_compare_valid_1 : lru_332; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4955 = 9'h14d == _GEN_14631 ? ~tag_compare_valid_1 : lru_333; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4956 = 9'h14e == _GEN_14631 ? ~tag_compare_valid_1 : lru_334; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4957 = 9'h14f == _GEN_14631 ? ~tag_compare_valid_1 : lru_335; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4958 = 9'h150 == _GEN_14631 ? ~tag_compare_valid_1 : lru_336; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4959 = 9'h151 == _GEN_14631 ? ~tag_compare_valid_1 : lru_337; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4960 = 9'h152 == _GEN_14631 ? ~tag_compare_valid_1 : lru_338; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4961 = 9'h153 == _GEN_14631 ? ~tag_compare_valid_1 : lru_339; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4962 = 9'h154 == _GEN_14631 ? ~tag_compare_valid_1 : lru_340; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4963 = 9'h155 == _GEN_14631 ? ~tag_compare_valid_1 : lru_341; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4964 = 9'h156 == _GEN_14631 ? ~tag_compare_valid_1 : lru_342; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4965 = 9'h157 == _GEN_14631 ? ~tag_compare_valid_1 : lru_343; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4966 = 9'h158 == _GEN_14631 ? ~tag_compare_valid_1 : lru_344; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4967 = 9'h159 == _GEN_14631 ? ~tag_compare_valid_1 : lru_345; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4968 = 9'h15a == _GEN_14631 ? ~tag_compare_valid_1 : lru_346; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4969 = 9'h15b == _GEN_14631 ? ~tag_compare_valid_1 : lru_347; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4970 = 9'h15c == _GEN_14631 ? ~tag_compare_valid_1 : lru_348; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4971 = 9'h15d == _GEN_14631 ? ~tag_compare_valid_1 : lru_349; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4972 = 9'h15e == _GEN_14631 ? ~tag_compare_valid_1 : lru_350; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4973 = 9'h15f == _GEN_14631 ? ~tag_compare_valid_1 : lru_351; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4974 = 9'h160 == _GEN_14631 ? ~tag_compare_valid_1 : lru_352; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4975 = 9'h161 == _GEN_14631 ? ~tag_compare_valid_1 : lru_353; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4976 = 9'h162 == _GEN_14631 ? ~tag_compare_valid_1 : lru_354; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4977 = 9'h163 == _GEN_14631 ? ~tag_compare_valid_1 : lru_355; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4978 = 9'h164 == _GEN_14631 ? ~tag_compare_valid_1 : lru_356; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4979 = 9'h165 == _GEN_14631 ? ~tag_compare_valid_1 : lru_357; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4980 = 9'h166 == _GEN_14631 ? ~tag_compare_valid_1 : lru_358; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4981 = 9'h167 == _GEN_14631 ? ~tag_compare_valid_1 : lru_359; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4982 = 9'h168 == _GEN_14631 ? ~tag_compare_valid_1 : lru_360; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4983 = 9'h169 == _GEN_14631 ? ~tag_compare_valid_1 : lru_361; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4984 = 9'h16a == _GEN_14631 ? ~tag_compare_valid_1 : lru_362; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4985 = 9'h16b == _GEN_14631 ? ~tag_compare_valid_1 : lru_363; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4986 = 9'h16c == _GEN_14631 ? ~tag_compare_valid_1 : lru_364; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4987 = 9'h16d == _GEN_14631 ? ~tag_compare_valid_1 : lru_365; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4988 = 9'h16e == _GEN_14631 ? ~tag_compare_valid_1 : lru_366; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4989 = 9'h16f == _GEN_14631 ? ~tag_compare_valid_1 : lru_367; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4990 = 9'h170 == _GEN_14631 ? ~tag_compare_valid_1 : lru_368; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4991 = 9'h171 == _GEN_14631 ? ~tag_compare_valid_1 : lru_369; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4992 = 9'h172 == _GEN_14631 ? ~tag_compare_valid_1 : lru_370; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4993 = 9'h173 == _GEN_14631 ? ~tag_compare_valid_1 : lru_371; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4994 = 9'h174 == _GEN_14631 ? ~tag_compare_valid_1 : lru_372; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4995 = 9'h175 == _GEN_14631 ? ~tag_compare_valid_1 : lru_373; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4996 = 9'h176 == _GEN_14631 ? ~tag_compare_valid_1 : lru_374; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4997 = 9'h177 == _GEN_14631 ? ~tag_compare_valid_1 : lru_375; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4998 = 9'h178 == _GEN_14631 ? ~tag_compare_valid_1 : lru_376; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_4999 = 9'h179 == _GEN_14631 ? ~tag_compare_valid_1 : lru_377; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5000 = 9'h17a == _GEN_14631 ? ~tag_compare_valid_1 : lru_378; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5001 = 9'h17b == _GEN_14631 ? ~tag_compare_valid_1 : lru_379; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5002 = 9'h17c == _GEN_14631 ? ~tag_compare_valid_1 : lru_380; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5003 = 9'h17d == _GEN_14631 ? ~tag_compare_valid_1 : lru_381; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5004 = 9'h17e == _GEN_14631 ? ~tag_compare_valid_1 : lru_382; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5005 = 9'h17f == _GEN_14631 ? ~tag_compare_valid_1 : lru_383; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5006 = 9'h180 == _GEN_14631 ? ~tag_compare_valid_1 : lru_384; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5007 = 9'h181 == _GEN_14631 ? ~tag_compare_valid_1 : lru_385; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5008 = 9'h182 == _GEN_14631 ? ~tag_compare_valid_1 : lru_386; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5009 = 9'h183 == _GEN_14631 ? ~tag_compare_valid_1 : lru_387; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5010 = 9'h184 == _GEN_14631 ? ~tag_compare_valid_1 : lru_388; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5011 = 9'h185 == _GEN_14631 ? ~tag_compare_valid_1 : lru_389; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5012 = 9'h186 == _GEN_14631 ? ~tag_compare_valid_1 : lru_390; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5013 = 9'h187 == _GEN_14631 ? ~tag_compare_valid_1 : lru_391; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5014 = 9'h188 == _GEN_14631 ? ~tag_compare_valid_1 : lru_392; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5015 = 9'h189 == _GEN_14631 ? ~tag_compare_valid_1 : lru_393; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5016 = 9'h18a == _GEN_14631 ? ~tag_compare_valid_1 : lru_394; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5017 = 9'h18b == _GEN_14631 ? ~tag_compare_valid_1 : lru_395; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5018 = 9'h18c == _GEN_14631 ? ~tag_compare_valid_1 : lru_396; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5019 = 9'h18d == _GEN_14631 ? ~tag_compare_valid_1 : lru_397; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5020 = 9'h18e == _GEN_14631 ? ~tag_compare_valid_1 : lru_398; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5021 = 9'h18f == _GEN_14631 ? ~tag_compare_valid_1 : lru_399; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5022 = 9'h190 == _GEN_14631 ? ~tag_compare_valid_1 : lru_400; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5023 = 9'h191 == _GEN_14631 ? ~tag_compare_valid_1 : lru_401; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5024 = 9'h192 == _GEN_14631 ? ~tag_compare_valid_1 : lru_402; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5025 = 9'h193 == _GEN_14631 ? ~tag_compare_valid_1 : lru_403; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5026 = 9'h194 == _GEN_14631 ? ~tag_compare_valid_1 : lru_404; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5027 = 9'h195 == _GEN_14631 ? ~tag_compare_valid_1 : lru_405; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5028 = 9'h196 == _GEN_14631 ? ~tag_compare_valid_1 : lru_406; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5029 = 9'h197 == _GEN_14631 ? ~tag_compare_valid_1 : lru_407; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5030 = 9'h198 == _GEN_14631 ? ~tag_compare_valid_1 : lru_408; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5031 = 9'h199 == _GEN_14631 ? ~tag_compare_valid_1 : lru_409; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5032 = 9'h19a == _GEN_14631 ? ~tag_compare_valid_1 : lru_410; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5033 = 9'h19b == _GEN_14631 ? ~tag_compare_valid_1 : lru_411; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5034 = 9'h19c == _GEN_14631 ? ~tag_compare_valid_1 : lru_412; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5035 = 9'h19d == _GEN_14631 ? ~tag_compare_valid_1 : lru_413; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5036 = 9'h19e == _GEN_14631 ? ~tag_compare_valid_1 : lru_414; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5037 = 9'h19f == _GEN_14631 ? ~tag_compare_valid_1 : lru_415; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5038 = 9'h1a0 == _GEN_14631 ? ~tag_compare_valid_1 : lru_416; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5039 = 9'h1a1 == _GEN_14631 ? ~tag_compare_valid_1 : lru_417; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5040 = 9'h1a2 == _GEN_14631 ? ~tag_compare_valid_1 : lru_418; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5041 = 9'h1a3 == _GEN_14631 ? ~tag_compare_valid_1 : lru_419; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5042 = 9'h1a4 == _GEN_14631 ? ~tag_compare_valid_1 : lru_420; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5043 = 9'h1a5 == _GEN_14631 ? ~tag_compare_valid_1 : lru_421; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5044 = 9'h1a6 == _GEN_14631 ? ~tag_compare_valid_1 : lru_422; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5045 = 9'h1a7 == _GEN_14631 ? ~tag_compare_valid_1 : lru_423; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5046 = 9'h1a8 == _GEN_14631 ? ~tag_compare_valid_1 : lru_424; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5047 = 9'h1a9 == _GEN_14631 ? ~tag_compare_valid_1 : lru_425; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5048 = 9'h1aa == _GEN_14631 ? ~tag_compare_valid_1 : lru_426; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5049 = 9'h1ab == _GEN_14631 ? ~tag_compare_valid_1 : lru_427; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5050 = 9'h1ac == _GEN_14631 ? ~tag_compare_valid_1 : lru_428; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5051 = 9'h1ad == _GEN_14631 ? ~tag_compare_valid_1 : lru_429; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5052 = 9'h1ae == _GEN_14631 ? ~tag_compare_valid_1 : lru_430; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5053 = 9'h1af == _GEN_14631 ? ~tag_compare_valid_1 : lru_431; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5054 = 9'h1b0 == _GEN_14631 ? ~tag_compare_valid_1 : lru_432; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5055 = 9'h1b1 == _GEN_14631 ? ~tag_compare_valid_1 : lru_433; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5056 = 9'h1b2 == _GEN_14631 ? ~tag_compare_valid_1 : lru_434; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5057 = 9'h1b3 == _GEN_14631 ? ~tag_compare_valid_1 : lru_435; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5058 = 9'h1b4 == _GEN_14631 ? ~tag_compare_valid_1 : lru_436; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5059 = 9'h1b5 == _GEN_14631 ? ~tag_compare_valid_1 : lru_437; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5060 = 9'h1b6 == _GEN_14631 ? ~tag_compare_valid_1 : lru_438; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5061 = 9'h1b7 == _GEN_14631 ? ~tag_compare_valid_1 : lru_439; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5062 = 9'h1b8 == _GEN_14631 ? ~tag_compare_valid_1 : lru_440; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5063 = 9'h1b9 == _GEN_14631 ? ~tag_compare_valid_1 : lru_441; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5064 = 9'h1ba == _GEN_14631 ? ~tag_compare_valid_1 : lru_442; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5065 = 9'h1bb == _GEN_14631 ? ~tag_compare_valid_1 : lru_443; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5066 = 9'h1bc == _GEN_14631 ? ~tag_compare_valid_1 : lru_444; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5067 = 9'h1bd == _GEN_14631 ? ~tag_compare_valid_1 : lru_445; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5068 = 9'h1be == _GEN_14631 ? ~tag_compare_valid_1 : lru_446; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5069 = 9'h1bf == _GEN_14631 ? ~tag_compare_valid_1 : lru_447; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5070 = 9'h1c0 == _GEN_14631 ? ~tag_compare_valid_1 : lru_448; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5071 = 9'h1c1 == _GEN_14631 ? ~tag_compare_valid_1 : lru_449; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5072 = 9'h1c2 == _GEN_14631 ? ~tag_compare_valid_1 : lru_450; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5073 = 9'h1c3 == _GEN_14631 ? ~tag_compare_valid_1 : lru_451; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5074 = 9'h1c4 == _GEN_14631 ? ~tag_compare_valid_1 : lru_452; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5075 = 9'h1c5 == _GEN_14631 ? ~tag_compare_valid_1 : lru_453; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5076 = 9'h1c6 == _GEN_14631 ? ~tag_compare_valid_1 : lru_454; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5077 = 9'h1c7 == _GEN_14631 ? ~tag_compare_valid_1 : lru_455; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5078 = 9'h1c8 == _GEN_14631 ? ~tag_compare_valid_1 : lru_456; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5079 = 9'h1c9 == _GEN_14631 ? ~tag_compare_valid_1 : lru_457; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5080 = 9'h1ca == _GEN_14631 ? ~tag_compare_valid_1 : lru_458; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5081 = 9'h1cb == _GEN_14631 ? ~tag_compare_valid_1 : lru_459; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5082 = 9'h1cc == _GEN_14631 ? ~tag_compare_valid_1 : lru_460; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5083 = 9'h1cd == _GEN_14631 ? ~tag_compare_valid_1 : lru_461; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5084 = 9'h1ce == _GEN_14631 ? ~tag_compare_valid_1 : lru_462; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5085 = 9'h1cf == _GEN_14631 ? ~tag_compare_valid_1 : lru_463; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5086 = 9'h1d0 == _GEN_14631 ? ~tag_compare_valid_1 : lru_464; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5087 = 9'h1d1 == _GEN_14631 ? ~tag_compare_valid_1 : lru_465; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5088 = 9'h1d2 == _GEN_14631 ? ~tag_compare_valid_1 : lru_466; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5089 = 9'h1d3 == _GEN_14631 ? ~tag_compare_valid_1 : lru_467; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5090 = 9'h1d4 == _GEN_14631 ? ~tag_compare_valid_1 : lru_468; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5091 = 9'h1d5 == _GEN_14631 ? ~tag_compare_valid_1 : lru_469; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5092 = 9'h1d6 == _GEN_14631 ? ~tag_compare_valid_1 : lru_470; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5093 = 9'h1d7 == _GEN_14631 ? ~tag_compare_valid_1 : lru_471; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5094 = 9'h1d8 == _GEN_14631 ? ~tag_compare_valid_1 : lru_472; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5095 = 9'h1d9 == _GEN_14631 ? ~tag_compare_valid_1 : lru_473; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5096 = 9'h1da == _GEN_14631 ? ~tag_compare_valid_1 : lru_474; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5097 = 9'h1db == _GEN_14631 ? ~tag_compare_valid_1 : lru_475; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5098 = 9'h1dc == _GEN_14631 ? ~tag_compare_valid_1 : lru_476; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5099 = 9'h1dd == _GEN_14631 ? ~tag_compare_valid_1 : lru_477; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5100 = 9'h1de == _GEN_14631 ? ~tag_compare_valid_1 : lru_478; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5101 = 9'h1df == _GEN_14631 ? ~tag_compare_valid_1 : lru_479; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5102 = 9'h1e0 == _GEN_14631 ? ~tag_compare_valid_1 : lru_480; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5103 = 9'h1e1 == _GEN_14631 ? ~tag_compare_valid_1 : lru_481; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5104 = 9'h1e2 == _GEN_14631 ? ~tag_compare_valid_1 : lru_482; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5105 = 9'h1e3 == _GEN_14631 ? ~tag_compare_valid_1 : lru_483; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5106 = 9'h1e4 == _GEN_14631 ? ~tag_compare_valid_1 : lru_484; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5107 = 9'h1e5 == _GEN_14631 ? ~tag_compare_valid_1 : lru_485; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5108 = 9'h1e6 == _GEN_14631 ? ~tag_compare_valid_1 : lru_486; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5109 = 9'h1e7 == _GEN_14631 ? ~tag_compare_valid_1 : lru_487; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5110 = 9'h1e8 == _GEN_14631 ? ~tag_compare_valid_1 : lru_488; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5111 = 9'h1e9 == _GEN_14631 ? ~tag_compare_valid_1 : lru_489; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5112 = 9'h1ea == _GEN_14631 ? ~tag_compare_valid_1 : lru_490; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5113 = 9'h1eb == _GEN_14631 ? ~tag_compare_valid_1 : lru_491; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5114 = 9'h1ec == _GEN_14631 ? ~tag_compare_valid_1 : lru_492; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5115 = 9'h1ed == _GEN_14631 ? ~tag_compare_valid_1 : lru_493; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5116 = 9'h1ee == _GEN_14631 ? ~tag_compare_valid_1 : lru_494; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5117 = 9'h1ef == _GEN_14631 ? ~tag_compare_valid_1 : lru_495; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5118 = 9'h1f0 == _GEN_14631 ? ~tag_compare_valid_1 : lru_496; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5119 = 9'h1f1 == _GEN_14631 ? ~tag_compare_valid_1 : lru_497; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5120 = 9'h1f2 == _GEN_14631 ? ~tag_compare_valid_1 : lru_498; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5121 = 9'h1f3 == _GEN_14631 ? ~tag_compare_valid_1 : lru_499; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5122 = 9'h1f4 == _GEN_14631 ? ~tag_compare_valid_1 : lru_500; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5123 = 9'h1f5 == _GEN_14631 ? ~tag_compare_valid_1 : lru_501; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5124 = 9'h1f6 == _GEN_14631 ? ~tag_compare_valid_1 : lru_502; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5125 = 9'h1f7 == _GEN_14631 ? ~tag_compare_valid_1 : lru_503; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5126 = 9'h1f8 == _GEN_14631 ? ~tag_compare_valid_1 : lru_504; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5127 = 9'h1f9 == _GEN_14631 ? ~tag_compare_valid_1 : lru_505; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5128 = 9'h1fa == _GEN_14631 ? ~tag_compare_valid_1 : lru_506; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5129 = 9'h1fb == _GEN_14631 ? ~tag_compare_valid_1 : lru_507; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5130 = 9'h1fc == _GEN_14631 ? ~tag_compare_valid_1 : lru_508; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5131 = 9'h1fd == _GEN_14631 ? ~tag_compare_valid_1 : lru_509; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5132 = 9'h1fe == _GEN_14631 ? ~tag_compare_valid_1 : lru_510; // @[ICache.scala 190:{21,21} 68:20]
  wire  _GEN_5133 = 9'h1ff == _GEN_14631 ? ~tag_compare_valid_1 : lru_511; // @[ICache.scala 190:{21,21} 68:20]
  wire [2:0] _GEN_5134 = io_cpu_cpu_stall ? 3'h4 : state; // @[ICache.scala 191:34 192:28 39:81]
  wire [31:0] _GEN_5135 = io_cpu_cpu_stall ? data_1_0 : saved_1_inst; // @[ICache.scala 113:22 191:34 193:28]
  wire  _GEN_5136 = io_cpu_cpu_stall ? cache_hit_available : saved_0_valid; // @[ICache.scala 113:22 191:34 194:28]
  wire  _GEN_5137 = io_cpu_cpu_stall ? inst_valid_1 : saved_1_valid; // @[ICache.scala 113:22 191:34 195:28]
  wire  _GEN_5138 = _T ? _GEN_4622 : lru_0; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5139 = _T ? _GEN_4623 : lru_1; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5140 = _T ? _GEN_4624 : lru_2; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5141 = _T ? _GEN_4625 : lru_3; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5142 = _T ? _GEN_4626 : lru_4; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5143 = _T ? _GEN_4627 : lru_5; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5144 = _T ? _GEN_4628 : lru_6; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5145 = _T ? _GEN_4629 : lru_7; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5146 = _T ? _GEN_4630 : lru_8; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5147 = _T ? _GEN_4631 : lru_9; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5148 = _T ? _GEN_4632 : lru_10; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5149 = _T ? _GEN_4633 : lru_11; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5150 = _T ? _GEN_4634 : lru_12; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5151 = _T ? _GEN_4635 : lru_13; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5152 = _T ? _GEN_4636 : lru_14; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5153 = _T ? _GEN_4637 : lru_15; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5154 = _T ? _GEN_4638 : lru_16; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5155 = _T ? _GEN_4639 : lru_17; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5156 = _T ? _GEN_4640 : lru_18; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5157 = _T ? _GEN_4641 : lru_19; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5158 = _T ? _GEN_4642 : lru_20; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5159 = _T ? _GEN_4643 : lru_21; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5160 = _T ? _GEN_4644 : lru_22; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5161 = _T ? _GEN_4645 : lru_23; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5162 = _T ? _GEN_4646 : lru_24; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5163 = _T ? _GEN_4647 : lru_25; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5164 = _T ? _GEN_4648 : lru_26; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5165 = _T ? _GEN_4649 : lru_27; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5166 = _T ? _GEN_4650 : lru_28; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5167 = _T ? _GEN_4651 : lru_29; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5168 = _T ? _GEN_4652 : lru_30; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5169 = _T ? _GEN_4653 : lru_31; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5170 = _T ? _GEN_4654 : lru_32; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5171 = _T ? _GEN_4655 : lru_33; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5172 = _T ? _GEN_4656 : lru_34; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5173 = _T ? _GEN_4657 : lru_35; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5174 = _T ? _GEN_4658 : lru_36; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5175 = _T ? _GEN_4659 : lru_37; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5176 = _T ? _GEN_4660 : lru_38; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5177 = _T ? _GEN_4661 : lru_39; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5178 = _T ? _GEN_4662 : lru_40; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5179 = _T ? _GEN_4663 : lru_41; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5180 = _T ? _GEN_4664 : lru_42; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5181 = _T ? _GEN_4665 : lru_43; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5182 = _T ? _GEN_4666 : lru_44; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5183 = _T ? _GEN_4667 : lru_45; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5184 = _T ? _GEN_4668 : lru_46; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5185 = _T ? _GEN_4669 : lru_47; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5186 = _T ? _GEN_4670 : lru_48; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5187 = _T ? _GEN_4671 : lru_49; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5188 = _T ? _GEN_4672 : lru_50; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5189 = _T ? _GEN_4673 : lru_51; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5190 = _T ? _GEN_4674 : lru_52; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5191 = _T ? _GEN_4675 : lru_53; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5192 = _T ? _GEN_4676 : lru_54; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5193 = _T ? _GEN_4677 : lru_55; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5194 = _T ? _GEN_4678 : lru_56; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5195 = _T ? _GEN_4679 : lru_57; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5196 = _T ? _GEN_4680 : lru_58; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5197 = _T ? _GEN_4681 : lru_59; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5198 = _T ? _GEN_4682 : lru_60; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5199 = _T ? _GEN_4683 : lru_61; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5200 = _T ? _GEN_4684 : lru_62; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5201 = _T ? _GEN_4685 : lru_63; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5202 = _T ? _GEN_4686 : lru_64; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5203 = _T ? _GEN_4687 : lru_65; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5204 = _T ? _GEN_4688 : lru_66; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5205 = _T ? _GEN_4689 : lru_67; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5206 = _T ? _GEN_4690 : lru_68; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5207 = _T ? _GEN_4691 : lru_69; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5208 = _T ? _GEN_4692 : lru_70; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5209 = _T ? _GEN_4693 : lru_71; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5210 = _T ? _GEN_4694 : lru_72; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5211 = _T ? _GEN_4695 : lru_73; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5212 = _T ? _GEN_4696 : lru_74; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5213 = _T ? _GEN_4697 : lru_75; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5214 = _T ? _GEN_4698 : lru_76; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5215 = _T ? _GEN_4699 : lru_77; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5216 = _T ? _GEN_4700 : lru_78; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5217 = _T ? _GEN_4701 : lru_79; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5218 = _T ? _GEN_4702 : lru_80; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5219 = _T ? _GEN_4703 : lru_81; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5220 = _T ? _GEN_4704 : lru_82; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5221 = _T ? _GEN_4705 : lru_83; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5222 = _T ? _GEN_4706 : lru_84; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5223 = _T ? _GEN_4707 : lru_85; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5224 = _T ? _GEN_4708 : lru_86; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5225 = _T ? _GEN_4709 : lru_87; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5226 = _T ? _GEN_4710 : lru_88; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5227 = _T ? _GEN_4711 : lru_89; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5228 = _T ? _GEN_4712 : lru_90; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5229 = _T ? _GEN_4713 : lru_91; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5230 = _T ? _GEN_4714 : lru_92; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5231 = _T ? _GEN_4715 : lru_93; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5232 = _T ? _GEN_4716 : lru_94; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5233 = _T ? _GEN_4717 : lru_95; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5234 = _T ? _GEN_4718 : lru_96; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5235 = _T ? _GEN_4719 : lru_97; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5236 = _T ? _GEN_4720 : lru_98; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5237 = _T ? _GEN_4721 : lru_99; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5238 = _T ? _GEN_4722 : lru_100; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5239 = _T ? _GEN_4723 : lru_101; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5240 = _T ? _GEN_4724 : lru_102; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5241 = _T ? _GEN_4725 : lru_103; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5242 = _T ? _GEN_4726 : lru_104; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5243 = _T ? _GEN_4727 : lru_105; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5244 = _T ? _GEN_4728 : lru_106; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5245 = _T ? _GEN_4729 : lru_107; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5246 = _T ? _GEN_4730 : lru_108; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5247 = _T ? _GEN_4731 : lru_109; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5248 = _T ? _GEN_4732 : lru_110; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5249 = _T ? _GEN_4733 : lru_111; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5250 = _T ? _GEN_4734 : lru_112; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5251 = _T ? _GEN_4735 : lru_113; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5252 = _T ? _GEN_4736 : lru_114; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5253 = _T ? _GEN_4737 : lru_115; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5254 = _T ? _GEN_4738 : lru_116; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5255 = _T ? _GEN_4739 : lru_117; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5256 = _T ? _GEN_4740 : lru_118; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5257 = _T ? _GEN_4741 : lru_119; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5258 = _T ? _GEN_4742 : lru_120; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5259 = _T ? _GEN_4743 : lru_121; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5260 = _T ? _GEN_4744 : lru_122; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5261 = _T ? _GEN_4745 : lru_123; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5262 = _T ? _GEN_4746 : lru_124; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5263 = _T ? _GEN_4747 : lru_125; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5264 = _T ? _GEN_4748 : lru_126; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5265 = _T ? _GEN_4749 : lru_127; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5266 = _T ? _GEN_4750 : lru_128; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5267 = _T ? _GEN_4751 : lru_129; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5268 = _T ? _GEN_4752 : lru_130; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5269 = _T ? _GEN_4753 : lru_131; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5270 = _T ? _GEN_4754 : lru_132; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5271 = _T ? _GEN_4755 : lru_133; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5272 = _T ? _GEN_4756 : lru_134; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5273 = _T ? _GEN_4757 : lru_135; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5274 = _T ? _GEN_4758 : lru_136; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5275 = _T ? _GEN_4759 : lru_137; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5276 = _T ? _GEN_4760 : lru_138; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5277 = _T ? _GEN_4761 : lru_139; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5278 = _T ? _GEN_4762 : lru_140; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5279 = _T ? _GEN_4763 : lru_141; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5280 = _T ? _GEN_4764 : lru_142; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5281 = _T ? _GEN_4765 : lru_143; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5282 = _T ? _GEN_4766 : lru_144; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5283 = _T ? _GEN_4767 : lru_145; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5284 = _T ? _GEN_4768 : lru_146; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5285 = _T ? _GEN_4769 : lru_147; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5286 = _T ? _GEN_4770 : lru_148; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5287 = _T ? _GEN_4771 : lru_149; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5288 = _T ? _GEN_4772 : lru_150; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5289 = _T ? _GEN_4773 : lru_151; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5290 = _T ? _GEN_4774 : lru_152; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5291 = _T ? _GEN_4775 : lru_153; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5292 = _T ? _GEN_4776 : lru_154; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5293 = _T ? _GEN_4777 : lru_155; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5294 = _T ? _GEN_4778 : lru_156; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5295 = _T ? _GEN_4779 : lru_157; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5296 = _T ? _GEN_4780 : lru_158; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5297 = _T ? _GEN_4781 : lru_159; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5298 = _T ? _GEN_4782 : lru_160; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5299 = _T ? _GEN_4783 : lru_161; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5300 = _T ? _GEN_4784 : lru_162; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5301 = _T ? _GEN_4785 : lru_163; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5302 = _T ? _GEN_4786 : lru_164; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5303 = _T ? _GEN_4787 : lru_165; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5304 = _T ? _GEN_4788 : lru_166; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5305 = _T ? _GEN_4789 : lru_167; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5306 = _T ? _GEN_4790 : lru_168; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5307 = _T ? _GEN_4791 : lru_169; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5308 = _T ? _GEN_4792 : lru_170; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5309 = _T ? _GEN_4793 : lru_171; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5310 = _T ? _GEN_4794 : lru_172; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5311 = _T ? _GEN_4795 : lru_173; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5312 = _T ? _GEN_4796 : lru_174; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5313 = _T ? _GEN_4797 : lru_175; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5314 = _T ? _GEN_4798 : lru_176; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5315 = _T ? _GEN_4799 : lru_177; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5316 = _T ? _GEN_4800 : lru_178; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5317 = _T ? _GEN_4801 : lru_179; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5318 = _T ? _GEN_4802 : lru_180; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5319 = _T ? _GEN_4803 : lru_181; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5320 = _T ? _GEN_4804 : lru_182; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5321 = _T ? _GEN_4805 : lru_183; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5322 = _T ? _GEN_4806 : lru_184; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5323 = _T ? _GEN_4807 : lru_185; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5324 = _T ? _GEN_4808 : lru_186; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5325 = _T ? _GEN_4809 : lru_187; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5326 = _T ? _GEN_4810 : lru_188; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5327 = _T ? _GEN_4811 : lru_189; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5328 = _T ? _GEN_4812 : lru_190; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5329 = _T ? _GEN_4813 : lru_191; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5330 = _T ? _GEN_4814 : lru_192; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5331 = _T ? _GEN_4815 : lru_193; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5332 = _T ? _GEN_4816 : lru_194; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5333 = _T ? _GEN_4817 : lru_195; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5334 = _T ? _GEN_4818 : lru_196; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5335 = _T ? _GEN_4819 : lru_197; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5336 = _T ? _GEN_4820 : lru_198; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5337 = _T ? _GEN_4821 : lru_199; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5338 = _T ? _GEN_4822 : lru_200; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5339 = _T ? _GEN_4823 : lru_201; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5340 = _T ? _GEN_4824 : lru_202; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5341 = _T ? _GEN_4825 : lru_203; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5342 = _T ? _GEN_4826 : lru_204; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5343 = _T ? _GEN_4827 : lru_205; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5344 = _T ? _GEN_4828 : lru_206; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5345 = _T ? _GEN_4829 : lru_207; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5346 = _T ? _GEN_4830 : lru_208; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5347 = _T ? _GEN_4831 : lru_209; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5348 = _T ? _GEN_4832 : lru_210; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5349 = _T ? _GEN_4833 : lru_211; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5350 = _T ? _GEN_4834 : lru_212; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5351 = _T ? _GEN_4835 : lru_213; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5352 = _T ? _GEN_4836 : lru_214; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5353 = _T ? _GEN_4837 : lru_215; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5354 = _T ? _GEN_4838 : lru_216; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5355 = _T ? _GEN_4839 : lru_217; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5356 = _T ? _GEN_4840 : lru_218; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5357 = _T ? _GEN_4841 : lru_219; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5358 = _T ? _GEN_4842 : lru_220; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5359 = _T ? _GEN_4843 : lru_221; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5360 = _T ? _GEN_4844 : lru_222; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5361 = _T ? _GEN_4845 : lru_223; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5362 = _T ? _GEN_4846 : lru_224; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5363 = _T ? _GEN_4847 : lru_225; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5364 = _T ? _GEN_4848 : lru_226; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5365 = _T ? _GEN_4849 : lru_227; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5366 = _T ? _GEN_4850 : lru_228; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5367 = _T ? _GEN_4851 : lru_229; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5368 = _T ? _GEN_4852 : lru_230; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5369 = _T ? _GEN_4853 : lru_231; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5370 = _T ? _GEN_4854 : lru_232; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5371 = _T ? _GEN_4855 : lru_233; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5372 = _T ? _GEN_4856 : lru_234; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5373 = _T ? _GEN_4857 : lru_235; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5374 = _T ? _GEN_4858 : lru_236; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5375 = _T ? _GEN_4859 : lru_237; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5376 = _T ? _GEN_4860 : lru_238; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5377 = _T ? _GEN_4861 : lru_239; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5378 = _T ? _GEN_4862 : lru_240; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5379 = _T ? _GEN_4863 : lru_241; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5380 = _T ? _GEN_4864 : lru_242; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5381 = _T ? _GEN_4865 : lru_243; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5382 = _T ? _GEN_4866 : lru_244; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5383 = _T ? _GEN_4867 : lru_245; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5384 = _T ? _GEN_4868 : lru_246; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5385 = _T ? _GEN_4869 : lru_247; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5386 = _T ? _GEN_4870 : lru_248; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5387 = _T ? _GEN_4871 : lru_249; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5388 = _T ? _GEN_4872 : lru_250; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5389 = _T ? _GEN_4873 : lru_251; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5390 = _T ? _GEN_4874 : lru_252; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5391 = _T ? _GEN_4875 : lru_253; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5392 = _T ? _GEN_4876 : lru_254; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5393 = _T ? _GEN_4877 : lru_255; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5394 = _T ? _GEN_4878 : lru_256; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5395 = _T ? _GEN_4879 : lru_257; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5396 = _T ? _GEN_4880 : lru_258; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5397 = _T ? _GEN_4881 : lru_259; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5398 = _T ? _GEN_4882 : lru_260; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5399 = _T ? _GEN_4883 : lru_261; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5400 = _T ? _GEN_4884 : lru_262; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5401 = _T ? _GEN_4885 : lru_263; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5402 = _T ? _GEN_4886 : lru_264; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5403 = _T ? _GEN_4887 : lru_265; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5404 = _T ? _GEN_4888 : lru_266; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5405 = _T ? _GEN_4889 : lru_267; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5406 = _T ? _GEN_4890 : lru_268; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5407 = _T ? _GEN_4891 : lru_269; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5408 = _T ? _GEN_4892 : lru_270; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5409 = _T ? _GEN_4893 : lru_271; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5410 = _T ? _GEN_4894 : lru_272; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5411 = _T ? _GEN_4895 : lru_273; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5412 = _T ? _GEN_4896 : lru_274; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5413 = _T ? _GEN_4897 : lru_275; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5414 = _T ? _GEN_4898 : lru_276; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5415 = _T ? _GEN_4899 : lru_277; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5416 = _T ? _GEN_4900 : lru_278; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5417 = _T ? _GEN_4901 : lru_279; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5418 = _T ? _GEN_4902 : lru_280; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5419 = _T ? _GEN_4903 : lru_281; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5420 = _T ? _GEN_4904 : lru_282; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5421 = _T ? _GEN_4905 : lru_283; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5422 = _T ? _GEN_4906 : lru_284; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5423 = _T ? _GEN_4907 : lru_285; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5424 = _T ? _GEN_4908 : lru_286; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5425 = _T ? _GEN_4909 : lru_287; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5426 = _T ? _GEN_4910 : lru_288; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5427 = _T ? _GEN_4911 : lru_289; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5428 = _T ? _GEN_4912 : lru_290; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5429 = _T ? _GEN_4913 : lru_291; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5430 = _T ? _GEN_4914 : lru_292; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5431 = _T ? _GEN_4915 : lru_293; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5432 = _T ? _GEN_4916 : lru_294; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5433 = _T ? _GEN_4917 : lru_295; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5434 = _T ? _GEN_4918 : lru_296; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5435 = _T ? _GEN_4919 : lru_297; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5436 = _T ? _GEN_4920 : lru_298; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5437 = _T ? _GEN_4921 : lru_299; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5438 = _T ? _GEN_4922 : lru_300; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5439 = _T ? _GEN_4923 : lru_301; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5440 = _T ? _GEN_4924 : lru_302; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5441 = _T ? _GEN_4925 : lru_303; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5442 = _T ? _GEN_4926 : lru_304; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5443 = _T ? _GEN_4927 : lru_305; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5444 = _T ? _GEN_4928 : lru_306; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5445 = _T ? _GEN_4929 : lru_307; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5446 = _T ? _GEN_4930 : lru_308; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5447 = _T ? _GEN_4931 : lru_309; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5448 = _T ? _GEN_4932 : lru_310; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5449 = _T ? _GEN_4933 : lru_311; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5450 = _T ? _GEN_4934 : lru_312; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5451 = _T ? _GEN_4935 : lru_313; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5452 = _T ? _GEN_4936 : lru_314; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5453 = _T ? _GEN_4937 : lru_315; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5454 = _T ? _GEN_4938 : lru_316; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5455 = _T ? _GEN_4939 : lru_317; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5456 = _T ? _GEN_4940 : lru_318; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5457 = _T ? _GEN_4941 : lru_319; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5458 = _T ? _GEN_4942 : lru_320; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5459 = _T ? _GEN_4943 : lru_321; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5460 = _T ? _GEN_4944 : lru_322; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5461 = _T ? _GEN_4945 : lru_323; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5462 = _T ? _GEN_4946 : lru_324; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5463 = _T ? _GEN_4947 : lru_325; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5464 = _T ? _GEN_4948 : lru_326; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5465 = _T ? _GEN_4949 : lru_327; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5466 = _T ? _GEN_4950 : lru_328; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5467 = _T ? _GEN_4951 : lru_329; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5468 = _T ? _GEN_4952 : lru_330; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5469 = _T ? _GEN_4953 : lru_331; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5470 = _T ? _GEN_4954 : lru_332; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5471 = _T ? _GEN_4955 : lru_333; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5472 = _T ? _GEN_4956 : lru_334; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5473 = _T ? _GEN_4957 : lru_335; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5474 = _T ? _GEN_4958 : lru_336; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5475 = _T ? _GEN_4959 : lru_337; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5476 = _T ? _GEN_4960 : lru_338; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5477 = _T ? _GEN_4961 : lru_339; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5478 = _T ? _GEN_4962 : lru_340; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5479 = _T ? _GEN_4963 : lru_341; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5480 = _T ? _GEN_4964 : lru_342; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5481 = _T ? _GEN_4965 : lru_343; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5482 = _T ? _GEN_4966 : lru_344; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5483 = _T ? _GEN_4967 : lru_345; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5484 = _T ? _GEN_4968 : lru_346; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5485 = _T ? _GEN_4969 : lru_347; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5486 = _T ? _GEN_4970 : lru_348; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5487 = _T ? _GEN_4971 : lru_349; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5488 = _T ? _GEN_4972 : lru_350; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5489 = _T ? _GEN_4973 : lru_351; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5490 = _T ? _GEN_4974 : lru_352; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5491 = _T ? _GEN_4975 : lru_353; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5492 = _T ? _GEN_4976 : lru_354; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5493 = _T ? _GEN_4977 : lru_355; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5494 = _T ? _GEN_4978 : lru_356; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5495 = _T ? _GEN_4979 : lru_357; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5496 = _T ? _GEN_4980 : lru_358; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5497 = _T ? _GEN_4981 : lru_359; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5498 = _T ? _GEN_4982 : lru_360; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5499 = _T ? _GEN_4983 : lru_361; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5500 = _T ? _GEN_4984 : lru_362; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5501 = _T ? _GEN_4985 : lru_363; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5502 = _T ? _GEN_4986 : lru_364; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5503 = _T ? _GEN_4987 : lru_365; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5504 = _T ? _GEN_4988 : lru_366; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5505 = _T ? _GEN_4989 : lru_367; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5506 = _T ? _GEN_4990 : lru_368; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5507 = _T ? _GEN_4991 : lru_369; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5508 = _T ? _GEN_4992 : lru_370; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5509 = _T ? _GEN_4993 : lru_371; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5510 = _T ? _GEN_4994 : lru_372; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5511 = _T ? _GEN_4995 : lru_373; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5512 = _T ? _GEN_4996 : lru_374; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5513 = _T ? _GEN_4997 : lru_375; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5514 = _T ? _GEN_4998 : lru_376; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5515 = _T ? _GEN_4999 : lru_377; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5516 = _T ? _GEN_5000 : lru_378; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5517 = _T ? _GEN_5001 : lru_379; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5518 = _T ? _GEN_5002 : lru_380; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5519 = _T ? _GEN_5003 : lru_381; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5520 = _T ? _GEN_5004 : lru_382; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5521 = _T ? _GEN_5005 : lru_383; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5522 = _T ? _GEN_5006 : lru_384; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5523 = _T ? _GEN_5007 : lru_385; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5524 = _T ? _GEN_5008 : lru_386; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5525 = _T ? _GEN_5009 : lru_387; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5526 = _T ? _GEN_5010 : lru_388; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5527 = _T ? _GEN_5011 : lru_389; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5528 = _T ? _GEN_5012 : lru_390; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5529 = _T ? _GEN_5013 : lru_391; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5530 = _T ? _GEN_5014 : lru_392; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5531 = _T ? _GEN_5015 : lru_393; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5532 = _T ? _GEN_5016 : lru_394; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5533 = _T ? _GEN_5017 : lru_395; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5534 = _T ? _GEN_5018 : lru_396; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5535 = _T ? _GEN_5019 : lru_397; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5536 = _T ? _GEN_5020 : lru_398; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5537 = _T ? _GEN_5021 : lru_399; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5538 = _T ? _GEN_5022 : lru_400; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5539 = _T ? _GEN_5023 : lru_401; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5540 = _T ? _GEN_5024 : lru_402; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5541 = _T ? _GEN_5025 : lru_403; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5542 = _T ? _GEN_5026 : lru_404; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5543 = _T ? _GEN_5027 : lru_405; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5544 = _T ? _GEN_5028 : lru_406; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5545 = _T ? _GEN_5029 : lru_407; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5546 = _T ? _GEN_5030 : lru_408; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5547 = _T ? _GEN_5031 : lru_409; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5548 = _T ? _GEN_5032 : lru_410; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5549 = _T ? _GEN_5033 : lru_411; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5550 = _T ? _GEN_5034 : lru_412; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5551 = _T ? _GEN_5035 : lru_413; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5552 = _T ? _GEN_5036 : lru_414; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5553 = _T ? _GEN_5037 : lru_415; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5554 = _T ? _GEN_5038 : lru_416; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5555 = _T ? _GEN_5039 : lru_417; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5556 = _T ? _GEN_5040 : lru_418; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5557 = _T ? _GEN_5041 : lru_419; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5558 = _T ? _GEN_5042 : lru_420; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5559 = _T ? _GEN_5043 : lru_421; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5560 = _T ? _GEN_5044 : lru_422; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5561 = _T ? _GEN_5045 : lru_423; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5562 = _T ? _GEN_5046 : lru_424; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5563 = _T ? _GEN_5047 : lru_425; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5564 = _T ? _GEN_5048 : lru_426; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5565 = _T ? _GEN_5049 : lru_427; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5566 = _T ? _GEN_5050 : lru_428; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5567 = _T ? _GEN_5051 : lru_429; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5568 = _T ? _GEN_5052 : lru_430; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5569 = _T ? _GEN_5053 : lru_431; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5570 = _T ? _GEN_5054 : lru_432; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5571 = _T ? _GEN_5055 : lru_433; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5572 = _T ? _GEN_5056 : lru_434; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5573 = _T ? _GEN_5057 : lru_435; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5574 = _T ? _GEN_5058 : lru_436; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5575 = _T ? _GEN_5059 : lru_437; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5576 = _T ? _GEN_5060 : lru_438; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5577 = _T ? _GEN_5061 : lru_439; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5578 = _T ? _GEN_5062 : lru_440; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5579 = _T ? _GEN_5063 : lru_441; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5580 = _T ? _GEN_5064 : lru_442; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5581 = _T ? _GEN_5065 : lru_443; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5582 = _T ? _GEN_5066 : lru_444; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5583 = _T ? _GEN_5067 : lru_445; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5584 = _T ? _GEN_5068 : lru_446; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5585 = _T ? _GEN_5069 : lru_447; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5586 = _T ? _GEN_5070 : lru_448; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5587 = _T ? _GEN_5071 : lru_449; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5588 = _T ? _GEN_5072 : lru_450; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5589 = _T ? _GEN_5073 : lru_451; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5590 = _T ? _GEN_5074 : lru_452; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5591 = _T ? _GEN_5075 : lru_453; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5592 = _T ? _GEN_5076 : lru_454; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5593 = _T ? _GEN_5077 : lru_455; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5594 = _T ? _GEN_5078 : lru_456; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5595 = _T ? _GEN_5079 : lru_457; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5596 = _T ? _GEN_5080 : lru_458; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5597 = _T ? _GEN_5081 : lru_459; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5598 = _T ? _GEN_5082 : lru_460; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5599 = _T ? _GEN_5083 : lru_461; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5600 = _T ? _GEN_5084 : lru_462; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5601 = _T ? _GEN_5085 : lru_463; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5602 = _T ? _GEN_5086 : lru_464; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5603 = _T ? _GEN_5087 : lru_465; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5604 = _T ? _GEN_5088 : lru_466; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5605 = _T ? _GEN_5089 : lru_467; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5606 = _T ? _GEN_5090 : lru_468; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5607 = _T ? _GEN_5091 : lru_469; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5608 = _T ? _GEN_5092 : lru_470; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5609 = _T ? _GEN_5093 : lru_471; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5610 = _T ? _GEN_5094 : lru_472; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5611 = _T ? _GEN_5095 : lru_473; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5612 = _T ? _GEN_5096 : lru_474; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5613 = _T ? _GEN_5097 : lru_475; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5614 = _T ? _GEN_5098 : lru_476; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5615 = _T ? _GEN_5099 : lru_477; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5616 = _T ? _GEN_5100 : lru_478; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5617 = _T ? _GEN_5101 : lru_479; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5618 = _T ? _GEN_5102 : lru_480; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5619 = _T ? _GEN_5103 : lru_481; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5620 = _T ? _GEN_5104 : lru_482; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5621 = _T ? _GEN_5105 : lru_483; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5622 = _T ? _GEN_5106 : lru_484; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5623 = _T ? _GEN_5107 : lru_485; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5624 = _T ? _GEN_5108 : lru_486; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5625 = _T ? _GEN_5109 : lru_487; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5626 = _T ? _GEN_5110 : lru_488; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5627 = _T ? _GEN_5111 : lru_489; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5628 = _T ? _GEN_5112 : lru_490; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5629 = _T ? _GEN_5113 : lru_491; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5630 = _T ? _GEN_5114 : lru_492; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5631 = _T ? _GEN_5115 : lru_493; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5632 = _T ? _GEN_5116 : lru_494; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5633 = _T ? _GEN_5117 : lru_495; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5634 = _T ? _GEN_5118 : lru_496; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5635 = _T ? _GEN_5119 : lru_497; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5636 = _T ? _GEN_5120 : lru_498; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5637 = _T ? _GEN_5121 : lru_499; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5638 = _T ? _GEN_5122 : lru_500; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5639 = _T ? _GEN_5123 : lru_501; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5640 = _T ? _GEN_5124 : lru_502; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5641 = _T ? _GEN_5125 : lru_503; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5642 = _T ? _GEN_5126 : lru_504; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5643 = _T ? _GEN_5127 : lru_505; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5644 = _T ? _GEN_5128 : lru_506; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5645 = _T ? _GEN_5129 : lru_507; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5646 = _T ? _GEN_5130 : lru_508; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5647 = _T ? _GEN_5131 : lru_509; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5648 = _T ? _GEN_5132 : lru_510; // @[ICache.scala 189:42 68:20]
  wire  _GEN_5649 = _T ? _GEN_5133 : lru_511; // @[ICache.scala 189:42 68:20]
  wire [2:0] _GEN_5650 = _T ? _GEN_5134 : state; // @[ICache.scala 189:42 39:81]
  wire [31:0] _GEN_5651 = _T ? _GEN_5135 : saved_1_inst; // @[ICache.scala 113:22 189:42]
  wire  _GEN_5652 = _T ? _GEN_5136 : saved_0_valid; // @[ICache.scala 113:22 189:42]
  wire  _GEN_5653 = _T ? _GEN_5137 : saved_1_valid; // @[ICache.scala 113:22 189:42]
  wire [2:0] _GEN_5654 = ~cache_hit ? 3'h3 : _GEN_5650; // @[ICache.scala 175:32 176:19]
  wire [31:0] _GEN_5655 = ~cache_hit ? _ar_addr_T_1 : ar_addr; // @[ICache.scala 175:32 177:19 149:24]
  wire [7:0] _GEN_5656 = ~cache_hit ? 8'hf : ar_len; // @[ICache.scala 175:32 178:19 149:24]
  wire [2:0] _GEN_5657 = ~cache_hit ? 3'h2 : ar_size; // @[ICache.scala 175:32 179:19 149:24]
  wire  _GEN_5658 = ~cache_hit | arvalid; // @[ICache.scala 175:32 180:19 150:24]
  wire [5:0] _GEN_5659 = ~cache_hit ? vset : rset; // @[ICache.scala 175:32 182:36 95:21]
  wire [3:0] _GEN_5660 = ~cache_hit ? _GEN_3592 : data_wstrb_0_0; // @[ICache.scala 175:32 61:27]
  wire [3:0] _GEN_5661 = ~cache_hit ? _GEN_3593 : data_wstrb_1_0; // @[ICache.scala 175:32 61:27]
  wire [3:0] _GEN_5662 = ~cache_hit ? _GEN_3594 : data_wstrb_0_1; // @[ICache.scala 175:32 61:27]
  wire [3:0] _GEN_5663 = ~cache_hit ? _GEN_3595 : data_wstrb_1_1; // @[ICache.scala 175:32 61:27]
  wire  _GEN_5664 = ~cache_hit ? _GEN_3596 : tag_wstrb_0; // @[ICache.scala 175:32 64:26]
  wire  _GEN_5665 = ~cache_hit ? _GEN_3597 : tag_wstrb_1; // @[ICache.scala 175:32 64:26]
  wire [19:0] _GEN_5666 = ~cache_hit ? inst_tag : tag_wdata; // @[ICache.scala 175:32 186:36 65:26]
  wire  _GEN_5667 = ~cache_hit ? _GEN_3598 : _GEN_1027; // @[ICache.scala 175:32]
  wire  _GEN_5668 = ~cache_hit ? _GEN_3599 : _GEN_1539; // @[ICache.scala 175:32]
  wire  _GEN_5669 = ~cache_hit ? _GEN_3600 : _GEN_1028; // @[ICache.scala 175:32]
  wire  _GEN_5670 = ~cache_hit ? _GEN_3601 : _GEN_1540; // @[ICache.scala 175:32]
  wire  _GEN_5671 = ~cache_hit ? _GEN_3602 : _GEN_1029; // @[ICache.scala 175:32]
  wire  _GEN_5672 = ~cache_hit ? _GEN_3603 : _GEN_1541; // @[ICache.scala 175:32]
  wire  _GEN_5673 = ~cache_hit ? _GEN_3604 : _GEN_1030; // @[ICache.scala 175:32]
  wire  _GEN_5674 = ~cache_hit ? _GEN_3605 : _GEN_1542; // @[ICache.scala 175:32]
  wire  _GEN_5675 = ~cache_hit ? _GEN_3606 : _GEN_1031; // @[ICache.scala 175:32]
  wire  _GEN_5676 = ~cache_hit ? _GEN_3607 : _GEN_1543; // @[ICache.scala 175:32]
  wire  _GEN_5677 = ~cache_hit ? _GEN_3608 : _GEN_1032; // @[ICache.scala 175:32]
  wire  _GEN_5678 = ~cache_hit ? _GEN_3609 : _GEN_1544; // @[ICache.scala 175:32]
  wire  _GEN_5679 = ~cache_hit ? _GEN_3610 : _GEN_1033; // @[ICache.scala 175:32]
  wire  _GEN_5680 = ~cache_hit ? _GEN_3611 : _GEN_1545; // @[ICache.scala 175:32]
  wire  _GEN_5681 = ~cache_hit ? _GEN_3612 : _GEN_1034; // @[ICache.scala 175:32]
  wire  _GEN_5682 = ~cache_hit ? _GEN_3613 : _GEN_1546; // @[ICache.scala 175:32]
  wire  _GEN_5683 = ~cache_hit ? _GEN_3614 : _GEN_1035; // @[ICache.scala 175:32]
  wire  _GEN_5684 = ~cache_hit ? _GEN_3615 : _GEN_1547; // @[ICache.scala 175:32]
  wire  _GEN_5685 = ~cache_hit ? _GEN_3616 : _GEN_1036; // @[ICache.scala 175:32]
  wire  _GEN_5686 = ~cache_hit ? _GEN_3617 : _GEN_1548; // @[ICache.scala 175:32]
  wire  _GEN_5687 = ~cache_hit ? _GEN_3618 : _GEN_1037; // @[ICache.scala 175:32]
  wire  _GEN_5688 = ~cache_hit ? _GEN_3619 : _GEN_1549; // @[ICache.scala 175:32]
  wire  _GEN_5689 = ~cache_hit ? _GEN_3620 : _GEN_1038; // @[ICache.scala 175:32]
  wire  _GEN_5690 = ~cache_hit ? _GEN_3621 : _GEN_1550; // @[ICache.scala 175:32]
  wire  _GEN_5691 = ~cache_hit ? _GEN_3622 : _GEN_1039; // @[ICache.scala 175:32]
  wire  _GEN_5692 = ~cache_hit ? _GEN_3623 : _GEN_1551; // @[ICache.scala 175:32]
  wire  _GEN_5693 = ~cache_hit ? _GEN_3624 : _GEN_1040; // @[ICache.scala 175:32]
  wire  _GEN_5694 = ~cache_hit ? _GEN_3625 : _GEN_1552; // @[ICache.scala 175:32]
  wire  _GEN_5695 = ~cache_hit ? _GEN_3626 : _GEN_1041; // @[ICache.scala 175:32]
  wire  _GEN_5696 = ~cache_hit ? _GEN_3627 : _GEN_1553; // @[ICache.scala 175:32]
  wire  _GEN_5697 = ~cache_hit ? _GEN_3628 : _GEN_1042; // @[ICache.scala 175:32]
  wire  _GEN_5698 = ~cache_hit ? _GEN_3629 : _GEN_1554; // @[ICache.scala 175:32]
  wire  _GEN_5699 = ~cache_hit ? _GEN_3630 : _GEN_1043; // @[ICache.scala 175:32]
  wire  _GEN_5700 = ~cache_hit ? _GEN_3631 : _GEN_1555; // @[ICache.scala 175:32]
  wire  _GEN_5701 = ~cache_hit ? _GEN_3632 : _GEN_1044; // @[ICache.scala 175:32]
  wire  _GEN_5702 = ~cache_hit ? _GEN_3633 : _GEN_1556; // @[ICache.scala 175:32]
  wire  _GEN_5703 = ~cache_hit ? _GEN_3634 : _GEN_1045; // @[ICache.scala 175:32]
  wire  _GEN_5704 = ~cache_hit ? _GEN_3635 : _GEN_1557; // @[ICache.scala 175:32]
  wire  _GEN_5705 = ~cache_hit ? _GEN_3636 : _GEN_1046; // @[ICache.scala 175:32]
  wire  _GEN_5706 = ~cache_hit ? _GEN_3637 : _GEN_1558; // @[ICache.scala 175:32]
  wire  _GEN_5707 = ~cache_hit ? _GEN_3638 : _GEN_1047; // @[ICache.scala 175:32]
  wire  _GEN_5708 = ~cache_hit ? _GEN_3639 : _GEN_1559; // @[ICache.scala 175:32]
  wire  _GEN_5709 = ~cache_hit ? _GEN_3640 : _GEN_1048; // @[ICache.scala 175:32]
  wire  _GEN_5710 = ~cache_hit ? _GEN_3641 : _GEN_1560; // @[ICache.scala 175:32]
  wire  _GEN_5711 = ~cache_hit ? _GEN_3642 : _GEN_1049; // @[ICache.scala 175:32]
  wire  _GEN_5712 = ~cache_hit ? _GEN_3643 : _GEN_1561; // @[ICache.scala 175:32]
  wire  _GEN_5713 = ~cache_hit ? _GEN_3644 : _GEN_1050; // @[ICache.scala 175:32]
  wire  _GEN_5714 = ~cache_hit ? _GEN_3645 : _GEN_1562; // @[ICache.scala 175:32]
  wire  _GEN_5715 = ~cache_hit ? _GEN_3646 : _GEN_1051; // @[ICache.scala 175:32]
  wire  _GEN_5716 = ~cache_hit ? _GEN_3647 : _GEN_1563; // @[ICache.scala 175:32]
  wire  _GEN_5717 = ~cache_hit ? _GEN_3648 : _GEN_1052; // @[ICache.scala 175:32]
  wire  _GEN_5718 = ~cache_hit ? _GEN_3649 : _GEN_1564; // @[ICache.scala 175:32]
  wire  _GEN_5719 = ~cache_hit ? _GEN_3650 : _GEN_1053; // @[ICache.scala 175:32]
  wire  _GEN_5720 = ~cache_hit ? _GEN_3651 : _GEN_1565; // @[ICache.scala 175:32]
  wire  _GEN_5721 = ~cache_hit ? _GEN_3652 : _GEN_1054; // @[ICache.scala 175:32]
  wire  _GEN_5722 = ~cache_hit ? _GEN_3653 : _GEN_1566; // @[ICache.scala 175:32]
  wire  _GEN_5723 = ~cache_hit ? _GEN_3654 : _GEN_1055; // @[ICache.scala 175:32]
  wire  _GEN_5724 = ~cache_hit ? _GEN_3655 : _GEN_1567; // @[ICache.scala 175:32]
  wire  _GEN_5725 = ~cache_hit ? _GEN_3656 : _GEN_1056; // @[ICache.scala 175:32]
  wire  _GEN_5726 = ~cache_hit ? _GEN_3657 : _GEN_1568; // @[ICache.scala 175:32]
  wire  _GEN_5727 = ~cache_hit ? _GEN_3658 : _GEN_1057; // @[ICache.scala 175:32]
  wire  _GEN_5728 = ~cache_hit ? _GEN_3659 : _GEN_1569; // @[ICache.scala 175:32]
  wire  _GEN_5729 = ~cache_hit ? _GEN_3660 : _GEN_1058; // @[ICache.scala 175:32]
  wire  _GEN_5730 = ~cache_hit ? _GEN_3661 : _GEN_1570; // @[ICache.scala 175:32]
  wire  _GEN_5731 = ~cache_hit ? _GEN_3662 : _GEN_1059; // @[ICache.scala 175:32]
  wire  _GEN_5732 = ~cache_hit ? _GEN_3663 : _GEN_1571; // @[ICache.scala 175:32]
  wire  _GEN_5733 = ~cache_hit ? _GEN_3664 : _GEN_1060; // @[ICache.scala 175:32]
  wire  _GEN_5734 = ~cache_hit ? _GEN_3665 : _GEN_1572; // @[ICache.scala 175:32]
  wire  _GEN_5735 = ~cache_hit ? _GEN_3666 : _GEN_1061; // @[ICache.scala 175:32]
  wire  _GEN_5736 = ~cache_hit ? _GEN_3667 : _GEN_1573; // @[ICache.scala 175:32]
  wire  _GEN_5737 = ~cache_hit ? _GEN_3668 : _GEN_1062; // @[ICache.scala 175:32]
  wire  _GEN_5738 = ~cache_hit ? _GEN_3669 : _GEN_1574; // @[ICache.scala 175:32]
  wire  _GEN_5739 = ~cache_hit ? _GEN_3670 : _GEN_1063; // @[ICache.scala 175:32]
  wire  _GEN_5740 = ~cache_hit ? _GEN_3671 : _GEN_1575; // @[ICache.scala 175:32]
  wire  _GEN_5741 = ~cache_hit ? _GEN_3672 : _GEN_1064; // @[ICache.scala 175:32]
  wire  _GEN_5742 = ~cache_hit ? _GEN_3673 : _GEN_1576; // @[ICache.scala 175:32]
  wire  _GEN_5743 = ~cache_hit ? _GEN_3674 : _GEN_1065; // @[ICache.scala 175:32]
  wire  _GEN_5744 = ~cache_hit ? _GEN_3675 : _GEN_1577; // @[ICache.scala 175:32]
  wire  _GEN_5745 = ~cache_hit ? _GEN_3676 : _GEN_1066; // @[ICache.scala 175:32]
  wire  _GEN_5746 = ~cache_hit ? _GEN_3677 : _GEN_1578; // @[ICache.scala 175:32]
  wire  _GEN_5747 = ~cache_hit ? _GEN_3678 : _GEN_1067; // @[ICache.scala 175:32]
  wire  _GEN_5748 = ~cache_hit ? _GEN_3679 : _GEN_1579; // @[ICache.scala 175:32]
  wire  _GEN_5749 = ~cache_hit ? _GEN_3680 : _GEN_1068; // @[ICache.scala 175:32]
  wire  _GEN_5750 = ~cache_hit ? _GEN_3681 : _GEN_1580; // @[ICache.scala 175:32]
  wire  _GEN_5751 = ~cache_hit ? _GEN_3682 : _GEN_1069; // @[ICache.scala 175:32]
  wire  _GEN_5752 = ~cache_hit ? _GEN_3683 : _GEN_1581; // @[ICache.scala 175:32]
  wire  _GEN_5753 = ~cache_hit ? _GEN_3684 : _GEN_1070; // @[ICache.scala 175:32]
  wire  _GEN_5754 = ~cache_hit ? _GEN_3685 : _GEN_1582; // @[ICache.scala 175:32]
  wire  _GEN_5755 = ~cache_hit ? _GEN_3686 : _GEN_1071; // @[ICache.scala 175:32]
  wire  _GEN_5756 = ~cache_hit ? _GEN_3687 : _GEN_1583; // @[ICache.scala 175:32]
  wire  _GEN_5757 = ~cache_hit ? _GEN_3688 : _GEN_1072; // @[ICache.scala 175:32]
  wire  _GEN_5758 = ~cache_hit ? _GEN_3689 : _GEN_1584; // @[ICache.scala 175:32]
  wire  _GEN_5759 = ~cache_hit ? _GEN_3690 : _GEN_1073; // @[ICache.scala 175:32]
  wire  _GEN_5760 = ~cache_hit ? _GEN_3691 : _GEN_1585; // @[ICache.scala 175:32]
  wire  _GEN_5761 = ~cache_hit ? _GEN_3692 : _GEN_1074; // @[ICache.scala 175:32]
  wire  _GEN_5762 = ~cache_hit ? _GEN_3693 : _GEN_1586; // @[ICache.scala 175:32]
  wire  _GEN_5763 = ~cache_hit ? _GEN_3694 : _GEN_1075; // @[ICache.scala 175:32]
  wire  _GEN_5764 = ~cache_hit ? _GEN_3695 : _GEN_1587; // @[ICache.scala 175:32]
  wire  _GEN_5765 = ~cache_hit ? _GEN_3696 : _GEN_1076; // @[ICache.scala 175:32]
  wire  _GEN_5766 = ~cache_hit ? _GEN_3697 : _GEN_1588; // @[ICache.scala 175:32]
  wire  _GEN_5767 = ~cache_hit ? _GEN_3698 : _GEN_1077; // @[ICache.scala 175:32]
  wire  _GEN_5768 = ~cache_hit ? _GEN_3699 : _GEN_1589; // @[ICache.scala 175:32]
  wire  _GEN_5769 = ~cache_hit ? _GEN_3700 : _GEN_1078; // @[ICache.scala 175:32]
  wire  _GEN_5770 = ~cache_hit ? _GEN_3701 : _GEN_1590; // @[ICache.scala 175:32]
  wire  _GEN_5771 = ~cache_hit ? _GEN_3702 : _GEN_1079; // @[ICache.scala 175:32]
  wire  _GEN_5772 = ~cache_hit ? _GEN_3703 : _GEN_1591; // @[ICache.scala 175:32]
  wire  _GEN_5773 = ~cache_hit ? _GEN_3704 : _GEN_1080; // @[ICache.scala 175:32]
  wire  _GEN_5774 = ~cache_hit ? _GEN_3705 : _GEN_1592; // @[ICache.scala 175:32]
  wire  _GEN_5775 = ~cache_hit ? _GEN_3706 : _GEN_1081; // @[ICache.scala 175:32]
  wire  _GEN_5776 = ~cache_hit ? _GEN_3707 : _GEN_1593; // @[ICache.scala 175:32]
  wire  _GEN_5777 = ~cache_hit ? _GEN_3708 : _GEN_1082; // @[ICache.scala 175:32]
  wire  _GEN_5778 = ~cache_hit ? _GEN_3709 : _GEN_1594; // @[ICache.scala 175:32]
  wire  _GEN_5779 = ~cache_hit ? _GEN_3710 : _GEN_1083; // @[ICache.scala 175:32]
  wire  _GEN_5780 = ~cache_hit ? _GEN_3711 : _GEN_1595; // @[ICache.scala 175:32]
  wire  _GEN_5781 = ~cache_hit ? _GEN_3712 : _GEN_1084; // @[ICache.scala 175:32]
  wire  _GEN_5782 = ~cache_hit ? _GEN_3713 : _GEN_1596; // @[ICache.scala 175:32]
  wire  _GEN_5783 = ~cache_hit ? _GEN_3714 : _GEN_1085; // @[ICache.scala 175:32]
  wire  _GEN_5784 = ~cache_hit ? _GEN_3715 : _GEN_1597; // @[ICache.scala 175:32]
  wire  _GEN_5785 = ~cache_hit ? _GEN_3716 : _GEN_1086; // @[ICache.scala 175:32]
  wire  _GEN_5786 = ~cache_hit ? _GEN_3717 : _GEN_1598; // @[ICache.scala 175:32]
  wire  _GEN_5787 = ~cache_hit ? _GEN_3718 : _GEN_1087; // @[ICache.scala 175:32]
  wire  _GEN_5788 = ~cache_hit ? _GEN_3719 : _GEN_1599; // @[ICache.scala 175:32]
  wire  _GEN_5789 = ~cache_hit ? _GEN_3720 : _GEN_1088; // @[ICache.scala 175:32]
  wire  _GEN_5790 = ~cache_hit ? _GEN_3721 : _GEN_1600; // @[ICache.scala 175:32]
  wire  _GEN_5791 = ~cache_hit ? _GEN_3722 : _GEN_1089; // @[ICache.scala 175:32]
  wire  _GEN_5792 = ~cache_hit ? _GEN_3723 : _GEN_1601; // @[ICache.scala 175:32]
  wire  _GEN_5793 = ~cache_hit ? _GEN_3724 : _GEN_1090; // @[ICache.scala 175:32]
  wire  _GEN_5794 = ~cache_hit ? _GEN_3725 : _GEN_1602; // @[ICache.scala 175:32]
  wire  _GEN_5795 = ~cache_hit ? _GEN_3726 : _GEN_1091; // @[ICache.scala 175:32]
  wire  _GEN_5796 = ~cache_hit ? _GEN_3727 : _GEN_1603; // @[ICache.scala 175:32]
  wire  _GEN_5797 = ~cache_hit ? _GEN_3728 : _GEN_1092; // @[ICache.scala 175:32]
  wire  _GEN_5798 = ~cache_hit ? _GEN_3729 : _GEN_1604; // @[ICache.scala 175:32]
  wire  _GEN_5799 = ~cache_hit ? _GEN_3730 : _GEN_1093; // @[ICache.scala 175:32]
  wire  _GEN_5800 = ~cache_hit ? _GEN_3731 : _GEN_1605; // @[ICache.scala 175:32]
  wire  _GEN_5801 = ~cache_hit ? _GEN_3732 : _GEN_1094; // @[ICache.scala 175:32]
  wire  _GEN_5802 = ~cache_hit ? _GEN_3733 : _GEN_1606; // @[ICache.scala 175:32]
  wire  _GEN_5803 = ~cache_hit ? _GEN_3734 : _GEN_1095; // @[ICache.scala 175:32]
  wire  _GEN_5804 = ~cache_hit ? _GEN_3735 : _GEN_1607; // @[ICache.scala 175:32]
  wire  _GEN_5805 = ~cache_hit ? _GEN_3736 : _GEN_1096; // @[ICache.scala 175:32]
  wire  _GEN_5806 = ~cache_hit ? _GEN_3737 : _GEN_1608; // @[ICache.scala 175:32]
  wire  _GEN_5807 = ~cache_hit ? _GEN_3738 : _GEN_1097; // @[ICache.scala 175:32]
  wire  _GEN_5808 = ~cache_hit ? _GEN_3739 : _GEN_1609; // @[ICache.scala 175:32]
  wire  _GEN_5809 = ~cache_hit ? _GEN_3740 : _GEN_1098; // @[ICache.scala 175:32]
  wire  _GEN_5810 = ~cache_hit ? _GEN_3741 : _GEN_1610; // @[ICache.scala 175:32]
  wire  _GEN_5811 = ~cache_hit ? _GEN_3742 : _GEN_1099; // @[ICache.scala 175:32]
  wire  _GEN_5812 = ~cache_hit ? _GEN_3743 : _GEN_1611; // @[ICache.scala 175:32]
  wire  _GEN_5813 = ~cache_hit ? _GEN_3744 : _GEN_1100; // @[ICache.scala 175:32]
  wire  _GEN_5814 = ~cache_hit ? _GEN_3745 : _GEN_1612; // @[ICache.scala 175:32]
  wire  _GEN_5815 = ~cache_hit ? _GEN_3746 : _GEN_1101; // @[ICache.scala 175:32]
  wire  _GEN_5816 = ~cache_hit ? _GEN_3747 : _GEN_1613; // @[ICache.scala 175:32]
  wire  _GEN_5817 = ~cache_hit ? _GEN_3748 : _GEN_1102; // @[ICache.scala 175:32]
  wire  _GEN_5818 = ~cache_hit ? _GEN_3749 : _GEN_1614; // @[ICache.scala 175:32]
  wire  _GEN_5819 = ~cache_hit ? _GEN_3750 : _GEN_1103; // @[ICache.scala 175:32]
  wire  _GEN_5820 = ~cache_hit ? _GEN_3751 : _GEN_1615; // @[ICache.scala 175:32]
  wire  _GEN_5821 = ~cache_hit ? _GEN_3752 : _GEN_1104; // @[ICache.scala 175:32]
  wire  _GEN_5822 = ~cache_hit ? _GEN_3753 : _GEN_1616; // @[ICache.scala 175:32]
  wire  _GEN_5823 = ~cache_hit ? _GEN_3754 : _GEN_1105; // @[ICache.scala 175:32]
  wire  _GEN_5824 = ~cache_hit ? _GEN_3755 : _GEN_1617; // @[ICache.scala 175:32]
  wire  _GEN_5825 = ~cache_hit ? _GEN_3756 : _GEN_1106; // @[ICache.scala 175:32]
  wire  _GEN_5826 = ~cache_hit ? _GEN_3757 : _GEN_1618; // @[ICache.scala 175:32]
  wire  _GEN_5827 = ~cache_hit ? _GEN_3758 : _GEN_1107; // @[ICache.scala 175:32]
  wire  _GEN_5828 = ~cache_hit ? _GEN_3759 : _GEN_1619; // @[ICache.scala 175:32]
  wire  _GEN_5829 = ~cache_hit ? _GEN_3760 : _GEN_1108; // @[ICache.scala 175:32]
  wire  _GEN_5830 = ~cache_hit ? _GEN_3761 : _GEN_1620; // @[ICache.scala 175:32]
  wire  _GEN_5831 = ~cache_hit ? _GEN_3762 : _GEN_1109; // @[ICache.scala 175:32]
  wire  _GEN_5832 = ~cache_hit ? _GEN_3763 : _GEN_1621; // @[ICache.scala 175:32]
  wire  _GEN_5833 = ~cache_hit ? _GEN_3764 : _GEN_1110; // @[ICache.scala 175:32]
  wire  _GEN_5834 = ~cache_hit ? _GEN_3765 : _GEN_1622; // @[ICache.scala 175:32]
  wire  _GEN_5835 = ~cache_hit ? _GEN_3766 : _GEN_1111; // @[ICache.scala 175:32]
  wire  _GEN_5836 = ~cache_hit ? _GEN_3767 : _GEN_1623; // @[ICache.scala 175:32]
  wire  _GEN_5837 = ~cache_hit ? _GEN_3768 : _GEN_1112; // @[ICache.scala 175:32]
  wire  _GEN_5838 = ~cache_hit ? _GEN_3769 : _GEN_1624; // @[ICache.scala 175:32]
  wire  _GEN_5839 = ~cache_hit ? _GEN_3770 : _GEN_1113; // @[ICache.scala 175:32]
  wire  _GEN_5840 = ~cache_hit ? _GEN_3771 : _GEN_1625; // @[ICache.scala 175:32]
  wire  _GEN_5841 = ~cache_hit ? _GEN_3772 : _GEN_1114; // @[ICache.scala 175:32]
  wire  _GEN_5842 = ~cache_hit ? _GEN_3773 : _GEN_1626; // @[ICache.scala 175:32]
  wire  _GEN_5843 = ~cache_hit ? _GEN_3774 : _GEN_1115; // @[ICache.scala 175:32]
  wire  _GEN_5844 = ~cache_hit ? _GEN_3775 : _GEN_1627; // @[ICache.scala 175:32]
  wire  _GEN_5845 = ~cache_hit ? _GEN_3776 : _GEN_1116; // @[ICache.scala 175:32]
  wire  _GEN_5846 = ~cache_hit ? _GEN_3777 : _GEN_1628; // @[ICache.scala 175:32]
  wire  _GEN_5847 = ~cache_hit ? _GEN_3778 : _GEN_1117; // @[ICache.scala 175:32]
  wire  _GEN_5848 = ~cache_hit ? _GEN_3779 : _GEN_1629; // @[ICache.scala 175:32]
  wire  _GEN_5849 = ~cache_hit ? _GEN_3780 : _GEN_1118; // @[ICache.scala 175:32]
  wire  _GEN_5850 = ~cache_hit ? _GEN_3781 : _GEN_1630; // @[ICache.scala 175:32]
  wire  _GEN_5851 = ~cache_hit ? _GEN_3782 : _GEN_1119; // @[ICache.scala 175:32]
  wire  _GEN_5852 = ~cache_hit ? _GEN_3783 : _GEN_1631; // @[ICache.scala 175:32]
  wire  _GEN_5853 = ~cache_hit ? _GEN_3784 : _GEN_1120; // @[ICache.scala 175:32]
  wire  _GEN_5854 = ~cache_hit ? _GEN_3785 : _GEN_1632; // @[ICache.scala 175:32]
  wire  _GEN_5855 = ~cache_hit ? _GEN_3786 : _GEN_1121; // @[ICache.scala 175:32]
  wire  _GEN_5856 = ~cache_hit ? _GEN_3787 : _GEN_1633; // @[ICache.scala 175:32]
  wire  _GEN_5857 = ~cache_hit ? _GEN_3788 : _GEN_1122; // @[ICache.scala 175:32]
  wire  _GEN_5858 = ~cache_hit ? _GEN_3789 : _GEN_1634; // @[ICache.scala 175:32]
  wire  _GEN_5859 = ~cache_hit ? _GEN_3790 : _GEN_1123; // @[ICache.scala 175:32]
  wire  _GEN_5860 = ~cache_hit ? _GEN_3791 : _GEN_1635; // @[ICache.scala 175:32]
  wire  _GEN_5861 = ~cache_hit ? _GEN_3792 : _GEN_1124; // @[ICache.scala 175:32]
  wire  _GEN_5862 = ~cache_hit ? _GEN_3793 : _GEN_1636; // @[ICache.scala 175:32]
  wire  _GEN_5863 = ~cache_hit ? _GEN_3794 : _GEN_1125; // @[ICache.scala 175:32]
  wire  _GEN_5864 = ~cache_hit ? _GEN_3795 : _GEN_1637; // @[ICache.scala 175:32]
  wire  _GEN_5865 = ~cache_hit ? _GEN_3796 : _GEN_1126; // @[ICache.scala 175:32]
  wire  _GEN_5866 = ~cache_hit ? _GEN_3797 : _GEN_1638; // @[ICache.scala 175:32]
  wire  _GEN_5867 = ~cache_hit ? _GEN_3798 : _GEN_1127; // @[ICache.scala 175:32]
  wire  _GEN_5868 = ~cache_hit ? _GEN_3799 : _GEN_1639; // @[ICache.scala 175:32]
  wire  _GEN_5869 = ~cache_hit ? _GEN_3800 : _GEN_1128; // @[ICache.scala 175:32]
  wire  _GEN_5870 = ~cache_hit ? _GEN_3801 : _GEN_1640; // @[ICache.scala 175:32]
  wire  _GEN_5871 = ~cache_hit ? _GEN_3802 : _GEN_1129; // @[ICache.scala 175:32]
  wire  _GEN_5872 = ~cache_hit ? _GEN_3803 : _GEN_1641; // @[ICache.scala 175:32]
  wire  _GEN_5873 = ~cache_hit ? _GEN_3804 : _GEN_1130; // @[ICache.scala 175:32]
  wire  _GEN_5874 = ~cache_hit ? _GEN_3805 : _GEN_1642; // @[ICache.scala 175:32]
  wire  _GEN_5875 = ~cache_hit ? _GEN_3806 : _GEN_1131; // @[ICache.scala 175:32]
  wire  _GEN_5876 = ~cache_hit ? _GEN_3807 : _GEN_1643; // @[ICache.scala 175:32]
  wire  _GEN_5877 = ~cache_hit ? _GEN_3808 : _GEN_1132; // @[ICache.scala 175:32]
  wire  _GEN_5878 = ~cache_hit ? _GEN_3809 : _GEN_1644; // @[ICache.scala 175:32]
  wire  _GEN_5879 = ~cache_hit ? _GEN_3810 : _GEN_1133; // @[ICache.scala 175:32]
  wire  _GEN_5880 = ~cache_hit ? _GEN_3811 : _GEN_1645; // @[ICache.scala 175:32]
  wire  _GEN_5881 = ~cache_hit ? _GEN_3812 : _GEN_1134; // @[ICache.scala 175:32]
  wire  _GEN_5882 = ~cache_hit ? _GEN_3813 : _GEN_1646; // @[ICache.scala 175:32]
  wire  _GEN_5883 = ~cache_hit ? _GEN_3814 : _GEN_1135; // @[ICache.scala 175:32]
  wire  _GEN_5884 = ~cache_hit ? _GEN_3815 : _GEN_1647; // @[ICache.scala 175:32]
  wire  _GEN_5885 = ~cache_hit ? _GEN_3816 : _GEN_1136; // @[ICache.scala 175:32]
  wire  _GEN_5886 = ~cache_hit ? _GEN_3817 : _GEN_1648; // @[ICache.scala 175:32]
  wire  _GEN_5887 = ~cache_hit ? _GEN_3818 : _GEN_1137; // @[ICache.scala 175:32]
  wire  _GEN_5888 = ~cache_hit ? _GEN_3819 : _GEN_1649; // @[ICache.scala 175:32]
  wire  _GEN_5889 = ~cache_hit ? _GEN_3820 : _GEN_1138; // @[ICache.scala 175:32]
  wire  _GEN_5890 = ~cache_hit ? _GEN_3821 : _GEN_1650; // @[ICache.scala 175:32]
  wire  _GEN_5891 = ~cache_hit ? _GEN_3822 : _GEN_1139; // @[ICache.scala 175:32]
  wire  _GEN_5892 = ~cache_hit ? _GEN_3823 : _GEN_1651; // @[ICache.scala 175:32]
  wire  _GEN_5893 = ~cache_hit ? _GEN_3824 : _GEN_1140; // @[ICache.scala 175:32]
  wire  _GEN_5894 = ~cache_hit ? _GEN_3825 : _GEN_1652; // @[ICache.scala 175:32]
  wire  _GEN_5895 = ~cache_hit ? _GEN_3826 : _GEN_1141; // @[ICache.scala 175:32]
  wire  _GEN_5896 = ~cache_hit ? _GEN_3827 : _GEN_1653; // @[ICache.scala 175:32]
  wire  _GEN_5897 = ~cache_hit ? _GEN_3828 : _GEN_1142; // @[ICache.scala 175:32]
  wire  _GEN_5898 = ~cache_hit ? _GEN_3829 : _GEN_1654; // @[ICache.scala 175:32]
  wire  _GEN_5899 = ~cache_hit ? _GEN_3830 : _GEN_1143; // @[ICache.scala 175:32]
  wire  _GEN_5900 = ~cache_hit ? _GEN_3831 : _GEN_1655; // @[ICache.scala 175:32]
  wire  _GEN_5901 = ~cache_hit ? _GEN_3832 : _GEN_1144; // @[ICache.scala 175:32]
  wire  _GEN_5902 = ~cache_hit ? _GEN_3833 : _GEN_1656; // @[ICache.scala 175:32]
  wire  _GEN_5903 = ~cache_hit ? _GEN_3834 : _GEN_1145; // @[ICache.scala 175:32]
  wire  _GEN_5904 = ~cache_hit ? _GEN_3835 : _GEN_1657; // @[ICache.scala 175:32]
  wire  _GEN_5905 = ~cache_hit ? _GEN_3836 : _GEN_1146; // @[ICache.scala 175:32]
  wire  _GEN_5906 = ~cache_hit ? _GEN_3837 : _GEN_1658; // @[ICache.scala 175:32]
  wire  _GEN_5907 = ~cache_hit ? _GEN_3838 : _GEN_1147; // @[ICache.scala 175:32]
  wire  _GEN_5908 = ~cache_hit ? _GEN_3839 : _GEN_1659; // @[ICache.scala 175:32]
  wire  _GEN_5909 = ~cache_hit ? _GEN_3840 : _GEN_1148; // @[ICache.scala 175:32]
  wire  _GEN_5910 = ~cache_hit ? _GEN_3841 : _GEN_1660; // @[ICache.scala 175:32]
  wire  _GEN_5911 = ~cache_hit ? _GEN_3842 : _GEN_1149; // @[ICache.scala 175:32]
  wire  _GEN_5912 = ~cache_hit ? _GEN_3843 : _GEN_1661; // @[ICache.scala 175:32]
  wire  _GEN_5913 = ~cache_hit ? _GEN_3844 : _GEN_1150; // @[ICache.scala 175:32]
  wire  _GEN_5914 = ~cache_hit ? _GEN_3845 : _GEN_1662; // @[ICache.scala 175:32]
  wire  _GEN_5915 = ~cache_hit ? _GEN_3846 : _GEN_1151; // @[ICache.scala 175:32]
  wire  _GEN_5916 = ~cache_hit ? _GEN_3847 : _GEN_1663; // @[ICache.scala 175:32]
  wire  _GEN_5917 = ~cache_hit ? _GEN_3848 : _GEN_1152; // @[ICache.scala 175:32]
  wire  _GEN_5918 = ~cache_hit ? _GEN_3849 : _GEN_1664; // @[ICache.scala 175:32]
  wire  _GEN_5919 = ~cache_hit ? _GEN_3850 : _GEN_1153; // @[ICache.scala 175:32]
  wire  _GEN_5920 = ~cache_hit ? _GEN_3851 : _GEN_1665; // @[ICache.scala 175:32]
  wire  _GEN_5921 = ~cache_hit ? _GEN_3852 : _GEN_1154; // @[ICache.scala 175:32]
  wire  _GEN_5922 = ~cache_hit ? _GEN_3853 : _GEN_1666; // @[ICache.scala 175:32]
  wire  _GEN_5923 = ~cache_hit ? _GEN_3854 : _GEN_1155; // @[ICache.scala 175:32]
  wire  _GEN_5924 = ~cache_hit ? _GEN_3855 : _GEN_1667; // @[ICache.scala 175:32]
  wire  _GEN_5925 = ~cache_hit ? _GEN_3856 : _GEN_1156; // @[ICache.scala 175:32]
  wire  _GEN_5926 = ~cache_hit ? _GEN_3857 : _GEN_1668; // @[ICache.scala 175:32]
  wire  _GEN_5927 = ~cache_hit ? _GEN_3858 : _GEN_1157; // @[ICache.scala 175:32]
  wire  _GEN_5928 = ~cache_hit ? _GEN_3859 : _GEN_1669; // @[ICache.scala 175:32]
  wire  _GEN_5929 = ~cache_hit ? _GEN_3860 : _GEN_1158; // @[ICache.scala 175:32]
  wire  _GEN_5930 = ~cache_hit ? _GEN_3861 : _GEN_1670; // @[ICache.scala 175:32]
  wire  _GEN_5931 = ~cache_hit ? _GEN_3862 : _GEN_1159; // @[ICache.scala 175:32]
  wire  _GEN_5932 = ~cache_hit ? _GEN_3863 : _GEN_1671; // @[ICache.scala 175:32]
  wire  _GEN_5933 = ~cache_hit ? _GEN_3864 : _GEN_1160; // @[ICache.scala 175:32]
  wire  _GEN_5934 = ~cache_hit ? _GEN_3865 : _GEN_1672; // @[ICache.scala 175:32]
  wire  _GEN_5935 = ~cache_hit ? _GEN_3866 : _GEN_1161; // @[ICache.scala 175:32]
  wire  _GEN_5936 = ~cache_hit ? _GEN_3867 : _GEN_1673; // @[ICache.scala 175:32]
  wire  _GEN_5937 = ~cache_hit ? _GEN_3868 : _GEN_1162; // @[ICache.scala 175:32]
  wire  _GEN_5938 = ~cache_hit ? _GEN_3869 : _GEN_1674; // @[ICache.scala 175:32]
  wire  _GEN_5939 = ~cache_hit ? _GEN_3870 : _GEN_1163; // @[ICache.scala 175:32]
  wire  _GEN_5940 = ~cache_hit ? _GEN_3871 : _GEN_1675; // @[ICache.scala 175:32]
  wire  _GEN_5941 = ~cache_hit ? _GEN_3872 : _GEN_1164; // @[ICache.scala 175:32]
  wire  _GEN_5942 = ~cache_hit ? _GEN_3873 : _GEN_1676; // @[ICache.scala 175:32]
  wire  _GEN_5943 = ~cache_hit ? _GEN_3874 : _GEN_1165; // @[ICache.scala 175:32]
  wire  _GEN_5944 = ~cache_hit ? _GEN_3875 : _GEN_1677; // @[ICache.scala 175:32]
  wire  _GEN_5945 = ~cache_hit ? _GEN_3876 : _GEN_1166; // @[ICache.scala 175:32]
  wire  _GEN_5946 = ~cache_hit ? _GEN_3877 : _GEN_1678; // @[ICache.scala 175:32]
  wire  _GEN_5947 = ~cache_hit ? _GEN_3878 : _GEN_1167; // @[ICache.scala 175:32]
  wire  _GEN_5948 = ~cache_hit ? _GEN_3879 : _GEN_1679; // @[ICache.scala 175:32]
  wire  _GEN_5949 = ~cache_hit ? _GEN_3880 : _GEN_1168; // @[ICache.scala 175:32]
  wire  _GEN_5950 = ~cache_hit ? _GEN_3881 : _GEN_1680; // @[ICache.scala 175:32]
  wire  _GEN_5951 = ~cache_hit ? _GEN_3882 : _GEN_1169; // @[ICache.scala 175:32]
  wire  _GEN_5952 = ~cache_hit ? _GEN_3883 : _GEN_1681; // @[ICache.scala 175:32]
  wire  _GEN_5953 = ~cache_hit ? _GEN_3884 : _GEN_1170; // @[ICache.scala 175:32]
  wire  _GEN_5954 = ~cache_hit ? _GEN_3885 : _GEN_1682; // @[ICache.scala 175:32]
  wire  _GEN_5955 = ~cache_hit ? _GEN_3886 : _GEN_1171; // @[ICache.scala 175:32]
  wire  _GEN_5956 = ~cache_hit ? _GEN_3887 : _GEN_1683; // @[ICache.scala 175:32]
  wire  _GEN_5957 = ~cache_hit ? _GEN_3888 : _GEN_1172; // @[ICache.scala 175:32]
  wire  _GEN_5958 = ~cache_hit ? _GEN_3889 : _GEN_1684; // @[ICache.scala 175:32]
  wire  _GEN_5959 = ~cache_hit ? _GEN_3890 : _GEN_1173; // @[ICache.scala 175:32]
  wire  _GEN_5960 = ~cache_hit ? _GEN_3891 : _GEN_1685; // @[ICache.scala 175:32]
  wire  _GEN_5961 = ~cache_hit ? _GEN_3892 : _GEN_1174; // @[ICache.scala 175:32]
  wire  _GEN_5962 = ~cache_hit ? _GEN_3893 : _GEN_1686; // @[ICache.scala 175:32]
  wire  _GEN_5963 = ~cache_hit ? _GEN_3894 : _GEN_1175; // @[ICache.scala 175:32]
  wire  _GEN_5964 = ~cache_hit ? _GEN_3895 : _GEN_1687; // @[ICache.scala 175:32]
  wire  _GEN_5965 = ~cache_hit ? _GEN_3896 : _GEN_1176; // @[ICache.scala 175:32]
  wire  _GEN_5966 = ~cache_hit ? _GEN_3897 : _GEN_1688; // @[ICache.scala 175:32]
  wire  _GEN_5967 = ~cache_hit ? _GEN_3898 : _GEN_1177; // @[ICache.scala 175:32]
  wire  _GEN_5968 = ~cache_hit ? _GEN_3899 : _GEN_1689; // @[ICache.scala 175:32]
  wire  _GEN_5969 = ~cache_hit ? _GEN_3900 : _GEN_1178; // @[ICache.scala 175:32]
  wire  _GEN_5970 = ~cache_hit ? _GEN_3901 : _GEN_1690; // @[ICache.scala 175:32]
  wire  _GEN_5971 = ~cache_hit ? _GEN_3902 : _GEN_1179; // @[ICache.scala 175:32]
  wire  _GEN_5972 = ~cache_hit ? _GEN_3903 : _GEN_1691; // @[ICache.scala 175:32]
  wire  _GEN_5973 = ~cache_hit ? _GEN_3904 : _GEN_1180; // @[ICache.scala 175:32]
  wire  _GEN_5974 = ~cache_hit ? _GEN_3905 : _GEN_1692; // @[ICache.scala 175:32]
  wire  _GEN_5975 = ~cache_hit ? _GEN_3906 : _GEN_1181; // @[ICache.scala 175:32]
  wire  _GEN_5976 = ~cache_hit ? _GEN_3907 : _GEN_1693; // @[ICache.scala 175:32]
  wire  _GEN_5977 = ~cache_hit ? _GEN_3908 : _GEN_1182; // @[ICache.scala 175:32]
  wire  _GEN_5978 = ~cache_hit ? _GEN_3909 : _GEN_1694; // @[ICache.scala 175:32]
  wire  _GEN_5979 = ~cache_hit ? _GEN_3910 : _GEN_1183; // @[ICache.scala 175:32]
  wire  _GEN_5980 = ~cache_hit ? _GEN_3911 : _GEN_1695; // @[ICache.scala 175:32]
  wire  _GEN_5981 = ~cache_hit ? _GEN_3912 : _GEN_1184; // @[ICache.scala 175:32]
  wire  _GEN_5982 = ~cache_hit ? _GEN_3913 : _GEN_1696; // @[ICache.scala 175:32]
  wire  _GEN_5983 = ~cache_hit ? _GEN_3914 : _GEN_1185; // @[ICache.scala 175:32]
  wire  _GEN_5984 = ~cache_hit ? _GEN_3915 : _GEN_1697; // @[ICache.scala 175:32]
  wire  _GEN_5985 = ~cache_hit ? _GEN_3916 : _GEN_1186; // @[ICache.scala 175:32]
  wire  _GEN_5986 = ~cache_hit ? _GEN_3917 : _GEN_1698; // @[ICache.scala 175:32]
  wire  _GEN_5987 = ~cache_hit ? _GEN_3918 : _GEN_1187; // @[ICache.scala 175:32]
  wire  _GEN_5988 = ~cache_hit ? _GEN_3919 : _GEN_1699; // @[ICache.scala 175:32]
  wire  _GEN_5989 = ~cache_hit ? _GEN_3920 : _GEN_1188; // @[ICache.scala 175:32]
  wire  _GEN_5990 = ~cache_hit ? _GEN_3921 : _GEN_1700; // @[ICache.scala 175:32]
  wire  _GEN_5991 = ~cache_hit ? _GEN_3922 : _GEN_1189; // @[ICache.scala 175:32]
  wire  _GEN_5992 = ~cache_hit ? _GEN_3923 : _GEN_1701; // @[ICache.scala 175:32]
  wire  _GEN_5993 = ~cache_hit ? _GEN_3924 : _GEN_1190; // @[ICache.scala 175:32]
  wire  _GEN_5994 = ~cache_hit ? _GEN_3925 : _GEN_1702; // @[ICache.scala 175:32]
  wire  _GEN_5995 = ~cache_hit ? _GEN_3926 : _GEN_1191; // @[ICache.scala 175:32]
  wire  _GEN_5996 = ~cache_hit ? _GEN_3927 : _GEN_1703; // @[ICache.scala 175:32]
  wire  _GEN_5997 = ~cache_hit ? _GEN_3928 : _GEN_1192; // @[ICache.scala 175:32]
  wire  _GEN_5998 = ~cache_hit ? _GEN_3929 : _GEN_1704; // @[ICache.scala 175:32]
  wire  _GEN_5999 = ~cache_hit ? _GEN_3930 : _GEN_1193; // @[ICache.scala 175:32]
  wire  _GEN_6000 = ~cache_hit ? _GEN_3931 : _GEN_1705; // @[ICache.scala 175:32]
  wire  _GEN_6001 = ~cache_hit ? _GEN_3932 : _GEN_1194; // @[ICache.scala 175:32]
  wire  _GEN_6002 = ~cache_hit ? _GEN_3933 : _GEN_1706; // @[ICache.scala 175:32]
  wire  _GEN_6003 = ~cache_hit ? _GEN_3934 : _GEN_1195; // @[ICache.scala 175:32]
  wire  _GEN_6004 = ~cache_hit ? _GEN_3935 : _GEN_1707; // @[ICache.scala 175:32]
  wire  _GEN_6005 = ~cache_hit ? _GEN_3936 : _GEN_1196; // @[ICache.scala 175:32]
  wire  _GEN_6006 = ~cache_hit ? _GEN_3937 : _GEN_1708; // @[ICache.scala 175:32]
  wire  _GEN_6007 = ~cache_hit ? _GEN_3938 : _GEN_1197; // @[ICache.scala 175:32]
  wire  _GEN_6008 = ~cache_hit ? _GEN_3939 : _GEN_1709; // @[ICache.scala 175:32]
  wire  _GEN_6009 = ~cache_hit ? _GEN_3940 : _GEN_1198; // @[ICache.scala 175:32]
  wire  _GEN_6010 = ~cache_hit ? _GEN_3941 : _GEN_1710; // @[ICache.scala 175:32]
  wire  _GEN_6011 = ~cache_hit ? _GEN_3942 : _GEN_1199; // @[ICache.scala 175:32]
  wire  _GEN_6012 = ~cache_hit ? _GEN_3943 : _GEN_1711; // @[ICache.scala 175:32]
  wire  _GEN_6013 = ~cache_hit ? _GEN_3944 : _GEN_1200; // @[ICache.scala 175:32]
  wire  _GEN_6014 = ~cache_hit ? _GEN_3945 : _GEN_1712; // @[ICache.scala 175:32]
  wire  _GEN_6015 = ~cache_hit ? _GEN_3946 : _GEN_1201; // @[ICache.scala 175:32]
  wire  _GEN_6016 = ~cache_hit ? _GEN_3947 : _GEN_1713; // @[ICache.scala 175:32]
  wire  _GEN_6017 = ~cache_hit ? _GEN_3948 : _GEN_1202; // @[ICache.scala 175:32]
  wire  _GEN_6018 = ~cache_hit ? _GEN_3949 : _GEN_1714; // @[ICache.scala 175:32]
  wire  _GEN_6019 = ~cache_hit ? _GEN_3950 : _GEN_1203; // @[ICache.scala 175:32]
  wire  _GEN_6020 = ~cache_hit ? _GEN_3951 : _GEN_1715; // @[ICache.scala 175:32]
  wire  _GEN_6021 = ~cache_hit ? _GEN_3952 : _GEN_1204; // @[ICache.scala 175:32]
  wire  _GEN_6022 = ~cache_hit ? _GEN_3953 : _GEN_1716; // @[ICache.scala 175:32]
  wire  _GEN_6023 = ~cache_hit ? _GEN_3954 : _GEN_1205; // @[ICache.scala 175:32]
  wire  _GEN_6024 = ~cache_hit ? _GEN_3955 : _GEN_1717; // @[ICache.scala 175:32]
  wire  _GEN_6025 = ~cache_hit ? _GEN_3956 : _GEN_1206; // @[ICache.scala 175:32]
  wire  _GEN_6026 = ~cache_hit ? _GEN_3957 : _GEN_1718; // @[ICache.scala 175:32]
  wire  _GEN_6027 = ~cache_hit ? _GEN_3958 : _GEN_1207; // @[ICache.scala 175:32]
  wire  _GEN_6028 = ~cache_hit ? _GEN_3959 : _GEN_1719; // @[ICache.scala 175:32]
  wire  _GEN_6029 = ~cache_hit ? _GEN_3960 : _GEN_1208; // @[ICache.scala 175:32]
  wire  _GEN_6030 = ~cache_hit ? _GEN_3961 : _GEN_1720; // @[ICache.scala 175:32]
  wire  _GEN_6031 = ~cache_hit ? _GEN_3962 : _GEN_1209; // @[ICache.scala 175:32]
  wire  _GEN_6032 = ~cache_hit ? _GEN_3963 : _GEN_1721; // @[ICache.scala 175:32]
  wire  _GEN_6033 = ~cache_hit ? _GEN_3964 : _GEN_1210; // @[ICache.scala 175:32]
  wire  _GEN_6034 = ~cache_hit ? _GEN_3965 : _GEN_1722; // @[ICache.scala 175:32]
  wire  _GEN_6035 = ~cache_hit ? _GEN_3966 : _GEN_1211; // @[ICache.scala 175:32]
  wire  _GEN_6036 = ~cache_hit ? _GEN_3967 : _GEN_1723; // @[ICache.scala 175:32]
  wire  _GEN_6037 = ~cache_hit ? _GEN_3968 : _GEN_1212; // @[ICache.scala 175:32]
  wire  _GEN_6038 = ~cache_hit ? _GEN_3969 : _GEN_1724; // @[ICache.scala 175:32]
  wire  _GEN_6039 = ~cache_hit ? _GEN_3970 : _GEN_1213; // @[ICache.scala 175:32]
  wire  _GEN_6040 = ~cache_hit ? _GEN_3971 : _GEN_1725; // @[ICache.scala 175:32]
  wire  _GEN_6041 = ~cache_hit ? _GEN_3972 : _GEN_1214; // @[ICache.scala 175:32]
  wire  _GEN_6042 = ~cache_hit ? _GEN_3973 : _GEN_1726; // @[ICache.scala 175:32]
  wire  _GEN_6043 = ~cache_hit ? _GEN_3974 : _GEN_1215; // @[ICache.scala 175:32]
  wire  _GEN_6044 = ~cache_hit ? _GEN_3975 : _GEN_1727; // @[ICache.scala 175:32]
  wire  _GEN_6045 = ~cache_hit ? _GEN_3976 : _GEN_1216; // @[ICache.scala 175:32]
  wire  _GEN_6046 = ~cache_hit ? _GEN_3977 : _GEN_1728; // @[ICache.scala 175:32]
  wire  _GEN_6047 = ~cache_hit ? _GEN_3978 : _GEN_1217; // @[ICache.scala 175:32]
  wire  _GEN_6048 = ~cache_hit ? _GEN_3979 : _GEN_1729; // @[ICache.scala 175:32]
  wire  _GEN_6049 = ~cache_hit ? _GEN_3980 : _GEN_1218; // @[ICache.scala 175:32]
  wire  _GEN_6050 = ~cache_hit ? _GEN_3981 : _GEN_1730; // @[ICache.scala 175:32]
  wire  _GEN_6051 = ~cache_hit ? _GEN_3982 : _GEN_1219; // @[ICache.scala 175:32]
  wire  _GEN_6052 = ~cache_hit ? _GEN_3983 : _GEN_1731; // @[ICache.scala 175:32]
  wire  _GEN_6053 = ~cache_hit ? _GEN_3984 : _GEN_1220; // @[ICache.scala 175:32]
  wire  _GEN_6054 = ~cache_hit ? _GEN_3985 : _GEN_1732; // @[ICache.scala 175:32]
  wire  _GEN_6055 = ~cache_hit ? _GEN_3986 : _GEN_1221; // @[ICache.scala 175:32]
  wire  _GEN_6056 = ~cache_hit ? _GEN_3987 : _GEN_1733; // @[ICache.scala 175:32]
  wire  _GEN_6057 = ~cache_hit ? _GEN_3988 : _GEN_1222; // @[ICache.scala 175:32]
  wire  _GEN_6058 = ~cache_hit ? _GEN_3989 : _GEN_1734; // @[ICache.scala 175:32]
  wire  _GEN_6059 = ~cache_hit ? _GEN_3990 : _GEN_1223; // @[ICache.scala 175:32]
  wire  _GEN_6060 = ~cache_hit ? _GEN_3991 : _GEN_1735; // @[ICache.scala 175:32]
  wire  _GEN_6061 = ~cache_hit ? _GEN_3992 : _GEN_1224; // @[ICache.scala 175:32]
  wire  _GEN_6062 = ~cache_hit ? _GEN_3993 : _GEN_1736; // @[ICache.scala 175:32]
  wire  _GEN_6063 = ~cache_hit ? _GEN_3994 : _GEN_1225; // @[ICache.scala 175:32]
  wire  _GEN_6064 = ~cache_hit ? _GEN_3995 : _GEN_1737; // @[ICache.scala 175:32]
  wire  _GEN_6065 = ~cache_hit ? _GEN_3996 : _GEN_1226; // @[ICache.scala 175:32]
  wire  _GEN_6066 = ~cache_hit ? _GEN_3997 : _GEN_1738; // @[ICache.scala 175:32]
  wire  _GEN_6067 = ~cache_hit ? _GEN_3998 : _GEN_1227; // @[ICache.scala 175:32]
  wire  _GEN_6068 = ~cache_hit ? _GEN_3999 : _GEN_1739; // @[ICache.scala 175:32]
  wire  _GEN_6069 = ~cache_hit ? _GEN_4000 : _GEN_1228; // @[ICache.scala 175:32]
  wire  _GEN_6070 = ~cache_hit ? _GEN_4001 : _GEN_1740; // @[ICache.scala 175:32]
  wire  _GEN_6071 = ~cache_hit ? _GEN_4002 : _GEN_1229; // @[ICache.scala 175:32]
  wire  _GEN_6072 = ~cache_hit ? _GEN_4003 : _GEN_1741; // @[ICache.scala 175:32]
  wire  _GEN_6073 = ~cache_hit ? _GEN_4004 : _GEN_1230; // @[ICache.scala 175:32]
  wire  _GEN_6074 = ~cache_hit ? _GEN_4005 : _GEN_1742; // @[ICache.scala 175:32]
  wire  _GEN_6075 = ~cache_hit ? _GEN_4006 : _GEN_1231; // @[ICache.scala 175:32]
  wire  _GEN_6076 = ~cache_hit ? _GEN_4007 : _GEN_1743; // @[ICache.scala 175:32]
  wire  _GEN_6077 = ~cache_hit ? _GEN_4008 : _GEN_1232; // @[ICache.scala 175:32]
  wire  _GEN_6078 = ~cache_hit ? _GEN_4009 : _GEN_1744; // @[ICache.scala 175:32]
  wire  _GEN_6079 = ~cache_hit ? _GEN_4010 : _GEN_1233; // @[ICache.scala 175:32]
  wire  _GEN_6080 = ~cache_hit ? _GEN_4011 : _GEN_1745; // @[ICache.scala 175:32]
  wire  _GEN_6081 = ~cache_hit ? _GEN_4012 : _GEN_1234; // @[ICache.scala 175:32]
  wire  _GEN_6082 = ~cache_hit ? _GEN_4013 : _GEN_1746; // @[ICache.scala 175:32]
  wire  _GEN_6083 = ~cache_hit ? _GEN_4014 : _GEN_1235; // @[ICache.scala 175:32]
  wire  _GEN_6084 = ~cache_hit ? _GEN_4015 : _GEN_1747; // @[ICache.scala 175:32]
  wire  _GEN_6085 = ~cache_hit ? _GEN_4016 : _GEN_1236; // @[ICache.scala 175:32]
  wire  _GEN_6086 = ~cache_hit ? _GEN_4017 : _GEN_1748; // @[ICache.scala 175:32]
  wire  _GEN_6087 = ~cache_hit ? _GEN_4018 : _GEN_1237; // @[ICache.scala 175:32]
  wire  _GEN_6088 = ~cache_hit ? _GEN_4019 : _GEN_1749; // @[ICache.scala 175:32]
  wire  _GEN_6089 = ~cache_hit ? _GEN_4020 : _GEN_1238; // @[ICache.scala 175:32]
  wire  _GEN_6090 = ~cache_hit ? _GEN_4021 : _GEN_1750; // @[ICache.scala 175:32]
  wire  _GEN_6091 = ~cache_hit ? _GEN_4022 : _GEN_1239; // @[ICache.scala 175:32]
  wire  _GEN_6092 = ~cache_hit ? _GEN_4023 : _GEN_1751; // @[ICache.scala 175:32]
  wire  _GEN_6093 = ~cache_hit ? _GEN_4024 : _GEN_1240; // @[ICache.scala 175:32]
  wire  _GEN_6094 = ~cache_hit ? _GEN_4025 : _GEN_1752; // @[ICache.scala 175:32]
  wire  _GEN_6095 = ~cache_hit ? _GEN_4026 : _GEN_1241; // @[ICache.scala 175:32]
  wire  _GEN_6096 = ~cache_hit ? _GEN_4027 : _GEN_1753; // @[ICache.scala 175:32]
  wire  _GEN_6097 = ~cache_hit ? _GEN_4028 : _GEN_1242; // @[ICache.scala 175:32]
  wire  _GEN_6098 = ~cache_hit ? _GEN_4029 : _GEN_1754; // @[ICache.scala 175:32]
  wire  _GEN_6099 = ~cache_hit ? _GEN_4030 : _GEN_1243; // @[ICache.scala 175:32]
  wire  _GEN_6100 = ~cache_hit ? _GEN_4031 : _GEN_1755; // @[ICache.scala 175:32]
  wire  _GEN_6101 = ~cache_hit ? _GEN_4032 : _GEN_1244; // @[ICache.scala 175:32]
  wire  _GEN_6102 = ~cache_hit ? _GEN_4033 : _GEN_1756; // @[ICache.scala 175:32]
  wire  _GEN_6103 = ~cache_hit ? _GEN_4034 : _GEN_1245; // @[ICache.scala 175:32]
  wire  _GEN_6104 = ~cache_hit ? _GEN_4035 : _GEN_1757; // @[ICache.scala 175:32]
  wire  _GEN_6105 = ~cache_hit ? _GEN_4036 : _GEN_1246; // @[ICache.scala 175:32]
  wire  _GEN_6106 = ~cache_hit ? _GEN_4037 : _GEN_1758; // @[ICache.scala 175:32]
  wire  _GEN_6107 = ~cache_hit ? _GEN_4038 : _GEN_1247; // @[ICache.scala 175:32]
  wire  _GEN_6108 = ~cache_hit ? _GEN_4039 : _GEN_1759; // @[ICache.scala 175:32]
  wire  _GEN_6109 = ~cache_hit ? _GEN_4040 : _GEN_1248; // @[ICache.scala 175:32]
  wire  _GEN_6110 = ~cache_hit ? _GEN_4041 : _GEN_1760; // @[ICache.scala 175:32]
  wire  _GEN_6111 = ~cache_hit ? _GEN_4042 : _GEN_1249; // @[ICache.scala 175:32]
  wire  _GEN_6112 = ~cache_hit ? _GEN_4043 : _GEN_1761; // @[ICache.scala 175:32]
  wire  _GEN_6113 = ~cache_hit ? _GEN_4044 : _GEN_1250; // @[ICache.scala 175:32]
  wire  _GEN_6114 = ~cache_hit ? _GEN_4045 : _GEN_1762; // @[ICache.scala 175:32]
  wire  _GEN_6115 = ~cache_hit ? _GEN_4046 : _GEN_1251; // @[ICache.scala 175:32]
  wire  _GEN_6116 = ~cache_hit ? _GEN_4047 : _GEN_1763; // @[ICache.scala 175:32]
  wire  _GEN_6117 = ~cache_hit ? _GEN_4048 : _GEN_1252; // @[ICache.scala 175:32]
  wire  _GEN_6118 = ~cache_hit ? _GEN_4049 : _GEN_1764; // @[ICache.scala 175:32]
  wire  _GEN_6119 = ~cache_hit ? _GEN_4050 : _GEN_1253; // @[ICache.scala 175:32]
  wire  _GEN_6120 = ~cache_hit ? _GEN_4051 : _GEN_1765; // @[ICache.scala 175:32]
  wire  _GEN_6121 = ~cache_hit ? _GEN_4052 : _GEN_1254; // @[ICache.scala 175:32]
  wire  _GEN_6122 = ~cache_hit ? _GEN_4053 : _GEN_1766; // @[ICache.scala 175:32]
  wire  _GEN_6123 = ~cache_hit ? _GEN_4054 : _GEN_1255; // @[ICache.scala 175:32]
  wire  _GEN_6124 = ~cache_hit ? _GEN_4055 : _GEN_1767; // @[ICache.scala 175:32]
  wire  _GEN_6125 = ~cache_hit ? _GEN_4056 : _GEN_1256; // @[ICache.scala 175:32]
  wire  _GEN_6126 = ~cache_hit ? _GEN_4057 : _GEN_1768; // @[ICache.scala 175:32]
  wire  _GEN_6127 = ~cache_hit ? _GEN_4058 : _GEN_1257; // @[ICache.scala 175:32]
  wire  _GEN_6128 = ~cache_hit ? _GEN_4059 : _GEN_1769; // @[ICache.scala 175:32]
  wire  _GEN_6129 = ~cache_hit ? _GEN_4060 : _GEN_1258; // @[ICache.scala 175:32]
  wire  _GEN_6130 = ~cache_hit ? _GEN_4061 : _GEN_1770; // @[ICache.scala 175:32]
  wire  _GEN_6131 = ~cache_hit ? _GEN_4062 : _GEN_1259; // @[ICache.scala 175:32]
  wire  _GEN_6132 = ~cache_hit ? _GEN_4063 : _GEN_1771; // @[ICache.scala 175:32]
  wire  _GEN_6133 = ~cache_hit ? _GEN_4064 : _GEN_1260; // @[ICache.scala 175:32]
  wire  _GEN_6134 = ~cache_hit ? _GEN_4065 : _GEN_1772; // @[ICache.scala 175:32]
  wire  _GEN_6135 = ~cache_hit ? _GEN_4066 : _GEN_1261; // @[ICache.scala 175:32]
  wire  _GEN_6136 = ~cache_hit ? _GEN_4067 : _GEN_1773; // @[ICache.scala 175:32]
  wire  _GEN_6137 = ~cache_hit ? _GEN_4068 : _GEN_1262; // @[ICache.scala 175:32]
  wire  _GEN_6138 = ~cache_hit ? _GEN_4069 : _GEN_1774; // @[ICache.scala 175:32]
  wire  _GEN_6139 = ~cache_hit ? _GEN_4070 : _GEN_1263; // @[ICache.scala 175:32]
  wire  _GEN_6140 = ~cache_hit ? _GEN_4071 : _GEN_1775; // @[ICache.scala 175:32]
  wire  _GEN_6141 = ~cache_hit ? _GEN_4072 : _GEN_1264; // @[ICache.scala 175:32]
  wire  _GEN_6142 = ~cache_hit ? _GEN_4073 : _GEN_1776; // @[ICache.scala 175:32]
  wire  _GEN_6143 = ~cache_hit ? _GEN_4074 : _GEN_1265; // @[ICache.scala 175:32]
  wire  _GEN_6144 = ~cache_hit ? _GEN_4075 : _GEN_1777; // @[ICache.scala 175:32]
  wire  _GEN_6145 = ~cache_hit ? _GEN_4076 : _GEN_1266; // @[ICache.scala 175:32]
  wire  _GEN_6146 = ~cache_hit ? _GEN_4077 : _GEN_1778; // @[ICache.scala 175:32]
  wire  _GEN_6147 = ~cache_hit ? _GEN_4078 : _GEN_1267; // @[ICache.scala 175:32]
  wire  _GEN_6148 = ~cache_hit ? _GEN_4079 : _GEN_1779; // @[ICache.scala 175:32]
  wire  _GEN_6149 = ~cache_hit ? _GEN_4080 : _GEN_1268; // @[ICache.scala 175:32]
  wire  _GEN_6150 = ~cache_hit ? _GEN_4081 : _GEN_1780; // @[ICache.scala 175:32]
  wire  _GEN_6151 = ~cache_hit ? _GEN_4082 : _GEN_1269; // @[ICache.scala 175:32]
  wire  _GEN_6152 = ~cache_hit ? _GEN_4083 : _GEN_1781; // @[ICache.scala 175:32]
  wire  _GEN_6153 = ~cache_hit ? _GEN_4084 : _GEN_1270; // @[ICache.scala 175:32]
  wire  _GEN_6154 = ~cache_hit ? _GEN_4085 : _GEN_1782; // @[ICache.scala 175:32]
  wire  _GEN_6155 = ~cache_hit ? _GEN_4086 : _GEN_1271; // @[ICache.scala 175:32]
  wire  _GEN_6156 = ~cache_hit ? _GEN_4087 : _GEN_1783; // @[ICache.scala 175:32]
  wire  _GEN_6157 = ~cache_hit ? _GEN_4088 : _GEN_1272; // @[ICache.scala 175:32]
  wire  _GEN_6158 = ~cache_hit ? _GEN_4089 : _GEN_1784; // @[ICache.scala 175:32]
  wire  _GEN_6159 = ~cache_hit ? _GEN_4090 : _GEN_1273; // @[ICache.scala 175:32]
  wire  _GEN_6160 = ~cache_hit ? _GEN_4091 : _GEN_1785; // @[ICache.scala 175:32]
  wire  _GEN_6161 = ~cache_hit ? _GEN_4092 : _GEN_1274; // @[ICache.scala 175:32]
  wire  _GEN_6162 = ~cache_hit ? _GEN_4093 : _GEN_1786; // @[ICache.scala 175:32]
  wire  _GEN_6163 = ~cache_hit ? _GEN_4094 : _GEN_1275; // @[ICache.scala 175:32]
  wire  _GEN_6164 = ~cache_hit ? _GEN_4095 : _GEN_1787; // @[ICache.scala 175:32]
  wire  _GEN_6165 = ~cache_hit ? _GEN_4096 : _GEN_1276; // @[ICache.scala 175:32]
  wire  _GEN_6166 = ~cache_hit ? _GEN_4097 : _GEN_1788; // @[ICache.scala 175:32]
  wire  _GEN_6167 = ~cache_hit ? _GEN_4098 : _GEN_1277; // @[ICache.scala 175:32]
  wire  _GEN_6168 = ~cache_hit ? _GEN_4099 : _GEN_1789; // @[ICache.scala 175:32]
  wire  _GEN_6169 = ~cache_hit ? _GEN_4100 : _GEN_1278; // @[ICache.scala 175:32]
  wire  _GEN_6170 = ~cache_hit ? _GEN_4101 : _GEN_1790; // @[ICache.scala 175:32]
  wire  _GEN_6171 = ~cache_hit ? _GEN_4102 : _GEN_1279; // @[ICache.scala 175:32]
  wire  _GEN_6172 = ~cache_hit ? _GEN_4103 : _GEN_1791; // @[ICache.scala 175:32]
  wire  _GEN_6173 = ~cache_hit ? _GEN_4104 : _GEN_1280; // @[ICache.scala 175:32]
  wire  _GEN_6174 = ~cache_hit ? _GEN_4105 : _GEN_1792; // @[ICache.scala 175:32]
  wire  _GEN_6175 = ~cache_hit ? _GEN_4106 : _GEN_1281; // @[ICache.scala 175:32]
  wire  _GEN_6176 = ~cache_hit ? _GEN_4107 : _GEN_1793; // @[ICache.scala 175:32]
  wire  _GEN_6177 = ~cache_hit ? _GEN_4108 : _GEN_1282; // @[ICache.scala 175:32]
  wire  _GEN_6178 = ~cache_hit ? _GEN_4109 : _GEN_1794; // @[ICache.scala 175:32]
  wire  _GEN_6179 = ~cache_hit ? _GEN_4110 : _GEN_1283; // @[ICache.scala 175:32]
  wire  _GEN_6180 = ~cache_hit ? _GEN_4111 : _GEN_1795; // @[ICache.scala 175:32]
  wire  _GEN_6181 = ~cache_hit ? _GEN_4112 : _GEN_1284; // @[ICache.scala 175:32]
  wire  _GEN_6182 = ~cache_hit ? _GEN_4113 : _GEN_1796; // @[ICache.scala 175:32]
  wire  _GEN_6183 = ~cache_hit ? _GEN_4114 : _GEN_1285; // @[ICache.scala 175:32]
  wire  _GEN_6184 = ~cache_hit ? _GEN_4115 : _GEN_1797; // @[ICache.scala 175:32]
  wire  _GEN_6185 = ~cache_hit ? _GEN_4116 : _GEN_1286; // @[ICache.scala 175:32]
  wire  _GEN_6186 = ~cache_hit ? _GEN_4117 : _GEN_1798; // @[ICache.scala 175:32]
  wire  _GEN_6187 = ~cache_hit ? _GEN_4118 : _GEN_1287; // @[ICache.scala 175:32]
  wire  _GEN_6188 = ~cache_hit ? _GEN_4119 : _GEN_1799; // @[ICache.scala 175:32]
  wire  _GEN_6189 = ~cache_hit ? _GEN_4120 : _GEN_1288; // @[ICache.scala 175:32]
  wire  _GEN_6190 = ~cache_hit ? _GEN_4121 : _GEN_1800; // @[ICache.scala 175:32]
  wire  _GEN_6191 = ~cache_hit ? _GEN_4122 : _GEN_1289; // @[ICache.scala 175:32]
  wire  _GEN_6192 = ~cache_hit ? _GEN_4123 : _GEN_1801; // @[ICache.scala 175:32]
  wire  _GEN_6193 = ~cache_hit ? _GEN_4124 : _GEN_1290; // @[ICache.scala 175:32]
  wire  _GEN_6194 = ~cache_hit ? _GEN_4125 : _GEN_1802; // @[ICache.scala 175:32]
  wire  _GEN_6195 = ~cache_hit ? _GEN_4126 : _GEN_1291; // @[ICache.scala 175:32]
  wire  _GEN_6196 = ~cache_hit ? _GEN_4127 : _GEN_1803; // @[ICache.scala 175:32]
  wire  _GEN_6197 = ~cache_hit ? _GEN_4128 : _GEN_1292; // @[ICache.scala 175:32]
  wire  _GEN_6198 = ~cache_hit ? _GEN_4129 : _GEN_1804; // @[ICache.scala 175:32]
  wire  _GEN_6199 = ~cache_hit ? _GEN_4130 : _GEN_1293; // @[ICache.scala 175:32]
  wire  _GEN_6200 = ~cache_hit ? _GEN_4131 : _GEN_1805; // @[ICache.scala 175:32]
  wire  _GEN_6201 = ~cache_hit ? _GEN_4132 : _GEN_1294; // @[ICache.scala 175:32]
  wire  _GEN_6202 = ~cache_hit ? _GEN_4133 : _GEN_1806; // @[ICache.scala 175:32]
  wire  _GEN_6203 = ~cache_hit ? _GEN_4134 : _GEN_1295; // @[ICache.scala 175:32]
  wire  _GEN_6204 = ~cache_hit ? _GEN_4135 : _GEN_1807; // @[ICache.scala 175:32]
  wire  _GEN_6205 = ~cache_hit ? _GEN_4136 : _GEN_1296; // @[ICache.scala 175:32]
  wire  _GEN_6206 = ~cache_hit ? _GEN_4137 : _GEN_1808; // @[ICache.scala 175:32]
  wire  _GEN_6207 = ~cache_hit ? _GEN_4138 : _GEN_1297; // @[ICache.scala 175:32]
  wire  _GEN_6208 = ~cache_hit ? _GEN_4139 : _GEN_1809; // @[ICache.scala 175:32]
  wire  _GEN_6209 = ~cache_hit ? _GEN_4140 : _GEN_1298; // @[ICache.scala 175:32]
  wire  _GEN_6210 = ~cache_hit ? _GEN_4141 : _GEN_1810; // @[ICache.scala 175:32]
  wire  _GEN_6211 = ~cache_hit ? _GEN_4142 : _GEN_1299; // @[ICache.scala 175:32]
  wire  _GEN_6212 = ~cache_hit ? _GEN_4143 : _GEN_1811; // @[ICache.scala 175:32]
  wire  _GEN_6213 = ~cache_hit ? _GEN_4144 : _GEN_1300; // @[ICache.scala 175:32]
  wire  _GEN_6214 = ~cache_hit ? _GEN_4145 : _GEN_1812; // @[ICache.scala 175:32]
  wire  _GEN_6215 = ~cache_hit ? _GEN_4146 : _GEN_1301; // @[ICache.scala 175:32]
  wire  _GEN_6216 = ~cache_hit ? _GEN_4147 : _GEN_1813; // @[ICache.scala 175:32]
  wire  _GEN_6217 = ~cache_hit ? _GEN_4148 : _GEN_1302; // @[ICache.scala 175:32]
  wire  _GEN_6218 = ~cache_hit ? _GEN_4149 : _GEN_1814; // @[ICache.scala 175:32]
  wire  _GEN_6219 = ~cache_hit ? _GEN_4150 : _GEN_1303; // @[ICache.scala 175:32]
  wire  _GEN_6220 = ~cache_hit ? _GEN_4151 : _GEN_1815; // @[ICache.scala 175:32]
  wire  _GEN_6221 = ~cache_hit ? _GEN_4152 : _GEN_1304; // @[ICache.scala 175:32]
  wire  _GEN_6222 = ~cache_hit ? _GEN_4153 : _GEN_1816; // @[ICache.scala 175:32]
  wire  _GEN_6223 = ~cache_hit ? _GEN_4154 : _GEN_1305; // @[ICache.scala 175:32]
  wire  _GEN_6224 = ~cache_hit ? _GEN_4155 : _GEN_1817; // @[ICache.scala 175:32]
  wire  _GEN_6225 = ~cache_hit ? _GEN_4156 : _GEN_1306; // @[ICache.scala 175:32]
  wire  _GEN_6226 = ~cache_hit ? _GEN_4157 : _GEN_1818; // @[ICache.scala 175:32]
  wire  _GEN_6227 = ~cache_hit ? _GEN_4158 : _GEN_1307; // @[ICache.scala 175:32]
  wire  _GEN_6228 = ~cache_hit ? _GEN_4159 : _GEN_1819; // @[ICache.scala 175:32]
  wire  _GEN_6229 = ~cache_hit ? _GEN_4160 : _GEN_1308; // @[ICache.scala 175:32]
  wire  _GEN_6230 = ~cache_hit ? _GEN_4161 : _GEN_1820; // @[ICache.scala 175:32]
  wire  _GEN_6231 = ~cache_hit ? _GEN_4162 : _GEN_1309; // @[ICache.scala 175:32]
  wire  _GEN_6232 = ~cache_hit ? _GEN_4163 : _GEN_1821; // @[ICache.scala 175:32]
  wire  _GEN_6233 = ~cache_hit ? _GEN_4164 : _GEN_1310; // @[ICache.scala 175:32]
  wire  _GEN_6234 = ~cache_hit ? _GEN_4165 : _GEN_1822; // @[ICache.scala 175:32]
  wire  _GEN_6235 = ~cache_hit ? _GEN_4166 : _GEN_1311; // @[ICache.scala 175:32]
  wire  _GEN_6236 = ~cache_hit ? _GEN_4167 : _GEN_1823; // @[ICache.scala 175:32]
  wire  _GEN_6237 = ~cache_hit ? _GEN_4168 : _GEN_1312; // @[ICache.scala 175:32]
  wire  _GEN_6238 = ~cache_hit ? _GEN_4169 : _GEN_1824; // @[ICache.scala 175:32]
  wire  _GEN_6239 = ~cache_hit ? _GEN_4170 : _GEN_1313; // @[ICache.scala 175:32]
  wire  _GEN_6240 = ~cache_hit ? _GEN_4171 : _GEN_1825; // @[ICache.scala 175:32]
  wire  _GEN_6241 = ~cache_hit ? _GEN_4172 : _GEN_1314; // @[ICache.scala 175:32]
  wire  _GEN_6242 = ~cache_hit ? _GEN_4173 : _GEN_1826; // @[ICache.scala 175:32]
  wire  _GEN_6243 = ~cache_hit ? _GEN_4174 : _GEN_1315; // @[ICache.scala 175:32]
  wire  _GEN_6244 = ~cache_hit ? _GEN_4175 : _GEN_1827; // @[ICache.scala 175:32]
  wire  _GEN_6245 = ~cache_hit ? _GEN_4176 : _GEN_1316; // @[ICache.scala 175:32]
  wire  _GEN_6246 = ~cache_hit ? _GEN_4177 : _GEN_1828; // @[ICache.scala 175:32]
  wire  _GEN_6247 = ~cache_hit ? _GEN_4178 : _GEN_1317; // @[ICache.scala 175:32]
  wire  _GEN_6248 = ~cache_hit ? _GEN_4179 : _GEN_1829; // @[ICache.scala 175:32]
  wire  _GEN_6249 = ~cache_hit ? _GEN_4180 : _GEN_1318; // @[ICache.scala 175:32]
  wire  _GEN_6250 = ~cache_hit ? _GEN_4181 : _GEN_1830; // @[ICache.scala 175:32]
  wire  _GEN_6251 = ~cache_hit ? _GEN_4182 : _GEN_1319; // @[ICache.scala 175:32]
  wire  _GEN_6252 = ~cache_hit ? _GEN_4183 : _GEN_1831; // @[ICache.scala 175:32]
  wire  _GEN_6253 = ~cache_hit ? _GEN_4184 : _GEN_1320; // @[ICache.scala 175:32]
  wire  _GEN_6254 = ~cache_hit ? _GEN_4185 : _GEN_1832; // @[ICache.scala 175:32]
  wire  _GEN_6255 = ~cache_hit ? _GEN_4186 : _GEN_1321; // @[ICache.scala 175:32]
  wire  _GEN_6256 = ~cache_hit ? _GEN_4187 : _GEN_1833; // @[ICache.scala 175:32]
  wire  _GEN_6257 = ~cache_hit ? _GEN_4188 : _GEN_1322; // @[ICache.scala 175:32]
  wire  _GEN_6258 = ~cache_hit ? _GEN_4189 : _GEN_1834; // @[ICache.scala 175:32]
  wire  _GEN_6259 = ~cache_hit ? _GEN_4190 : _GEN_1323; // @[ICache.scala 175:32]
  wire  _GEN_6260 = ~cache_hit ? _GEN_4191 : _GEN_1835; // @[ICache.scala 175:32]
  wire  _GEN_6261 = ~cache_hit ? _GEN_4192 : _GEN_1324; // @[ICache.scala 175:32]
  wire  _GEN_6262 = ~cache_hit ? _GEN_4193 : _GEN_1836; // @[ICache.scala 175:32]
  wire  _GEN_6263 = ~cache_hit ? _GEN_4194 : _GEN_1325; // @[ICache.scala 175:32]
  wire  _GEN_6264 = ~cache_hit ? _GEN_4195 : _GEN_1837; // @[ICache.scala 175:32]
  wire  _GEN_6265 = ~cache_hit ? _GEN_4196 : _GEN_1326; // @[ICache.scala 175:32]
  wire  _GEN_6266 = ~cache_hit ? _GEN_4197 : _GEN_1838; // @[ICache.scala 175:32]
  wire  _GEN_6267 = ~cache_hit ? _GEN_4198 : _GEN_1327; // @[ICache.scala 175:32]
  wire  _GEN_6268 = ~cache_hit ? _GEN_4199 : _GEN_1839; // @[ICache.scala 175:32]
  wire  _GEN_6269 = ~cache_hit ? _GEN_4200 : _GEN_1328; // @[ICache.scala 175:32]
  wire  _GEN_6270 = ~cache_hit ? _GEN_4201 : _GEN_1840; // @[ICache.scala 175:32]
  wire  _GEN_6271 = ~cache_hit ? _GEN_4202 : _GEN_1329; // @[ICache.scala 175:32]
  wire  _GEN_6272 = ~cache_hit ? _GEN_4203 : _GEN_1841; // @[ICache.scala 175:32]
  wire  _GEN_6273 = ~cache_hit ? _GEN_4204 : _GEN_1330; // @[ICache.scala 175:32]
  wire  _GEN_6274 = ~cache_hit ? _GEN_4205 : _GEN_1842; // @[ICache.scala 175:32]
  wire  _GEN_6275 = ~cache_hit ? _GEN_4206 : _GEN_1331; // @[ICache.scala 175:32]
  wire  _GEN_6276 = ~cache_hit ? _GEN_4207 : _GEN_1843; // @[ICache.scala 175:32]
  wire  _GEN_6277 = ~cache_hit ? _GEN_4208 : _GEN_1332; // @[ICache.scala 175:32]
  wire  _GEN_6278 = ~cache_hit ? _GEN_4209 : _GEN_1844; // @[ICache.scala 175:32]
  wire  _GEN_6279 = ~cache_hit ? _GEN_4210 : _GEN_1333; // @[ICache.scala 175:32]
  wire  _GEN_6280 = ~cache_hit ? _GEN_4211 : _GEN_1845; // @[ICache.scala 175:32]
  wire  _GEN_6281 = ~cache_hit ? _GEN_4212 : _GEN_1334; // @[ICache.scala 175:32]
  wire  _GEN_6282 = ~cache_hit ? _GEN_4213 : _GEN_1846; // @[ICache.scala 175:32]
  wire  _GEN_6283 = ~cache_hit ? _GEN_4214 : _GEN_1335; // @[ICache.scala 175:32]
  wire  _GEN_6284 = ~cache_hit ? _GEN_4215 : _GEN_1847; // @[ICache.scala 175:32]
  wire  _GEN_6285 = ~cache_hit ? _GEN_4216 : _GEN_1336; // @[ICache.scala 175:32]
  wire  _GEN_6286 = ~cache_hit ? _GEN_4217 : _GEN_1848; // @[ICache.scala 175:32]
  wire  _GEN_6287 = ~cache_hit ? _GEN_4218 : _GEN_1337; // @[ICache.scala 175:32]
  wire  _GEN_6288 = ~cache_hit ? _GEN_4219 : _GEN_1849; // @[ICache.scala 175:32]
  wire  _GEN_6289 = ~cache_hit ? _GEN_4220 : _GEN_1338; // @[ICache.scala 175:32]
  wire  _GEN_6290 = ~cache_hit ? _GEN_4221 : _GEN_1850; // @[ICache.scala 175:32]
  wire  _GEN_6291 = ~cache_hit ? _GEN_4222 : _GEN_1339; // @[ICache.scala 175:32]
  wire  _GEN_6292 = ~cache_hit ? _GEN_4223 : _GEN_1851; // @[ICache.scala 175:32]
  wire  _GEN_6293 = ~cache_hit ? _GEN_4224 : _GEN_1340; // @[ICache.scala 175:32]
  wire  _GEN_6294 = ~cache_hit ? _GEN_4225 : _GEN_1852; // @[ICache.scala 175:32]
  wire  _GEN_6295 = ~cache_hit ? _GEN_4226 : _GEN_1341; // @[ICache.scala 175:32]
  wire  _GEN_6296 = ~cache_hit ? _GEN_4227 : _GEN_1853; // @[ICache.scala 175:32]
  wire  _GEN_6297 = ~cache_hit ? _GEN_4228 : _GEN_1342; // @[ICache.scala 175:32]
  wire  _GEN_6298 = ~cache_hit ? _GEN_4229 : _GEN_1854; // @[ICache.scala 175:32]
  wire  _GEN_6299 = ~cache_hit ? _GEN_4230 : _GEN_1343; // @[ICache.scala 175:32]
  wire  _GEN_6300 = ~cache_hit ? _GEN_4231 : _GEN_1855; // @[ICache.scala 175:32]
  wire  _GEN_6301 = ~cache_hit ? _GEN_4232 : _GEN_1344; // @[ICache.scala 175:32]
  wire  _GEN_6302 = ~cache_hit ? _GEN_4233 : _GEN_1856; // @[ICache.scala 175:32]
  wire  _GEN_6303 = ~cache_hit ? _GEN_4234 : _GEN_1345; // @[ICache.scala 175:32]
  wire  _GEN_6304 = ~cache_hit ? _GEN_4235 : _GEN_1857; // @[ICache.scala 175:32]
  wire  _GEN_6305 = ~cache_hit ? _GEN_4236 : _GEN_1346; // @[ICache.scala 175:32]
  wire  _GEN_6306 = ~cache_hit ? _GEN_4237 : _GEN_1858; // @[ICache.scala 175:32]
  wire  _GEN_6307 = ~cache_hit ? _GEN_4238 : _GEN_1347; // @[ICache.scala 175:32]
  wire  _GEN_6308 = ~cache_hit ? _GEN_4239 : _GEN_1859; // @[ICache.scala 175:32]
  wire  _GEN_6309 = ~cache_hit ? _GEN_4240 : _GEN_1348; // @[ICache.scala 175:32]
  wire  _GEN_6310 = ~cache_hit ? _GEN_4241 : _GEN_1860; // @[ICache.scala 175:32]
  wire  _GEN_6311 = ~cache_hit ? _GEN_4242 : _GEN_1349; // @[ICache.scala 175:32]
  wire  _GEN_6312 = ~cache_hit ? _GEN_4243 : _GEN_1861; // @[ICache.scala 175:32]
  wire  _GEN_6313 = ~cache_hit ? _GEN_4244 : _GEN_1350; // @[ICache.scala 175:32]
  wire  _GEN_6314 = ~cache_hit ? _GEN_4245 : _GEN_1862; // @[ICache.scala 175:32]
  wire  _GEN_6315 = ~cache_hit ? _GEN_4246 : _GEN_1351; // @[ICache.scala 175:32]
  wire  _GEN_6316 = ~cache_hit ? _GEN_4247 : _GEN_1863; // @[ICache.scala 175:32]
  wire  _GEN_6317 = ~cache_hit ? _GEN_4248 : _GEN_1352; // @[ICache.scala 175:32]
  wire  _GEN_6318 = ~cache_hit ? _GEN_4249 : _GEN_1864; // @[ICache.scala 175:32]
  wire  _GEN_6319 = ~cache_hit ? _GEN_4250 : _GEN_1353; // @[ICache.scala 175:32]
  wire  _GEN_6320 = ~cache_hit ? _GEN_4251 : _GEN_1865; // @[ICache.scala 175:32]
  wire  _GEN_6321 = ~cache_hit ? _GEN_4252 : _GEN_1354; // @[ICache.scala 175:32]
  wire  _GEN_6322 = ~cache_hit ? _GEN_4253 : _GEN_1866; // @[ICache.scala 175:32]
  wire  _GEN_6323 = ~cache_hit ? _GEN_4254 : _GEN_1355; // @[ICache.scala 175:32]
  wire  _GEN_6324 = ~cache_hit ? _GEN_4255 : _GEN_1867; // @[ICache.scala 175:32]
  wire  _GEN_6325 = ~cache_hit ? _GEN_4256 : _GEN_1356; // @[ICache.scala 175:32]
  wire  _GEN_6326 = ~cache_hit ? _GEN_4257 : _GEN_1868; // @[ICache.scala 175:32]
  wire  _GEN_6327 = ~cache_hit ? _GEN_4258 : _GEN_1357; // @[ICache.scala 175:32]
  wire  _GEN_6328 = ~cache_hit ? _GEN_4259 : _GEN_1869; // @[ICache.scala 175:32]
  wire  _GEN_6329 = ~cache_hit ? _GEN_4260 : _GEN_1358; // @[ICache.scala 175:32]
  wire  _GEN_6330 = ~cache_hit ? _GEN_4261 : _GEN_1870; // @[ICache.scala 175:32]
  wire  _GEN_6331 = ~cache_hit ? _GEN_4262 : _GEN_1359; // @[ICache.scala 175:32]
  wire  _GEN_6332 = ~cache_hit ? _GEN_4263 : _GEN_1871; // @[ICache.scala 175:32]
  wire  _GEN_6333 = ~cache_hit ? _GEN_4264 : _GEN_1360; // @[ICache.scala 175:32]
  wire  _GEN_6334 = ~cache_hit ? _GEN_4265 : _GEN_1872; // @[ICache.scala 175:32]
  wire  _GEN_6335 = ~cache_hit ? _GEN_4266 : _GEN_1361; // @[ICache.scala 175:32]
  wire  _GEN_6336 = ~cache_hit ? _GEN_4267 : _GEN_1873; // @[ICache.scala 175:32]
  wire  _GEN_6337 = ~cache_hit ? _GEN_4268 : _GEN_1362; // @[ICache.scala 175:32]
  wire  _GEN_6338 = ~cache_hit ? _GEN_4269 : _GEN_1874; // @[ICache.scala 175:32]
  wire  _GEN_6339 = ~cache_hit ? _GEN_4270 : _GEN_1363; // @[ICache.scala 175:32]
  wire  _GEN_6340 = ~cache_hit ? _GEN_4271 : _GEN_1875; // @[ICache.scala 175:32]
  wire  _GEN_6341 = ~cache_hit ? _GEN_4272 : _GEN_1364; // @[ICache.scala 175:32]
  wire  _GEN_6342 = ~cache_hit ? _GEN_4273 : _GEN_1876; // @[ICache.scala 175:32]
  wire  _GEN_6343 = ~cache_hit ? _GEN_4274 : _GEN_1365; // @[ICache.scala 175:32]
  wire  _GEN_6344 = ~cache_hit ? _GEN_4275 : _GEN_1877; // @[ICache.scala 175:32]
  wire  _GEN_6345 = ~cache_hit ? _GEN_4276 : _GEN_1366; // @[ICache.scala 175:32]
  wire  _GEN_6346 = ~cache_hit ? _GEN_4277 : _GEN_1878; // @[ICache.scala 175:32]
  wire  _GEN_6347 = ~cache_hit ? _GEN_4278 : _GEN_1367; // @[ICache.scala 175:32]
  wire  _GEN_6348 = ~cache_hit ? _GEN_4279 : _GEN_1879; // @[ICache.scala 175:32]
  wire  _GEN_6349 = ~cache_hit ? _GEN_4280 : _GEN_1368; // @[ICache.scala 175:32]
  wire  _GEN_6350 = ~cache_hit ? _GEN_4281 : _GEN_1880; // @[ICache.scala 175:32]
  wire  _GEN_6351 = ~cache_hit ? _GEN_4282 : _GEN_1369; // @[ICache.scala 175:32]
  wire  _GEN_6352 = ~cache_hit ? _GEN_4283 : _GEN_1881; // @[ICache.scala 175:32]
  wire  _GEN_6353 = ~cache_hit ? _GEN_4284 : _GEN_1370; // @[ICache.scala 175:32]
  wire  _GEN_6354 = ~cache_hit ? _GEN_4285 : _GEN_1882; // @[ICache.scala 175:32]
  wire  _GEN_6355 = ~cache_hit ? _GEN_4286 : _GEN_1371; // @[ICache.scala 175:32]
  wire  _GEN_6356 = ~cache_hit ? _GEN_4287 : _GEN_1883; // @[ICache.scala 175:32]
  wire  _GEN_6357 = ~cache_hit ? _GEN_4288 : _GEN_1372; // @[ICache.scala 175:32]
  wire  _GEN_6358 = ~cache_hit ? _GEN_4289 : _GEN_1884; // @[ICache.scala 175:32]
  wire  _GEN_6359 = ~cache_hit ? _GEN_4290 : _GEN_1373; // @[ICache.scala 175:32]
  wire  _GEN_6360 = ~cache_hit ? _GEN_4291 : _GEN_1885; // @[ICache.scala 175:32]
  wire  _GEN_6361 = ~cache_hit ? _GEN_4292 : _GEN_1374; // @[ICache.scala 175:32]
  wire  _GEN_6362 = ~cache_hit ? _GEN_4293 : _GEN_1886; // @[ICache.scala 175:32]
  wire  _GEN_6363 = ~cache_hit ? _GEN_4294 : _GEN_1375; // @[ICache.scala 175:32]
  wire  _GEN_6364 = ~cache_hit ? _GEN_4295 : _GEN_1887; // @[ICache.scala 175:32]
  wire  _GEN_6365 = ~cache_hit ? _GEN_4296 : _GEN_1376; // @[ICache.scala 175:32]
  wire  _GEN_6366 = ~cache_hit ? _GEN_4297 : _GEN_1888; // @[ICache.scala 175:32]
  wire  _GEN_6367 = ~cache_hit ? _GEN_4298 : _GEN_1377; // @[ICache.scala 175:32]
  wire  _GEN_6368 = ~cache_hit ? _GEN_4299 : _GEN_1889; // @[ICache.scala 175:32]
  wire  _GEN_6369 = ~cache_hit ? _GEN_4300 : _GEN_1378; // @[ICache.scala 175:32]
  wire  _GEN_6370 = ~cache_hit ? _GEN_4301 : _GEN_1890; // @[ICache.scala 175:32]
  wire  _GEN_6371 = ~cache_hit ? _GEN_4302 : _GEN_1379; // @[ICache.scala 175:32]
  wire  _GEN_6372 = ~cache_hit ? _GEN_4303 : _GEN_1891; // @[ICache.scala 175:32]
  wire  _GEN_6373 = ~cache_hit ? _GEN_4304 : _GEN_1380; // @[ICache.scala 175:32]
  wire  _GEN_6374 = ~cache_hit ? _GEN_4305 : _GEN_1892; // @[ICache.scala 175:32]
  wire  _GEN_6375 = ~cache_hit ? _GEN_4306 : _GEN_1381; // @[ICache.scala 175:32]
  wire  _GEN_6376 = ~cache_hit ? _GEN_4307 : _GEN_1893; // @[ICache.scala 175:32]
  wire  _GEN_6377 = ~cache_hit ? _GEN_4308 : _GEN_1382; // @[ICache.scala 175:32]
  wire  _GEN_6378 = ~cache_hit ? _GEN_4309 : _GEN_1894; // @[ICache.scala 175:32]
  wire  _GEN_6379 = ~cache_hit ? _GEN_4310 : _GEN_1383; // @[ICache.scala 175:32]
  wire  _GEN_6380 = ~cache_hit ? _GEN_4311 : _GEN_1895; // @[ICache.scala 175:32]
  wire  _GEN_6381 = ~cache_hit ? _GEN_4312 : _GEN_1384; // @[ICache.scala 175:32]
  wire  _GEN_6382 = ~cache_hit ? _GEN_4313 : _GEN_1896; // @[ICache.scala 175:32]
  wire  _GEN_6383 = ~cache_hit ? _GEN_4314 : _GEN_1385; // @[ICache.scala 175:32]
  wire  _GEN_6384 = ~cache_hit ? _GEN_4315 : _GEN_1897; // @[ICache.scala 175:32]
  wire  _GEN_6385 = ~cache_hit ? _GEN_4316 : _GEN_1386; // @[ICache.scala 175:32]
  wire  _GEN_6386 = ~cache_hit ? _GEN_4317 : _GEN_1898; // @[ICache.scala 175:32]
  wire  _GEN_6387 = ~cache_hit ? _GEN_4318 : _GEN_1387; // @[ICache.scala 175:32]
  wire  _GEN_6388 = ~cache_hit ? _GEN_4319 : _GEN_1899; // @[ICache.scala 175:32]
  wire  _GEN_6389 = ~cache_hit ? _GEN_4320 : _GEN_1388; // @[ICache.scala 175:32]
  wire  _GEN_6390 = ~cache_hit ? _GEN_4321 : _GEN_1900; // @[ICache.scala 175:32]
  wire  _GEN_6391 = ~cache_hit ? _GEN_4322 : _GEN_1389; // @[ICache.scala 175:32]
  wire  _GEN_6392 = ~cache_hit ? _GEN_4323 : _GEN_1901; // @[ICache.scala 175:32]
  wire  _GEN_6393 = ~cache_hit ? _GEN_4324 : _GEN_1390; // @[ICache.scala 175:32]
  wire  _GEN_6394 = ~cache_hit ? _GEN_4325 : _GEN_1902; // @[ICache.scala 175:32]
  wire  _GEN_6395 = ~cache_hit ? _GEN_4326 : _GEN_1391; // @[ICache.scala 175:32]
  wire  _GEN_6396 = ~cache_hit ? _GEN_4327 : _GEN_1903; // @[ICache.scala 175:32]
  wire  _GEN_6397 = ~cache_hit ? _GEN_4328 : _GEN_1392; // @[ICache.scala 175:32]
  wire  _GEN_6398 = ~cache_hit ? _GEN_4329 : _GEN_1904; // @[ICache.scala 175:32]
  wire  _GEN_6399 = ~cache_hit ? _GEN_4330 : _GEN_1393; // @[ICache.scala 175:32]
  wire  _GEN_6400 = ~cache_hit ? _GEN_4331 : _GEN_1905; // @[ICache.scala 175:32]
  wire  _GEN_6401 = ~cache_hit ? _GEN_4332 : _GEN_1394; // @[ICache.scala 175:32]
  wire  _GEN_6402 = ~cache_hit ? _GEN_4333 : _GEN_1906; // @[ICache.scala 175:32]
  wire  _GEN_6403 = ~cache_hit ? _GEN_4334 : _GEN_1395; // @[ICache.scala 175:32]
  wire  _GEN_6404 = ~cache_hit ? _GEN_4335 : _GEN_1907; // @[ICache.scala 175:32]
  wire  _GEN_6405 = ~cache_hit ? _GEN_4336 : _GEN_1396; // @[ICache.scala 175:32]
  wire  _GEN_6406 = ~cache_hit ? _GEN_4337 : _GEN_1908; // @[ICache.scala 175:32]
  wire  _GEN_6407 = ~cache_hit ? _GEN_4338 : _GEN_1397; // @[ICache.scala 175:32]
  wire  _GEN_6408 = ~cache_hit ? _GEN_4339 : _GEN_1909; // @[ICache.scala 175:32]
  wire  _GEN_6409 = ~cache_hit ? _GEN_4340 : _GEN_1398; // @[ICache.scala 175:32]
  wire  _GEN_6410 = ~cache_hit ? _GEN_4341 : _GEN_1910; // @[ICache.scala 175:32]
  wire  _GEN_6411 = ~cache_hit ? _GEN_4342 : _GEN_1399; // @[ICache.scala 175:32]
  wire  _GEN_6412 = ~cache_hit ? _GEN_4343 : _GEN_1911; // @[ICache.scala 175:32]
  wire  _GEN_6413 = ~cache_hit ? _GEN_4344 : _GEN_1400; // @[ICache.scala 175:32]
  wire  _GEN_6414 = ~cache_hit ? _GEN_4345 : _GEN_1912; // @[ICache.scala 175:32]
  wire  _GEN_6415 = ~cache_hit ? _GEN_4346 : _GEN_1401; // @[ICache.scala 175:32]
  wire  _GEN_6416 = ~cache_hit ? _GEN_4347 : _GEN_1913; // @[ICache.scala 175:32]
  wire  _GEN_6417 = ~cache_hit ? _GEN_4348 : _GEN_1402; // @[ICache.scala 175:32]
  wire  _GEN_6418 = ~cache_hit ? _GEN_4349 : _GEN_1914; // @[ICache.scala 175:32]
  wire  _GEN_6419 = ~cache_hit ? _GEN_4350 : _GEN_1403; // @[ICache.scala 175:32]
  wire  _GEN_6420 = ~cache_hit ? _GEN_4351 : _GEN_1915; // @[ICache.scala 175:32]
  wire  _GEN_6421 = ~cache_hit ? _GEN_4352 : _GEN_1404; // @[ICache.scala 175:32]
  wire  _GEN_6422 = ~cache_hit ? _GEN_4353 : _GEN_1916; // @[ICache.scala 175:32]
  wire  _GEN_6423 = ~cache_hit ? _GEN_4354 : _GEN_1405; // @[ICache.scala 175:32]
  wire  _GEN_6424 = ~cache_hit ? _GEN_4355 : _GEN_1917; // @[ICache.scala 175:32]
  wire  _GEN_6425 = ~cache_hit ? _GEN_4356 : _GEN_1406; // @[ICache.scala 175:32]
  wire  _GEN_6426 = ~cache_hit ? _GEN_4357 : _GEN_1918; // @[ICache.scala 175:32]
  wire  _GEN_6427 = ~cache_hit ? _GEN_4358 : _GEN_1407; // @[ICache.scala 175:32]
  wire  _GEN_6428 = ~cache_hit ? _GEN_4359 : _GEN_1919; // @[ICache.scala 175:32]
  wire  _GEN_6429 = ~cache_hit ? _GEN_4360 : _GEN_1408; // @[ICache.scala 175:32]
  wire  _GEN_6430 = ~cache_hit ? _GEN_4361 : _GEN_1920; // @[ICache.scala 175:32]
  wire  _GEN_6431 = ~cache_hit ? _GEN_4362 : _GEN_1409; // @[ICache.scala 175:32]
  wire  _GEN_6432 = ~cache_hit ? _GEN_4363 : _GEN_1921; // @[ICache.scala 175:32]
  wire  _GEN_6433 = ~cache_hit ? _GEN_4364 : _GEN_1410; // @[ICache.scala 175:32]
  wire  _GEN_6434 = ~cache_hit ? _GEN_4365 : _GEN_1922; // @[ICache.scala 175:32]
  wire  _GEN_6435 = ~cache_hit ? _GEN_4366 : _GEN_1411; // @[ICache.scala 175:32]
  wire  _GEN_6436 = ~cache_hit ? _GEN_4367 : _GEN_1923; // @[ICache.scala 175:32]
  wire  _GEN_6437 = ~cache_hit ? _GEN_4368 : _GEN_1412; // @[ICache.scala 175:32]
  wire  _GEN_6438 = ~cache_hit ? _GEN_4369 : _GEN_1924; // @[ICache.scala 175:32]
  wire  _GEN_6439 = ~cache_hit ? _GEN_4370 : _GEN_1413; // @[ICache.scala 175:32]
  wire  _GEN_6440 = ~cache_hit ? _GEN_4371 : _GEN_1925; // @[ICache.scala 175:32]
  wire  _GEN_6441 = ~cache_hit ? _GEN_4372 : _GEN_1414; // @[ICache.scala 175:32]
  wire  _GEN_6442 = ~cache_hit ? _GEN_4373 : _GEN_1926; // @[ICache.scala 175:32]
  wire  _GEN_6443 = ~cache_hit ? _GEN_4374 : _GEN_1415; // @[ICache.scala 175:32]
  wire  _GEN_6444 = ~cache_hit ? _GEN_4375 : _GEN_1927; // @[ICache.scala 175:32]
  wire  _GEN_6445 = ~cache_hit ? _GEN_4376 : _GEN_1416; // @[ICache.scala 175:32]
  wire  _GEN_6446 = ~cache_hit ? _GEN_4377 : _GEN_1928; // @[ICache.scala 175:32]
  wire  _GEN_6447 = ~cache_hit ? _GEN_4378 : _GEN_1417; // @[ICache.scala 175:32]
  wire  _GEN_6448 = ~cache_hit ? _GEN_4379 : _GEN_1929; // @[ICache.scala 175:32]
  wire  _GEN_6449 = ~cache_hit ? _GEN_4380 : _GEN_1418; // @[ICache.scala 175:32]
  wire  _GEN_6450 = ~cache_hit ? _GEN_4381 : _GEN_1930; // @[ICache.scala 175:32]
  wire  _GEN_6451 = ~cache_hit ? _GEN_4382 : _GEN_1419; // @[ICache.scala 175:32]
  wire  _GEN_6452 = ~cache_hit ? _GEN_4383 : _GEN_1931; // @[ICache.scala 175:32]
  wire  _GEN_6453 = ~cache_hit ? _GEN_4384 : _GEN_1420; // @[ICache.scala 175:32]
  wire  _GEN_6454 = ~cache_hit ? _GEN_4385 : _GEN_1932; // @[ICache.scala 175:32]
  wire  _GEN_6455 = ~cache_hit ? _GEN_4386 : _GEN_1421; // @[ICache.scala 175:32]
  wire  _GEN_6456 = ~cache_hit ? _GEN_4387 : _GEN_1933; // @[ICache.scala 175:32]
  wire  _GEN_6457 = ~cache_hit ? _GEN_4388 : _GEN_1422; // @[ICache.scala 175:32]
  wire  _GEN_6458 = ~cache_hit ? _GEN_4389 : _GEN_1934; // @[ICache.scala 175:32]
  wire  _GEN_6459 = ~cache_hit ? _GEN_4390 : _GEN_1423; // @[ICache.scala 175:32]
  wire  _GEN_6460 = ~cache_hit ? _GEN_4391 : _GEN_1935; // @[ICache.scala 175:32]
  wire  _GEN_6461 = ~cache_hit ? _GEN_4392 : _GEN_1424; // @[ICache.scala 175:32]
  wire  _GEN_6462 = ~cache_hit ? _GEN_4393 : _GEN_1936; // @[ICache.scala 175:32]
  wire  _GEN_6463 = ~cache_hit ? _GEN_4394 : _GEN_1425; // @[ICache.scala 175:32]
  wire  _GEN_6464 = ~cache_hit ? _GEN_4395 : _GEN_1937; // @[ICache.scala 175:32]
  wire  _GEN_6465 = ~cache_hit ? _GEN_4396 : _GEN_1426; // @[ICache.scala 175:32]
  wire  _GEN_6466 = ~cache_hit ? _GEN_4397 : _GEN_1938; // @[ICache.scala 175:32]
  wire  _GEN_6467 = ~cache_hit ? _GEN_4398 : _GEN_1427; // @[ICache.scala 175:32]
  wire  _GEN_6468 = ~cache_hit ? _GEN_4399 : _GEN_1939; // @[ICache.scala 175:32]
  wire  _GEN_6469 = ~cache_hit ? _GEN_4400 : _GEN_1428; // @[ICache.scala 175:32]
  wire  _GEN_6470 = ~cache_hit ? _GEN_4401 : _GEN_1940; // @[ICache.scala 175:32]
  wire  _GEN_6471 = ~cache_hit ? _GEN_4402 : _GEN_1429; // @[ICache.scala 175:32]
  wire  _GEN_6472 = ~cache_hit ? _GEN_4403 : _GEN_1941; // @[ICache.scala 175:32]
  wire  _GEN_6473 = ~cache_hit ? _GEN_4404 : _GEN_1430; // @[ICache.scala 175:32]
  wire  _GEN_6474 = ~cache_hit ? _GEN_4405 : _GEN_1942; // @[ICache.scala 175:32]
  wire  _GEN_6475 = ~cache_hit ? _GEN_4406 : _GEN_1431; // @[ICache.scala 175:32]
  wire  _GEN_6476 = ~cache_hit ? _GEN_4407 : _GEN_1943; // @[ICache.scala 175:32]
  wire  _GEN_6477 = ~cache_hit ? _GEN_4408 : _GEN_1432; // @[ICache.scala 175:32]
  wire  _GEN_6478 = ~cache_hit ? _GEN_4409 : _GEN_1944; // @[ICache.scala 175:32]
  wire  _GEN_6479 = ~cache_hit ? _GEN_4410 : _GEN_1433; // @[ICache.scala 175:32]
  wire  _GEN_6480 = ~cache_hit ? _GEN_4411 : _GEN_1945; // @[ICache.scala 175:32]
  wire  _GEN_6481 = ~cache_hit ? _GEN_4412 : _GEN_1434; // @[ICache.scala 175:32]
  wire  _GEN_6482 = ~cache_hit ? _GEN_4413 : _GEN_1946; // @[ICache.scala 175:32]
  wire  _GEN_6483 = ~cache_hit ? _GEN_4414 : _GEN_1435; // @[ICache.scala 175:32]
  wire  _GEN_6484 = ~cache_hit ? _GEN_4415 : _GEN_1947; // @[ICache.scala 175:32]
  wire  _GEN_6485 = ~cache_hit ? _GEN_4416 : _GEN_1436; // @[ICache.scala 175:32]
  wire  _GEN_6486 = ~cache_hit ? _GEN_4417 : _GEN_1948; // @[ICache.scala 175:32]
  wire  _GEN_6487 = ~cache_hit ? _GEN_4418 : _GEN_1437; // @[ICache.scala 175:32]
  wire  _GEN_6488 = ~cache_hit ? _GEN_4419 : _GEN_1949; // @[ICache.scala 175:32]
  wire  _GEN_6489 = ~cache_hit ? _GEN_4420 : _GEN_1438; // @[ICache.scala 175:32]
  wire  _GEN_6490 = ~cache_hit ? _GEN_4421 : _GEN_1950; // @[ICache.scala 175:32]
  wire  _GEN_6491 = ~cache_hit ? _GEN_4422 : _GEN_1439; // @[ICache.scala 175:32]
  wire  _GEN_6492 = ~cache_hit ? _GEN_4423 : _GEN_1951; // @[ICache.scala 175:32]
  wire  _GEN_6493 = ~cache_hit ? _GEN_4424 : _GEN_1440; // @[ICache.scala 175:32]
  wire  _GEN_6494 = ~cache_hit ? _GEN_4425 : _GEN_1952; // @[ICache.scala 175:32]
  wire  _GEN_6495 = ~cache_hit ? _GEN_4426 : _GEN_1441; // @[ICache.scala 175:32]
  wire  _GEN_6496 = ~cache_hit ? _GEN_4427 : _GEN_1953; // @[ICache.scala 175:32]
  wire  _GEN_6497 = ~cache_hit ? _GEN_4428 : _GEN_1442; // @[ICache.scala 175:32]
  wire  _GEN_6498 = ~cache_hit ? _GEN_4429 : _GEN_1954; // @[ICache.scala 175:32]
  wire  _GEN_6499 = ~cache_hit ? _GEN_4430 : _GEN_1443; // @[ICache.scala 175:32]
  wire  _GEN_6500 = ~cache_hit ? _GEN_4431 : _GEN_1955; // @[ICache.scala 175:32]
  wire  _GEN_6501 = ~cache_hit ? _GEN_4432 : _GEN_1444; // @[ICache.scala 175:32]
  wire  _GEN_6502 = ~cache_hit ? _GEN_4433 : _GEN_1956; // @[ICache.scala 175:32]
  wire  _GEN_6503 = ~cache_hit ? _GEN_4434 : _GEN_1445; // @[ICache.scala 175:32]
  wire  _GEN_6504 = ~cache_hit ? _GEN_4435 : _GEN_1957; // @[ICache.scala 175:32]
  wire  _GEN_6505 = ~cache_hit ? _GEN_4436 : _GEN_1446; // @[ICache.scala 175:32]
  wire  _GEN_6506 = ~cache_hit ? _GEN_4437 : _GEN_1958; // @[ICache.scala 175:32]
  wire  _GEN_6507 = ~cache_hit ? _GEN_4438 : _GEN_1447; // @[ICache.scala 175:32]
  wire  _GEN_6508 = ~cache_hit ? _GEN_4439 : _GEN_1959; // @[ICache.scala 175:32]
  wire  _GEN_6509 = ~cache_hit ? _GEN_4440 : _GEN_1448; // @[ICache.scala 175:32]
  wire  _GEN_6510 = ~cache_hit ? _GEN_4441 : _GEN_1960; // @[ICache.scala 175:32]
  wire  _GEN_6511 = ~cache_hit ? _GEN_4442 : _GEN_1449; // @[ICache.scala 175:32]
  wire  _GEN_6512 = ~cache_hit ? _GEN_4443 : _GEN_1961; // @[ICache.scala 175:32]
  wire  _GEN_6513 = ~cache_hit ? _GEN_4444 : _GEN_1450; // @[ICache.scala 175:32]
  wire  _GEN_6514 = ~cache_hit ? _GEN_4445 : _GEN_1962; // @[ICache.scala 175:32]
  wire  _GEN_6515 = ~cache_hit ? _GEN_4446 : _GEN_1451; // @[ICache.scala 175:32]
  wire  _GEN_6516 = ~cache_hit ? _GEN_4447 : _GEN_1963; // @[ICache.scala 175:32]
  wire  _GEN_6517 = ~cache_hit ? _GEN_4448 : _GEN_1452; // @[ICache.scala 175:32]
  wire  _GEN_6518 = ~cache_hit ? _GEN_4449 : _GEN_1964; // @[ICache.scala 175:32]
  wire  _GEN_6519 = ~cache_hit ? _GEN_4450 : _GEN_1453; // @[ICache.scala 175:32]
  wire  _GEN_6520 = ~cache_hit ? _GEN_4451 : _GEN_1965; // @[ICache.scala 175:32]
  wire  _GEN_6521 = ~cache_hit ? _GEN_4452 : _GEN_1454; // @[ICache.scala 175:32]
  wire  _GEN_6522 = ~cache_hit ? _GEN_4453 : _GEN_1966; // @[ICache.scala 175:32]
  wire  _GEN_6523 = ~cache_hit ? _GEN_4454 : _GEN_1455; // @[ICache.scala 175:32]
  wire  _GEN_6524 = ~cache_hit ? _GEN_4455 : _GEN_1967; // @[ICache.scala 175:32]
  wire  _GEN_6525 = ~cache_hit ? _GEN_4456 : _GEN_1456; // @[ICache.scala 175:32]
  wire  _GEN_6526 = ~cache_hit ? _GEN_4457 : _GEN_1968; // @[ICache.scala 175:32]
  wire  _GEN_6527 = ~cache_hit ? _GEN_4458 : _GEN_1457; // @[ICache.scala 175:32]
  wire  _GEN_6528 = ~cache_hit ? _GEN_4459 : _GEN_1969; // @[ICache.scala 175:32]
  wire  _GEN_6529 = ~cache_hit ? _GEN_4460 : _GEN_1458; // @[ICache.scala 175:32]
  wire  _GEN_6530 = ~cache_hit ? _GEN_4461 : _GEN_1970; // @[ICache.scala 175:32]
  wire  _GEN_6531 = ~cache_hit ? _GEN_4462 : _GEN_1459; // @[ICache.scala 175:32]
  wire  _GEN_6532 = ~cache_hit ? _GEN_4463 : _GEN_1971; // @[ICache.scala 175:32]
  wire  _GEN_6533 = ~cache_hit ? _GEN_4464 : _GEN_1460; // @[ICache.scala 175:32]
  wire  _GEN_6534 = ~cache_hit ? _GEN_4465 : _GEN_1972; // @[ICache.scala 175:32]
  wire  _GEN_6535 = ~cache_hit ? _GEN_4466 : _GEN_1461; // @[ICache.scala 175:32]
  wire  _GEN_6536 = ~cache_hit ? _GEN_4467 : _GEN_1973; // @[ICache.scala 175:32]
  wire  _GEN_6537 = ~cache_hit ? _GEN_4468 : _GEN_1462; // @[ICache.scala 175:32]
  wire  _GEN_6538 = ~cache_hit ? _GEN_4469 : _GEN_1974; // @[ICache.scala 175:32]
  wire  _GEN_6539 = ~cache_hit ? _GEN_4470 : _GEN_1463; // @[ICache.scala 175:32]
  wire  _GEN_6540 = ~cache_hit ? _GEN_4471 : _GEN_1975; // @[ICache.scala 175:32]
  wire  _GEN_6541 = ~cache_hit ? _GEN_4472 : _GEN_1464; // @[ICache.scala 175:32]
  wire  _GEN_6542 = ~cache_hit ? _GEN_4473 : _GEN_1976; // @[ICache.scala 175:32]
  wire  _GEN_6543 = ~cache_hit ? _GEN_4474 : _GEN_1465; // @[ICache.scala 175:32]
  wire  _GEN_6544 = ~cache_hit ? _GEN_4475 : _GEN_1977; // @[ICache.scala 175:32]
  wire  _GEN_6545 = ~cache_hit ? _GEN_4476 : _GEN_1466; // @[ICache.scala 175:32]
  wire  _GEN_6546 = ~cache_hit ? _GEN_4477 : _GEN_1978; // @[ICache.scala 175:32]
  wire  _GEN_6547 = ~cache_hit ? _GEN_4478 : _GEN_1467; // @[ICache.scala 175:32]
  wire  _GEN_6548 = ~cache_hit ? _GEN_4479 : _GEN_1979; // @[ICache.scala 175:32]
  wire  _GEN_6549 = ~cache_hit ? _GEN_4480 : _GEN_1468; // @[ICache.scala 175:32]
  wire  _GEN_6550 = ~cache_hit ? _GEN_4481 : _GEN_1980; // @[ICache.scala 175:32]
  wire  _GEN_6551 = ~cache_hit ? _GEN_4482 : _GEN_1469; // @[ICache.scala 175:32]
  wire  _GEN_6552 = ~cache_hit ? _GEN_4483 : _GEN_1981; // @[ICache.scala 175:32]
  wire  _GEN_6553 = ~cache_hit ? _GEN_4484 : _GEN_1470; // @[ICache.scala 175:32]
  wire  _GEN_6554 = ~cache_hit ? _GEN_4485 : _GEN_1982; // @[ICache.scala 175:32]
  wire  _GEN_6555 = ~cache_hit ? _GEN_4486 : _GEN_1471; // @[ICache.scala 175:32]
  wire  _GEN_6556 = ~cache_hit ? _GEN_4487 : _GEN_1983; // @[ICache.scala 175:32]
  wire  _GEN_6557 = ~cache_hit ? _GEN_4488 : _GEN_1472; // @[ICache.scala 175:32]
  wire  _GEN_6558 = ~cache_hit ? _GEN_4489 : _GEN_1984; // @[ICache.scala 175:32]
  wire  _GEN_6559 = ~cache_hit ? _GEN_4490 : _GEN_1473; // @[ICache.scala 175:32]
  wire  _GEN_6560 = ~cache_hit ? _GEN_4491 : _GEN_1985; // @[ICache.scala 175:32]
  wire  _GEN_6561 = ~cache_hit ? _GEN_4492 : _GEN_1474; // @[ICache.scala 175:32]
  wire  _GEN_6562 = ~cache_hit ? _GEN_4493 : _GEN_1986; // @[ICache.scala 175:32]
  wire  _GEN_6563 = ~cache_hit ? _GEN_4494 : _GEN_1475; // @[ICache.scala 175:32]
  wire  _GEN_6564 = ~cache_hit ? _GEN_4495 : _GEN_1987; // @[ICache.scala 175:32]
  wire  _GEN_6565 = ~cache_hit ? _GEN_4496 : _GEN_1476; // @[ICache.scala 175:32]
  wire  _GEN_6566 = ~cache_hit ? _GEN_4497 : _GEN_1988; // @[ICache.scala 175:32]
  wire  _GEN_6567 = ~cache_hit ? _GEN_4498 : _GEN_1477; // @[ICache.scala 175:32]
  wire  _GEN_6568 = ~cache_hit ? _GEN_4499 : _GEN_1989; // @[ICache.scala 175:32]
  wire  _GEN_6569 = ~cache_hit ? _GEN_4500 : _GEN_1478; // @[ICache.scala 175:32]
  wire  _GEN_6570 = ~cache_hit ? _GEN_4501 : _GEN_1990; // @[ICache.scala 175:32]
  wire  _GEN_6571 = ~cache_hit ? _GEN_4502 : _GEN_1479; // @[ICache.scala 175:32]
  wire  _GEN_6572 = ~cache_hit ? _GEN_4503 : _GEN_1991; // @[ICache.scala 175:32]
  wire  _GEN_6573 = ~cache_hit ? _GEN_4504 : _GEN_1480; // @[ICache.scala 175:32]
  wire  _GEN_6574 = ~cache_hit ? _GEN_4505 : _GEN_1992; // @[ICache.scala 175:32]
  wire  _GEN_6575 = ~cache_hit ? _GEN_4506 : _GEN_1481; // @[ICache.scala 175:32]
  wire  _GEN_6576 = ~cache_hit ? _GEN_4507 : _GEN_1993; // @[ICache.scala 175:32]
  wire  _GEN_6577 = ~cache_hit ? _GEN_4508 : _GEN_1482; // @[ICache.scala 175:32]
  wire  _GEN_6578 = ~cache_hit ? _GEN_4509 : _GEN_1994; // @[ICache.scala 175:32]
  wire  _GEN_6579 = ~cache_hit ? _GEN_4510 : _GEN_1483; // @[ICache.scala 175:32]
  wire  _GEN_6580 = ~cache_hit ? _GEN_4511 : _GEN_1995; // @[ICache.scala 175:32]
  wire  _GEN_6581 = ~cache_hit ? _GEN_4512 : _GEN_1484; // @[ICache.scala 175:32]
  wire  _GEN_6582 = ~cache_hit ? _GEN_4513 : _GEN_1996; // @[ICache.scala 175:32]
  wire  _GEN_6583 = ~cache_hit ? _GEN_4514 : _GEN_1485; // @[ICache.scala 175:32]
  wire  _GEN_6584 = ~cache_hit ? _GEN_4515 : _GEN_1997; // @[ICache.scala 175:32]
  wire  _GEN_6585 = ~cache_hit ? _GEN_4516 : _GEN_1486; // @[ICache.scala 175:32]
  wire  _GEN_6586 = ~cache_hit ? _GEN_4517 : _GEN_1998; // @[ICache.scala 175:32]
  wire  _GEN_6587 = ~cache_hit ? _GEN_4518 : _GEN_1487; // @[ICache.scala 175:32]
  wire  _GEN_6588 = ~cache_hit ? _GEN_4519 : _GEN_1999; // @[ICache.scala 175:32]
  wire  _GEN_6589 = ~cache_hit ? _GEN_4520 : _GEN_1488; // @[ICache.scala 175:32]
  wire  _GEN_6590 = ~cache_hit ? _GEN_4521 : _GEN_2000; // @[ICache.scala 175:32]
  wire  _GEN_6591 = ~cache_hit ? _GEN_4522 : _GEN_1489; // @[ICache.scala 175:32]
  wire  _GEN_6592 = ~cache_hit ? _GEN_4523 : _GEN_2001; // @[ICache.scala 175:32]
  wire  _GEN_6593 = ~cache_hit ? _GEN_4524 : _GEN_1490; // @[ICache.scala 175:32]
  wire  _GEN_6594 = ~cache_hit ? _GEN_4525 : _GEN_2002; // @[ICache.scala 175:32]
  wire  _GEN_6595 = ~cache_hit ? _GEN_4526 : _GEN_1491; // @[ICache.scala 175:32]
  wire  _GEN_6596 = ~cache_hit ? _GEN_4527 : _GEN_2003; // @[ICache.scala 175:32]
  wire  _GEN_6597 = ~cache_hit ? _GEN_4528 : _GEN_1492; // @[ICache.scala 175:32]
  wire  _GEN_6598 = ~cache_hit ? _GEN_4529 : _GEN_2004; // @[ICache.scala 175:32]
  wire  _GEN_6599 = ~cache_hit ? _GEN_4530 : _GEN_1493; // @[ICache.scala 175:32]
  wire  _GEN_6600 = ~cache_hit ? _GEN_4531 : _GEN_2005; // @[ICache.scala 175:32]
  wire  _GEN_6601 = ~cache_hit ? _GEN_4532 : _GEN_1494; // @[ICache.scala 175:32]
  wire  _GEN_6602 = ~cache_hit ? _GEN_4533 : _GEN_2006; // @[ICache.scala 175:32]
  wire  _GEN_6603 = ~cache_hit ? _GEN_4534 : _GEN_1495; // @[ICache.scala 175:32]
  wire  _GEN_6604 = ~cache_hit ? _GEN_4535 : _GEN_2007; // @[ICache.scala 175:32]
  wire  _GEN_6605 = ~cache_hit ? _GEN_4536 : _GEN_1496; // @[ICache.scala 175:32]
  wire  _GEN_6606 = ~cache_hit ? _GEN_4537 : _GEN_2008; // @[ICache.scala 175:32]
  wire  _GEN_6607 = ~cache_hit ? _GEN_4538 : _GEN_1497; // @[ICache.scala 175:32]
  wire  _GEN_6608 = ~cache_hit ? _GEN_4539 : _GEN_2009; // @[ICache.scala 175:32]
  wire  _GEN_6609 = ~cache_hit ? _GEN_4540 : _GEN_1498; // @[ICache.scala 175:32]
  wire  _GEN_6610 = ~cache_hit ? _GEN_4541 : _GEN_2010; // @[ICache.scala 175:32]
  wire  _GEN_6611 = ~cache_hit ? _GEN_4542 : _GEN_1499; // @[ICache.scala 175:32]
  wire  _GEN_6612 = ~cache_hit ? _GEN_4543 : _GEN_2011; // @[ICache.scala 175:32]
  wire  _GEN_6613 = ~cache_hit ? _GEN_4544 : _GEN_1500; // @[ICache.scala 175:32]
  wire  _GEN_6614 = ~cache_hit ? _GEN_4545 : _GEN_2012; // @[ICache.scala 175:32]
  wire  _GEN_6615 = ~cache_hit ? _GEN_4546 : _GEN_1501; // @[ICache.scala 175:32]
  wire  _GEN_6616 = ~cache_hit ? _GEN_4547 : _GEN_2013; // @[ICache.scala 175:32]
  wire  _GEN_6617 = ~cache_hit ? _GEN_4548 : _GEN_1502; // @[ICache.scala 175:32]
  wire  _GEN_6618 = ~cache_hit ? _GEN_4549 : _GEN_2014; // @[ICache.scala 175:32]
  wire  _GEN_6619 = ~cache_hit ? _GEN_4550 : _GEN_1503; // @[ICache.scala 175:32]
  wire  _GEN_6620 = ~cache_hit ? _GEN_4551 : _GEN_2015; // @[ICache.scala 175:32]
  wire  _GEN_6621 = ~cache_hit ? _GEN_4552 : _GEN_1504; // @[ICache.scala 175:32]
  wire  _GEN_6622 = ~cache_hit ? _GEN_4553 : _GEN_2016; // @[ICache.scala 175:32]
  wire  _GEN_6623 = ~cache_hit ? _GEN_4554 : _GEN_1505; // @[ICache.scala 175:32]
  wire  _GEN_6624 = ~cache_hit ? _GEN_4555 : _GEN_2017; // @[ICache.scala 175:32]
  wire  _GEN_6625 = ~cache_hit ? _GEN_4556 : _GEN_1506; // @[ICache.scala 175:32]
  wire  _GEN_6626 = ~cache_hit ? _GEN_4557 : _GEN_2018; // @[ICache.scala 175:32]
  wire  _GEN_6627 = ~cache_hit ? _GEN_4558 : _GEN_1507; // @[ICache.scala 175:32]
  wire  _GEN_6628 = ~cache_hit ? _GEN_4559 : _GEN_2019; // @[ICache.scala 175:32]
  wire  _GEN_6629 = ~cache_hit ? _GEN_4560 : _GEN_1508; // @[ICache.scala 175:32]
  wire  _GEN_6630 = ~cache_hit ? _GEN_4561 : _GEN_2020; // @[ICache.scala 175:32]
  wire  _GEN_6631 = ~cache_hit ? _GEN_4562 : _GEN_1509; // @[ICache.scala 175:32]
  wire  _GEN_6632 = ~cache_hit ? _GEN_4563 : _GEN_2021; // @[ICache.scala 175:32]
  wire  _GEN_6633 = ~cache_hit ? _GEN_4564 : _GEN_1510; // @[ICache.scala 175:32]
  wire  _GEN_6634 = ~cache_hit ? _GEN_4565 : _GEN_2022; // @[ICache.scala 175:32]
  wire  _GEN_6635 = ~cache_hit ? _GEN_4566 : _GEN_1511; // @[ICache.scala 175:32]
  wire  _GEN_6636 = ~cache_hit ? _GEN_4567 : _GEN_2023; // @[ICache.scala 175:32]
  wire  _GEN_6637 = ~cache_hit ? _GEN_4568 : _GEN_1512; // @[ICache.scala 175:32]
  wire  _GEN_6638 = ~cache_hit ? _GEN_4569 : _GEN_2024; // @[ICache.scala 175:32]
  wire  _GEN_6639 = ~cache_hit ? _GEN_4570 : _GEN_1513; // @[ICache.scala 175:32]
  wire  _GEN_6640 = ~cache_hit ? _GEN_4571 : _GEN_2025; // @[ICache.scala 175:32]
  wire  _GEN_6641 = ~cache_hit ? _GEN_4572 : _GEN_1514; // @[ICache.scala 175:32]
  wire  _GEN_6642 = ~cache_hit ? _GEN_4573 : _GEN_2026; // @[ICache.scala 175:32]
  wire  _GEN_6643 = ~cache_hit ? _GEN_4574 : _GEN_1515; // @[ICache.scala 175:32]
  wire  _GEN_6644 = ~cache_hit ? _GEN_4575 : _GEN_2027; // @[ICache.scala 175:32]
  wire  _GEN_6645 = ~cache_hit ? _GEN_4576 : _GEN_1516; // @[ICache.scala 175:32]
  wire  _GEN_6646 = ~cache_hit ? _GEN_4577 : _GEN_2028; // @[ICache.scala 175:32]
  wire  _GEN_6647 = ~cache_hit ? _GEN_4578 : _GEN_1517; // @[ICache.scala 175:32]
  wire  _GEN_6648 = ~cache_hit ? _GEN_4579 : _GEN_2029; // @[ICache.scala 175:32]
  wire  _GEN_6649 = ~cache_hit ? _GEN_4580 : _GEN_1518; // @[ICache.scala 175:32]
  wire  _GEN_6650 = ~cache_hit ? _GEN_4581 : _GEN_2030; // @[ICache.scala 175:32]
  wire  _GEN_6651 = ~cache_hit ? _GEN_4582 : _GEN_1519; // @[ICache.scala 175:32]
  wire  _GEN_6652 = ~cache_hit ? _GEN_4583 : _GEN_2031; // @[ICache.scala 175:32]
  wire  _GEN_6653 = ~cache_hit ? _GEN_4584 : _GEN_1520; // @[ICache.scala 175:32]
  wire  _GEN_6654 = ~cache_hit ? _GEN_4585 : _GEN_2032; // @[ICache.scala 175:32]
  wire  _GEN_6655 = ~cache_hit ? _GEN_4586 : _GEN_1521; // @[ICache.scala 175:32]
  wire  _GEN_6656 = ~cache_hit ? _GEN_4587 : _GEN_2033; // @[ICache.scala 175:32]
  wire  _GEN_6657 = ~cache_hit ? _GEN_4588 : _GEN_1522; // @[ICache.scala 175:32]
  wire  _GEN_6658 = ~cache_hit ? _GEN_4589 : _GEN_2034; // @[ICache.scala 175:32]
  wire  _GEN_6659 = ~cache_hit ? _GEN_4590 : _GEN_1523; // @[ICache.scala 175:32]
  wire  _GEN_6660 = ~cache_hit ? _GEN_4591 : _GEN_2035; // @[ICache.scala 175:32]
  wire  _GEN_6661 = ~cache_hit ? _GEN_4592 : _GEN_1524; // @[ICache.scala 175:32]
  wire  _GEN_6662 = ~cache_hit ? _GEN_4593 : _GEN_2036; // @[ICache.scala 175:32]
  wire  _GEN_6663 = ~cache_hit ? _GEN_4594 : _GEN_1525; // @[ICache.scala 175:32]
  wire  _GEN_6664 = ~cache_hit ? _GEN_4595 : _GEN_2037; // @[ICache.scala 175:32]
  wire  _GEN_6665 = ~cache_hit ? _GEN_4596 : _GEN_1526; // @[ICache.scala 175:32]
  wire  _GEN_6666 = ~cache_hit ? _GEN_4597 : _GEN_2038; // @[ICache.scala 175:32]
  wire  _GEN_6667 = ~cache_hit ? _GEN_4598 : _GEN_1527; // @[ICache.scala 175:32]
  wire  _GEN_6668 = ~cache_hit ? _GEN_4599 : _GEN_2039; // @[ICache.scala 175:32]
  wire  _GEN_6669 = ~cache_hit ? _GEN_4600 : _GEN_1528; // @[ICache.scala 175:32]
  wire  _GEN_6670 = ~cache_hit ? _GEN_4601 : _GEN_2040; // @[ICache.scala 175:32]
  wire  _GEN_6671 = ~cache_hit ? _GEN_4602 : _GEN_1529; // @[ICache.scala 175:32]
  wire  _GEN_6672 = ~cache_hit ? _GEN_4603 : _GEN_2041; // @[ICache.scala 175:32]
  wire  _GEN_6673 = ~cache_hit ? _GEN_4604 : _GEN_1530; // @[ICache.scala 175:32]
  wire  _GEN_6674 = ~cache_hit ? _GEN_4605 : _GEN_2042; // @[ICache.scala 175:32]
  wire  _GEN_6675 = ~cache_hit ? _GEN_4606 : _GEN_1531; // @[ICache.scala 175:32]
  wire  _GEN_6676 = ~cache_hit ? _GEN_4607 : _GEN_2043; // @[ICache.scala 175:32]
  wire  _GEN_6677 = ~cache_hit ? _GEN_4608 : _GEN_1532; // @[ICache.scala 175:32]
  wire  _GEN_6678 = ~cache_hit ? _GEN_4609 : _GEN_2044; // @[ICache.scala 175:32]
  wire  _GEN_6679 = ~cache_hit ? _GEN_4610 : _GEN_1533; // @[ICache.scala 175:32]
  wire  _GEN_6680 = ~cache_hit ? _GEN_4611 : _GEN_2045; // @[ICache.scala 175:32]
  wire  _GEN_6681 = ~cache_hit ? _GEN_4612 : _GEN_1534; // @[ICache.scala 175:32]
  wire  _GEN_6682 = ~cache_hit ? _GEN_4613 : _GEN_2046; // @[ICache.scala 175:32]
  wire  _GEN_6683 = ~cache_hit ? _GEN_4614 : _GEN_1535; // @[ICache.scala 175:32]
  wire  _GEN_6684 = ~cache_hit ? _GEN_4615 : _GEN_2047; // @[ICache.scala 175:32]
  wire  _GEN_6685 = ~cache_hit ? _GEN_4616 : _GEN_1536; // @[ICache.scala 175:32]
  wire  _GEN_6686 = ~cache_hit ? _GEN_4617 : _GEN_2048; // @[ICache.scala 175:32]
  wire  _GEN_6687 = ~cache_hit ? _GEN_4618 : _GEN_1537; // @[ICache.scala 175:32]
  wire  _GEN_6688 = ~cache_hit ? _GEN_4619 : _GEN_2049; // @[ICache.scala 175:32]
  wire  _GEN_6689 = ~cache_hit ? _GEN_4620 : _GEN_1538; // @[ICache.scala 175:32]
  wire  _GEN_6690 = ~cache_hit ? _GEN_4621 : _GEN_2050; // @[ICache.scala 175:32]
  wire [4:0] _GEN_6691 = ~cache_hit ? 5'h0 : axi_cnt_value; // @[ICache.scala 175:32 Counter.scala 98:11 61:40]
  wire  _GEN_6692 = ~cache_hit ? lru_0 : _GEN_5138; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6693 = ~cache_hit ? lru_1 : _GEN_5139; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6694 = ~cache_hit ? lru_2 : _GEN_5140; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6695 = ~cache_hit ? lru_3 : _GEN_5141; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6696 = ~cache_hit ? lru_4 : _GEN_5142; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6697 = ~cache_hit ? lru_5 : _GEN_5143; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6698 = ~cache_hit ? lru_6 : _GEN_5144; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6699 = ~cache_hit ? lru_7 : _GEN_5145; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6700 = ~cache_hit ? lru_8 : _GEN_5146; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6701 = ~cache_hit ? lru_9 : _GEN_5147; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6702 = ~cache_hit ? lru_10 : _GEN_5148; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6703 = ~cache_hit ? lru_11 : _GEN_5149; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6704 = ~cache_hit ? lru_12 : _GEN_5150; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6705 = ~cache_hit ? lru_13 : _GEN_5151; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6706 = ~cache_hit ? lru_14 : _GEN_5152; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6707 = ~cache_hit ? lru_15 : _GEN_5153; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6708 = ~cache_hit ? lru_16 : _GEN_5154; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6709 = ~cache_hit ? lru_17 : _GEN_5155; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6710 = ~cache_hit ? lru_18 : _GEN_5156; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6711 = ~cache_hit ? lru_19 : _GEN_5157; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6712 = ~cache_hit ? lru_20 : _GEN_5158; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6713 = ~cache_hit ? lru_21 : _GEN_5159; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6714 = ~cache_hit ? lru_22 : _GEN_5160; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6715 = ~cache_hit ? lru_23 : _GEN_5161; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6716 = ~cache_hit ? lru_24 : _GEN_5162; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6717 = ~cache_hit ? lru_25 : _GEN_5163; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6718 = ~cache_hit ? lru_26 : _GEN_5164; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6719 = ~cache_hit ? lru_27 : _GEN_5165; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6720 = ~cache_hit ? lru_28 : _GEN_5166; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6721 = ~cache_hit ? lru_29 : _GEN_5167; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6722 = ~cache_hit ? lru_30 : _GEN_5168; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6723 = ~cache_hit ? lru_31 : _GEN_5169; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6724 = ~cache_hit ? lru_32 : _GEN_5170; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6725 = ~cache_hit ? lru_33 : _GEN_5171; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6726 = ~cache_hit ? lru_34 : _GEN_5172; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6727 = ~cache_hit ? lru_35 : _GEN_5173; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6728 = ~cache_hit ? lru_36 : _GEN_5174; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6729 = ~cache_hit ? lru_37 : _GEN_5175; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6730 = ~cache_hit ? lru_38 : _GEN_5176; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6731 = ~cache_hit ? lru_39 : _GEN_5177; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6732 = ~cache_hit ? lru_40 : _GEN_5178; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6733 = ~cache_hit ? lru_41 : _GEN_5179; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6734 = ~cache_hit ? lru_42 : _GEN_5180; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6735 = ~cache_hit ? lru_43 : _GEN_5181; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6736 = ~cache_hit ? lru_44 : _GEN_5182; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6737 = ~cache_hit ? lru_45 : _GEN_5183; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6738 = ~cache_hit ? lru_46 : _GEN_5184; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6739 = ~cache_hit ? lru_47 : _GEN_5185; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6740 = ~cache_hit ? lru_48 : _GEN_5186; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6741 = ~cache_hit ? lru_49 : _GEN_5187; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6742 = ~cache_hit ? lru_50 : _GEN_5188; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6743 = ~cache_hit ? lru_51 : _GEN_5189; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6744 = ~cache_hit ? lru_52 : _GEN_5190; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6745 = ~cache_hit ? lru_53 : _GEN_5191; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6746 = ~cache_hit ? lru_54 : _GEN_5192; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6747 = ~cache_hit ? lru_55 : _GEN_5193; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6748 = ~cache_hit ? lru_56 : _GEN_5194; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6749 = ~cache_hit ? lru_57 : _GEN_5195; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6750 = ~cache_hit ? lru_58 : _GEN_5196; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6751 = ~cache_hit ? lru_59 : _GEN_5197; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6752 = ~cache_hit ? lru_60 : _GEN_5198; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6753 = ~cache_hit ? lru_61 : _GEN_5199; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6754 = ~cache_hit ? lru_62 : _GEN_5200; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6755 = ~cache_hit ? lru_63 : _GEN_5201; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6756 = ~cache_hit ? lru_64 : _GEN_5202; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6757 = ~cache_hit ? lru_65 : _GEN_5203; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6758 = ~cache_hit ? lru_66 : _GEN_5204; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6759 = ~cache_hit ? lru_67 : _GEN_5205; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6760 = ~cache_hit ? lru_68 : _GEN_5206; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6761 = ~cache_hit ? lru_69 : _GEN_5207; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6762 = ~cache_hit ? lru_70 : _GEN_5208; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6763 = ~cache_hit ? lru_71 : _GEN_5209; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6764 = ~cache_hit ? lru_72 : _GEN_5210; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6765 = ~cache_hit ? lru_73 : _GEN_5211; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6766 = ~cache_hit ? lru_74 : _GEN_5212; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6767 = ~cache_hit ? lru_75 : _GEN_5213; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6768 = ~cache_hit ? lru_76 : _GEN_5214; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6769 = ~cache_hit ? lru_77 : _GEN_5215; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6770 = ~cache_hit ? lru_78 : _GEN_5216; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6771 = ~cache_hit ? lru_79 : _GEN_5217; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6772 = ~cache_hit ? lru_80 : _GEN_5218; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6773 = ~cache_hit ? lru_81 : _GEN_5219; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6774 = ~cache_hit ? lru_82 : _GEN_5220; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6775 = ~cache_hit ? lru_83 : _GEN_5221; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6776 = ~cache_hit ? lru_84 : _GEN_5222; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6777 = ~cache_hit ? lru_85 : _GEN_5223; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6778 = ~cache_hit ? lru_86 : _GEN_5224; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6779 = ~cache_hit ? lru_87 : _GEN_5225; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6780 = ~cache_hit ? lru_88 : _GEN_5226; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6781 = ~cache_hit ? lru_89 : _GEN_5227; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6782 = ~cache_hit ? lru_90 : _GEN_5228; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6783 = ~cache_hit ? lru_91 : _GEN_5229; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6784 = ~cache_hit ? lru_92 : _GEN_5230; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6785 = ~cache_hit ? lru_93 : _GEN_5231; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6786 = ~cache_hit ? lru_94 : _GEN_5232; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6787 = ~cache_hit ? lru_95 : _GEN_5233; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6788 = ~cache_hit ? lru_96 : _GEN_5234; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6789 = ~cache_hit ? lru_97 : _GEN_5235; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6790 = ~cache_hit ? lru_98 : _GEN_5236; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6791 = ~cache_hit ? lru_99 : _GEN_5237; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6792 = ~cache_hit ? lru_100 : _GEN_5238; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6793 = ~cache_hit ? lru_101 : _GEN_5239; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6794 = ~cache_hit ? lru_102 : _GEN_5240; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6795 = ~cache_hit ? lru_103 : _GEN_5241; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6796 = ~cache_hit ? lru_104 : _GEN_5242; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6797 = ~cache_hit ? lru_105 : _GEN_5243; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6798 = ~cache_hit ? lru_106 : _GEN_5244; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6799 = ~cache_hit ? lru_107 : _GEN_5245; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6800 = ~cache_hit ? lru_108 : _GEN_5246; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6801 = ~cache_hit ? lru_109 : _GEN_5247; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6802 = ~cache_hit ? lru_110 : _GEN_5248; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6803 = ~cache_hit ? lru_111 : _GEN_5249; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6804 = ~cache_hit ? lru_112 : _GEN_5250; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6805 = ~cache_hit ? lru_113 : _GEN_5251; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6806 = ~cache_hit ? lru_114 : _GEN_5252; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6807 = ~cache_hit ? lru_115 : _GEN_5253; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6808 = ~cache_hit ? lru_116 : _GEN_5254; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6809 = ~cache_hit ? lru_117 : _GEN_5255; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6810 = ~cache_hit ? lru_118 : _GEN_5256; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6811 = ~cache_hit ? lru_119 : _GEN_5257; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6812 = ~cache_hit ? lru_120 : _GEN_5258; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6813 = ~cache_hit ? lru_121 : _GEN_5259; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6814 = ~cache_hit ? lru_122 : _GEN_5260; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6815 = ~cache_hit ? lru_123 : _GEN_5261; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6816 = ~cache_hit ? lru_124 : _GEN_5262; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6817 = ~cache_hit ? lru_125 : _GEN_5263; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6818 = ~cache_hit ? lru_126 : _GEN_5264; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6819 = ~cache_hit ? lru_127 : _GEN_5265; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6820 = ~cache_hit ? lru_128 : _GEN_5266; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6821 = ~cache_hit ? lru_129 : _GEN_5267; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6822 = ~cache_hit ? lru_130 : _GEN_5268; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6823 = ~cache_hit ? lru_131 : _GEN_5269; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6824 = ~cache_hit ? lru_132 : _GEN_5270; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6825 = ~cache_hit ? lru_133 : _GEN_5271; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6826 = ~cache_hit ? lru_134 : _GEN_5272; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6827 = ~cache_hit ? lru_135 : _GEN_5273; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6828 = ~cache_hit ? lru_136 : _GEN_5274; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6829 = ~cache_hit ? lru_137 : _GEN_5275; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6830 = ~cache_hit ? lru_138 : _GEN_5276; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6831 = ~cache_hit ? lru_139 : _GEN_5277; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6832 = ~cache_hit ? lru_140 : _GEN_5278; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6833 = ~cache_hit ? lru_141 : _GEN_5279; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6834 = ~cache_hit ? lru_142 : _GEN_5280; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6835 = ~cache_hit ? lru_143 : _GEN_5281; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6836 = ~cache_hit ? lru_144 : _GEN_5282; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6837 = ~cache_hit ? lru_145 : _GEN_5283; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6838 = ~cache_hit ? lru_146 : _GEN_5284; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6839 = ~cache_hit ? lru_147 : _GEN_5285; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6840 = ~cache_hit ? lru_148 : _GEN_5286; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6841 = ~cache_hit ? lru_149 : _GEN_5287; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6842 = ~cache_hit ? lru_150 : _GEN_5288; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6843 = ~cache_hit ? lru_151 : _GEN_5289; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6844 = ~cache_hit ? lru_152 : _GEN_5290; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6845 = ~cache_hit ? lru_153 : _GEN_5291; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6846 = ~cache_hit ? lru_154 : _GEN_5292; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6847 = ~cache_hit ? lru_155 : _GEN_5293; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6848 = ~cache_hit ? lru_156 : _GEN_5294; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6849 = ~cache_hit ? lru_157 : _GEN_5295; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6850 = ~cache_hit ? lru_158 : _GEN_5296; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6851 = ~cache_hit ? lru_159 : _GEN_5297; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6852 = ~cache_hit ? lru_160 : _GEN_5298; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6853 = ~cache_hit ? lru_161 : _GEN_5299; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6854 = ~cache_hit ? lru_162 : _GEN_5300; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6855 = ~cache_hit ? lru_163 : _GEN_5301; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6856 = ~cache_hit ? lru_164 : _GEN_5302; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6857 = ~cache_hit ? lru_165 : _GEN_5303; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6858 = ~cache_hit ? lru_166 : _GEN_5304; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6859 = ~cache_hit ? lru_167 : _GEN_5305; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6860 = ~cache_hit ? lru_168 : _GEN_5306; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6861 = ~cache_hit ? lru_169 : _GEN_5307; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6862 = ~cache_hit ? lru_170 : _GEN_5308; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6863 = ~cache_hit ? lru_171 : _GEN_5309; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6864 = ~cache_hit ? lru_172 : _GEN_5310; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6865 = ~cache_hit ? lru_173 : _GEN_5311; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6866 = ~cache_hit ? lru_174 : _GEN_5312; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6867 = ~cache_hit ? lru_175 : _GEN_5313; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6868 = ~cache_hit ? lru_176 : _GEN_5314; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6869 = ~cache_hit ? lru_177 : _GEN_5315; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6870 = ~cache_hit ? lru_178 : _GEN_5316; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6871 = ~cache_hit ? lru_179 : _GEN_5317; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6872 = ~cache_hit ? lru_180 : _GEN_5318; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6873 = ~cache_hit ? lru_181 : _GEN_5319; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6874 = ~cache_hit ? lru_182 : _GEN_5320; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6875 = ~cache_hit ? lru_183 : _GEN_5321; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6876 = ~cache_hit ? lru_184 : _GEN_5322; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6877 = ~cache_hit ? lru_185 : _GEN_5323; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6878 = ~cache_hit ? lru_186 : _GEN_5324; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6879 = ~cache_hit ? lru_187 : _GEN_5325; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6880 = ~cache_hit ? lru_188 : _GEN_5326; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6881 = ~cache_hit ? lru_189 : _GEN_5327; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6882 = ~cache_hit ? lru_190 : _GEN_5328; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6883 = ~cache_hit ? lru_191 : _GEN_5329; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6884 = ~cache_hit ? lru_192 : _GEN_5330; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6885 = ~cache_hit ? lru_193 : _GEN_5331; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6886 = ~cache_hit ? lru_194 : _GEN_5332; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6887 = ~cache_hit ? lru_195 : _GEN_5333; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6888 = ~cache_hit ? lru_196 : _GEN_5334; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6889 = ~cache_hit ? lru_197 : _GEN_5335; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6890 = ~cache_hit ? lru_198 : _GEN_5336; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6891 = ~cache_hit ? lru_199 : _GEN_5337; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6892 = ~cache_hit ? lru_200 : _GEN_5338; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6893 = ~cache_hit ? lru_201 : _GEN_5339; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6894 = ~cache_hit ? lru_202 : _GEN_5340; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6895 = ~cache_hit ? lru_203 : _GEN_5341; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6896 = ~cache_hit ? lru_204 : _GEN_5342; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6897 = ~cache_hit ? lru_205 : _GEN_5343; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6898 = ~cache_hit ? lru_206 : _GEN_5344; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6899 = ~cache_hit ? lru_207 : _GEN_5345; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6900 = ~cache_hit ? lru_208 : _GEN_5346; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6901 = ~cache_hit ? lru_209 : _GEN_5347; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6902 = ~cache_hit ? lru_210 : _GEN_5348; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6903 = ~cache_hit ? lru_211 : _GEN_5349; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6904 = ~cache_hit ? lru_212 : _GEN_5350; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6905 = ~cache_hit ? lru_213 : _GEN_5351; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6906 = ~cache_hit ? lru_214 : _GEN_5352; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6907 = ~cache_hit ? lru_215 : _GEN_5353; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6908 = ~cache_hit ? lru_216 : _GEN_5354; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6909 = ~cache_hit ? lru_217 : _GEN_5355; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6910 = ~cache_hit ? lru_218 : _GEN_5356; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6911 = ~cache_hit ? lru_219 : _GEN_5357; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6912 = ~cache_hit ? lru_220 : _GEN_5358; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6913 = ~cache_hit ? lru_221 : _GEN_5359; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6914 = ~cache_hit ? lru_222 : _GEN_5360; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6915 = ~cache_hit ? lru_223 : _GEN_5361; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6916 = ~cache_hit ? lru_224 : _GEN_5362; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6917 = ~cache_hit ? lru_225 : _GEN_5363; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6918 = ~cache_hit ? lru_226 : _GEN_5364; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6919 = ~cache_hit ? lru_227 : _GEN_5365; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6920 = ~cache_hit ? lru_228 : _GEN_5366; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6921 = ~cache_hit ? lru_229 : _GEN_5367; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6922 = ~cache_hit ? lru_230 : _GEN_5368; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6923 = ~cache_hit ? lru_231 : _GEN_5369; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6924 = ~cache_hit ? lru_232 : _GEN_5370; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6925 = ~cache_hit ? lru_233 : _GEN_5371; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6926 = ~cache_hit ? lru_234 : _GEN_5372; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6927 = ~cache_hit ? lru_235 : _GEN_5373; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6928 = ~cache_hit ? lru_236 : _GEN_5374; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6929 = ~cache_hit ? lru_237 : _GEN_5375; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6930 = ~cache_hit ? lru_238 : _GEN_5376; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6931 = ~cache_hit ? lru_239 : _GEN_5377; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6932 = ~cache_hit ? lru_240 : _GEN_5378; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6933 = ~cache_hit ? lru_241 : _GEN_5379; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6934 = ~cache_hit ? lru_242 : _GEN_5380; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6935 = ~cache_hit ? lru_243 : _GEN_5381; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6936 = ~cache_hit ? lru_244 : _GEN_5382; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6937 = ~cache_hit ? lru_245 : _GEN_5383; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6938 = ~cache_hit ? lru_246 : _GEN_5384; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6939 = ~cache_hit ? lru_247 : _GEN_5385; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6940 = ~cache_hit ? lru_248 : _GEN_5386; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6941 = ~cache_hit ? lru_249 : _GEN_5387; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6942 = ~cache_hit ? lru_250 : _GEN_5388; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6943 = ~cache_hit ? lru_251 : _GEN_5389; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6944 = ~cache_hit ? lru_252 : _GEN_5390; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6945 = ~cache_hit ? lru_253 : _GEN_5391; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6946 = ~cache_hit ? lru_254 : _GEN_5392; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6947 = ~cache_hit ? lru_255 : _GEN_5393; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6948 = ~cache_hit ? lru_256 : _GEN_5394; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6949 = ~cache_hit ? lru_257 : _GEN_5395; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6950 = ~cache_hit ? lru_258 : _GEN_5396; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6951 = ~cache_hit ? lru_259 : _GEN_5397; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6952 = ~cache_hit ? lru_260 : _GEN_5398; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6953 = ~cache_hit ? lru_261 : _GEN_5399; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6954 = ~cache_hit ? lru_262 : _GEN_5400; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6955 = ~cache_hit ? lru_263 : _GEN_5401; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6956 = ~cache_hit ? lru_264 : _GEN_5402; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6957 = ~cache_hit ? lru_265 : _GEN_5403; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6958 = ~cache_hit ? lru_266 : _GEN_5404; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6959 = ~cache_hit ? lru_267 : _GEN_5405; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6960 = ~cache_hit ? lru_268 : _GEN_5406; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6961 = ~cache_hit ? lru_269 : _GEN_5407; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6962 = ~cache_hit ? lru_270 : _GEN_5408; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6963 = ~cache_hit ? lru_271 : _GEN_5409; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6964 = ~cache_hit ? lru_272 : _GEN_5410; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6965 = ~cache_hit ? lru_273 : _GEN_5411; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6966 = ~cache_hit ? lru_274 : _GEN_5412; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6967 = ~cache_hit ? lru_275 : _GEN_5413; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6968 = ~cache_hit ? lru_276 : _GEN_5414; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6969 = ~cache_hit ? lru_277 : _GEN_5415; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6970 = ~cache_hit ? lru_278 : _GEN_5416; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6971 = ~cache_hit ? lru_279 : _GEN_5417; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6972 = ~cache_hit ? lru_280 : _GEN_5418; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6973 = ~cache_hit ? lru_281 : _GEN_5419; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6974 = ~cache_hit ? lru_282 : _GEN_5420; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6975 = ~cache_hit ? lru_283 : _GEN_5421; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6976 = ~cache_hit ? lru_284 : _GEN_5422; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6977 = ~cache_hit ? lru_285 : _GEN_5423; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6978 = ~cache_hit ? lru_286 : _GEN_5424; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6979 = ~cache_hit ? lru_287 : _GEN_5425; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6980 = ~cache_hit ? lru_288 : _GEN_5426; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6981 = ~cache_hit ? lru_289 : _GEN_5427; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6982 = ~cache_hit ? lru_290 : _GEN_5428; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6983 = ~cache_hit ? lru_291 : _GEN_5429; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6984 = ~cache_hit ? lru_292 : _GEN_5430; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6985 = ~cache_hit ? lru_293 : _GEN_5431; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6986 = ~cache_hit ? lru_294 : _GEN_5432; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6987 = ~cache_hit ? lru_295 : _GEN_5433; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6988 = ~cache_hit ? lru_296 : _GEN_5434; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6989 = ~cache_hit ? lru_297 : _GEN_5435; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6990 = ~cache_hit ? lru_298 : _GEN_5436; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6991 = ~cache_hit ? lru_299 : _GEN_5437; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6992 = ~cache_hit ? lru_300 : _GEN_5438; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6993 = ~cache_hit ? lru_301 : _GEN_5439; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6994 = ~cache_hit ? lru_302 : _GEN_5440; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6995 = ~cache_hit ? lru_303 : _GEN_5441; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6996 = ~cache_hit ? lru_304 : _GEN_5442; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6997 = ~cache_hit ? lru_305 : _GEN_5443; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6998 = ~cache_hit ? lru_306 : _GEN_5444; // @[ICache.scala 175:32 68:20]
  wire  _GEN_6999 = ~cache_hit ? lru_307 : _GEN_5445; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7000 = ~cache_hit ? lru_308 : _GEN_5446; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7001 = ~cache_hit ? lru_309 : _GEN_5447; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7002 = ~cache_hit ? lru_310 : _GEN_5448; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7003 = ~cache_hit ? lru_311 : _GEN_5449; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7004 = ~cache_hit ? lru_312 : _GEN_5450; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7005 = ~cache_hit ? lru_313 : _GEN_5451; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7006 = ~cache_hit ? lru_314 : _GEN_5452; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7007 = ~cache_hit ? lru_315 : _GEN_5453; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7008 = ~cache_hit ? lru_316 : _GEN_5454; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7009 = ~cache_hit ? lru_317 : _GEN_5455; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7010 = ~cache_hit ? lru_318 : _GEN_5456; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7011 = ~cache_hit ? lru_319 : _GEN_5457; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7012 = ~cache_hit ? lru_320 : _GEN_5458; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7013 = ~cache_hit ? lru_321 : _GEN_5459; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7014 = ~cache_hit ? lru_322 : _GEN_5460; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7015 = ~cache_hit ? lru_323 : _GEN_5461; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7016 = ~cache_hit ? lru_324 : _GEN_5462; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7017 = ~cache_hit ? lru_325 : _GEN_5463; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7018 = ~cache_hit ? lru_326 : _GEN_5464; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7019 = ~cache_hit ? lru_327 : _GEN_5465; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7020 = ~cache_hit ? lru_328 : _GEN_5466; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7021 = ~cache_hit ? lru_329 : _GEN_5467; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7022 = ~cache_hit ? lru_330 : _GEN_5468; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7023 = ~cache_hit ? lru_331 : _GEN_5469; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7024 = ~cache_hit ? lru_332 : _GEN_5470; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7025 = ~cache_hit ? lru_333 : _GEN_5471; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7026 = ~cache_hit ? lru_334 : _GEN_5472; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7027 = ~cache_hit ? lru_335 : _GEN_5473; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7028 = ~cache_hit ? lru_336 : _GEN_5474; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7029 = ~cache_hit ? lru_337 : _GEN_5475; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7030 = ~cache_hit ? lru_338 : _GEN_5476; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7031 = ~cache_hit ? lru_339 : _GEN_5477; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7032 = ~cache_hit ? lru_340 : _GEN_5478; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7033 = ~cache_hit ? lru_341 : _GEN_5479; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7034 = ~cache_hit ? lru_342 : _GEN_5480; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7035 = ~cache_hit ? lru_343 : _GEN_5481; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7036 = ~cache_hit ? lru_344 : _GEN_5482; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7037 = ~cache_hit ? lru_345 : _GEN_5483; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7038 = ~cache_hit ? lru_346 : _GEN_5484; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7039 = ~cache_hit ? lru_347 : _GEN_5485; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7040 = ~cache_hit ? lru_348 : _GEN_5486; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7041 = ~cache_hit ? lru_349 : _GEN_5487; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7042 = ~cache_hit ? lru_350 : _GEN_5488; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7043 = ~cache_hit ? lru_351 : _GEN_5489; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7044 = ~cache_hit ? lru_352 : _GEN_5490; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7045 = ~cache_hit ? lru_353 : _GEN_5491; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7046 = ~cache_hit ? lru_354 : _GEN_5492; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7047 = ~cache_hit ? lru_355 : _GEN_5493; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7048 = ~cache_hit ? lru_356 : _GEN_5494; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7049 = ~cache_hit ? lru_357 : _GEN_5495; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7050 = ~cache_hit ? lru_358 : _GEN_5496; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7051 = ~cache_hit ? lru_359 : _GEN_5497; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7052 = ~cache_hit ? lru_360 : _GEN_5498; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7053 = ~cache_hit ? lru_361 : _GEN_5499; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7054 = ~cache_hit ? lru_362 : _GEN_5500; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7055 = ~cache_hit ? lru_363 : _GEN_5501; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7056 = ~cache_hit ? lru_364 : _GEN_5502; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7057 = ~cache_hit ? lru_365 : _GEN_5503; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7058 = ~cache_hit ? lru_366 : _GEN_5504; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7059 = ~cache_hit ? lru_367 : _GEN_5505; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7060 = ~cache_hit ? lru_368 : _GEN_5506; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7061 = ~cache_hit ? lru_369 : _GEN_5507; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7062 = ~cache_hit ? lru_370 : _GEN_5508; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7063 = ~cache_hit ? lru_371 : _GEN_5509; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7064 = ~cache_hit ? lru_372 : _GEN_5510; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7065 = ~cache_hit ? lru_373 : _GEN_5511; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7066 = ~cache_hit ? lru_374 : _GEN_5512; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7067 = ~cache_hit ? lru_375 : _GEN_5513; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7068 = ~cache_hit ? lru_376 : _GEN_5514; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7069 = ~cache_hit ? lru_377 : _GEN_5515; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7070 = ~cache_hit ? lru_378 : _GEN_5516; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7071 = ~cache_hit ? lru_379 : _GEN_5517; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7072 = ~cache_hit ? lru_380 : _GEN_5518; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7073 = ~cache_hit ? lru_381 : _GEN_5519; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7074 = ~cache_hit ? lru_382 : _GEN_5520; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7075 = ~cache_hit ? lru_383 : _GEN_5521; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7076 = ~cache_hit ? lru_384 : _GEN_5522; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7077 = ~cache_hit ? lru_385 : _GEN_5523; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7078 = ~cache_hit ? lru_386 : _GEN_5524; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7079 = ~cache_hit ? lru_387 : _GEN_5525; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7080 = ~cache_hit ? lru_388 : _GEN_5526; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7081 = ~cache_hit ? lru_389 : _GEN_5527; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7082 = ~cache_hit ? lru_390 : _GEN_5528; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7083 = ~cache_hit ? lru_391 : _GEN_5529; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7084 = ~cache_hit ? lru_392 : _GEN_5530; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7085 = ~cache_hit ? lru_393 : _GEN_5531; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7086 = ~cache_hit ? lru_394 : _GEN_5532; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7087 = ~cache_hit ? lru_395 : _GEN_5533; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7088 = ~cache_hit ? lru_396 : _GEN_5534; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7089 = ~cache_hit ? lru_397 : _GEN_5535; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7090 = ~cache_hit ? lru_398 : _GEN_5536; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7091 = ~cache_hit ? lru_399 : _GEN_5537; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7092 = ~cache_hit ? lru_400 : _GEN_5538; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7093 = ~cache_hit ? lru_401 : _GEN_5539; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7094 = ~cache_hit ? lru_402 : _GEN_5540; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7095 = ~cache_hit ? lru_403 : _GEN_5541; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7096 = ~cache_hit ? lru_404 : _GEN_5542; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7097 = ~cache_hit ? lru_405 : _GEN_5543; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7098 = ~cache_hit ? lru_406 : _GEN_5544; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7099 = ~cache_hit ? lru_407 : _GEN_5545; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7100 = ~cache_hit ? lru_408 : _GEN_5546; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7101 = ~cache_hit ? lru_409 : _GEN_5547; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7102 = ~cache_hit ? lru_410 : _GEN_5548; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7103 = ~cache_hit ? lru_411 : _GEN_5549; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7104 = ~cache_hit ? lru_412 : _GEN_5550; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7105 = ~cache_hit ? lru_413 : _GEN_5551; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7106 = ~cache_hit ? lru_414 : _GEN_5552; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7107 = ~cache_hit ? lru_415 : _GEN_5553; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7108 = ~cache_hit ? lru_416 : _GEN_5554; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7109 = ~cache_hit ? lru_417 : _GEN_5555; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7110 = ~cache_hit ? lru_418 : _GEN_5556; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7111 = ~cache_hit ? lru_419 : _GEN_5557; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7112 = ~cache_hit ? lru_420 : _GEN_5558; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7113 = ~cache_hit ? lru_421 : _GEN_5559; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7114 = ~cache_hit ? lru_422 : _GEN_5560; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7115 = ~cache_hit ? lru_423 : _GEN_5561; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7116 = ~cache_hit ? lru_424 : _GEN_5562; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7117 = ~cache_hit ? lru_425 : _GEN_5563; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7118 = ~cache_hit ? lru_426 : _GEN_5564; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7119 = ~cache_hit ? lru_427 : _GEN_5565; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7120 = ~cache_hit ? lru_428 : _GEN_5566; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7121 = ~cache_hit ? lru_429 : _GEN_5567; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7122 = ~cache_hit ? lru_430 : _GEN_5568; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7123 = ~cache_hit ? lru_431 : _GEN_5569; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7124 = ~cache_hit ? lru_432 : _GEN_5570; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7125 = ~cache_hit ? lru_433 : _GEN_5571; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7126 = ~cache_hit ? lru_434 : _GEN_5572; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7127 = ~cache_hit ? lru_435 : _GEN_5573; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7128 = ~cache_hit ? lru_436 : _GEN_5574; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7129 = ~cache_hit ? lru_437 : _GEN_5575; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7130 = ~cache_hit ? lru_438 : _GEN_5576; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7131 = ~cache_hit ? lru_439 : _GEN_5577; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7132 = ~cache_hit ? lru_440 : _GEN_5578; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7133 = ~cache_hit ? lru_441 : _GEN_5579; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7134 = ~cache_hit ? lru_442 : _GEN_5580; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7135 = ~cache_hit ? lru_443 : _GEN_5581; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7136 = ~cache_hit ? lru_444 : _GEN_5582; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7137 = ~cache_hit ? lru_445 : _GEN_5583; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7138 = ~cache_hit ? lru_446 : _GEN_5584; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7139 = ~cache_hit ? lru_447 : _GEN_5585; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7140 = ~cache_hit ? lru_448 : _GEN_5586; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7141 = ~cache_hit ? lru_449 : _GEN_5587; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7142 = ~cache_hit ? lru_450 : _GEN_5588; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7143 = ~cache_hit ? lru_451 : _GEN_5589; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7144 = ~cache_hit ? lru_452 : _GEN_5590; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7145 = ~cache_hit ? lru_453 : _GEN_5591; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7146 = ~cache_hit ? lru_454 : _GEN_5592; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7147 = ~cache_hit ? lru_455 : _GEN_5593; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7148 = ~cache_hit ? lru_456 : _GEN_5594; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7149 = ~cache_hit ? lru_457 : _GEN_5595; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7150 = ~cache_hit ? lru_458 : _GEN_5596; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7151 = ~cache_hit ? lru_459 : _GEN_5597; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7152 = ~cache_hit ? lru_460 : _GEN_5598; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7153 = ~cache_hit ? lru_461 : _GEN_5599; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7154 = ~cache_hit ? lru_462 : _GEN_5600; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7155 = ~cache_hit ? lru_463 : _GEN_5601; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7156 = ~cache_hit ? lru_464 : _GEN_5602; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7157 = ~cache_hit ? lru_465 : _GEN_5603; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7158 = ~cache_hit ? lru_466 : _GEN_5604; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7159 = ~cache_hit ? lru_467 : _GEN_5605; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7160 = ~cache_hit ? lru_468 : _GEN_5606; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7161 = ~cache_hit ? lru_469 : _GEN_5607; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7162 = ~cache_hit ? lru_470 : _GEN_5608; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7163 = ~cache_hit ? lru_471 : _GEN_5609; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7164 = ~cache_hit ? lru_472 : _GEN_5610; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7165 = ~cache_hit ? lru_473 : _GEN_5611; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7166 = ~cache_hit ? lru_474 : _GEN_5612; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7167 = ~cache_hit ? lru_475 : _GEN_5613; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7168 = ~cache_hit ? lru_476 : _GEN_5614; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7169 = ~cache_hit ? lru_477 : _GEN_5615; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7170 = ~cache_hit ? lru_478 : _GEN_5616; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7171 = ~cache_hit ? lru_479 : _GEN_5617; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7172 = ~cache_hit ? lru_480 : _GEN_5618; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7173 = ~cache_hit ? lru_481 : _GEN_5619; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7174 = ~cache_hit ? lru_482 : _GEN_5620; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7175 = ~cache_hit ? lru_483 : _GEN_5621; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7176 = ~cache_hit ? lru_484 : _GEN_5622; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7177 = ~cache_hit ? lru_485 : _GEN_5623; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7178 = ~cache_hit ? lru_486 : _GEN_5624; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7179 = ~cache_hit ? lru_487 : _GEN_5625; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7180 = ~cache_hit ? lru_488 : _GEN_5626; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7181 = ~cache_hit ? lru_489 : _GEN_5627; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7182 = ~cache_hit ? lru_490 : _GEN_5628; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7183 = ~cache_hit ? lru_491 : _GEN_5629; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7184 = ~cache_hit ? lru_492 : _GEN_5630; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7185 = ~cache_hit ? lru_493 : _GEN_5631; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7186 = ~cache_hit ? lru_494 : _GEN_5632; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7187 = ~cache_hit ? lru_495 : _GEN_5633; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7188 = ~cache_hit ? lru_496 : _GEN_5634; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7189 = ~cache_hit ? lru_497 : _GEN_5635; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7190 = ~cache_hit ? lru_498 : _GEN_5636; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7191 = ~cache_hit ? lru_499 : _GEN_5637; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7192 = ~cache_hit ? lru_500 : _GEN_5638; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7193 = ~cache_hit ? lru_501 : _GEN_5639; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7194 = ~cache_hit ? lru_502 : _GEN_5640; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7195 = ~cache_hit ? lru_503 : _GEN_5641; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7196 = ~cache_hit ? lru_504 : _GEN_5642; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7197 = ~cache_hit ? lru_505 : _GEN_5643; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7198 = ~cache_hit ? lru_506 : _GEN_5644; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7199 = ~cache_hit ? lru_507 : _GEN_5645; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7200 = ~cache_hit ? lru_508 : _GEN_5646; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7201 = ~cache_hit ? lru_509 : _GEN_5647; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7202 = ~cache_hit ? lru_510 : _GEN_5648; // @[ICache.scala 175:32 68:20]
  wire  _GEN_7203 = ~cache_hit ? lru_511 : _GEN_5649; // @[ICache.scala 175:32 68:20]
  wire [31:0] _GEN_7204 = ~cache_hit ? saved_1_inst : _GEN_5651; // @[ICache.scala 113:22 175:32]
  wire  _GEN_7205 = ~cache_hit ? saved_0_valid : _GEN_5652; // @[ICache.scala 113:22 175:32]
  wire  _GEN_7206 = ~cache_hit ? saved_1_valid : _GEN_5653; // @[ICache.scala 113:22 175:32]
  wire [2:0] _GEN_7207 = uncached ? 3'h2 : _GEN_5654; // @[ICache.scala 169:30 170:19]
  wire [31:0] _GEN_7208 = uncached ? inst_pa : _GEN_5655; // @[ICache.scala 169:30 171:19]
  wire [7:0] _GEN_7209 = uncached ? 8'h0 : _GEN_5656; // @[ICache.scala 169:30 172:19]
  wire [2:0] _GEN_7210 = uncached ? 3'h2 : _GEN_5657; // @[ICache.scala 169:30 173:19]
  wire  _GEN_7211 = uncached | _GEN_5658; // @[ICache.scala 169:30 174:19]
  wire [5:0] _GEN_7212 = uncached ? rset : _GEN_5659; // @[ICache.scala 169:30 95:21]
  wire [3:0] _GEN_7213 = uncached ? data_wstrb_0_0 : _GEN_5660; // @[ICache.scala 169:30 61:27]
  wire [3:0] _GEN_7214 = uncached ? data_wstrb_1_0 : _GEN_5661; // @[ICache.scala 169:30 61:27]
  wire [3:0] _GEN_7215 = uncached ? data_wstrb_0_1 : _GEN_5662; // @[ICache.scala 169:30 61:27]
  wire [3:0] _GEN_7216 = uncached ? data_wstrb_1_1 : _GEN_5663; // @[ICache.scala 169:30 61:27]
  wire  _GEN_7217 = uncached ? tag_wstrb_0 : _GEN_5664; // @[ICache.scala 169:30 64:26]
  wire  _GEN_7218 = uncached ? tag_wstrb_1 : _GEN_5665; // @[ICache.scala 169:30 64:26]
  wire [19:0] _GEN_7219 = uncached ? tag_wdata : _GEN_5666; // @[ICache.scala 169:30 65:26]
  wire  _GEN_7220 = uncached ? _GEN_1027 : _GEN_5667; // @[ICache.scala 169:30]
  wire  _GEN_7221 = uncached ? _GEN_1539 : _GEN_5668; // @[ICache.scala 169:30]
  wire  _GEN_7222 = uncached ? _GEN_1028 : _GEN_5669; // @[ICache.scala 169:30]
  wire  _GEN_7223 = uncached ? _GEN_1540 : _GEN_5670; // @[ICache.scala 169:30]
  wire  _GEN_7224 = uncached ? _GEN_1029 : _GEN_5671; // @[ICache.scala 169:30]
  wire  _GEN_7225 = uncached ? _GEN_1541 : _GEN_5672; // @[ICache.scala 169:30]
  wire  _GEN_7226 = uncached ? _GEN_1030 : _GEN_5673; // @[ICache.scala 169:30]
  wire  _GEN_7227 = uncached ? _GEN_1542 : _GEN_5674; // @[ICache.scala 169:30]
  wire  _GEN_7228 = uncached ? _GEN_1031 : _GEN_5675; // @[ICache.scala 169:30]
  wire  _GEN_7229 = uncached ? _GEN_1543 : _GEN_5676; // @[ICache.scala 169:30]
  wire  _GEN_7230 = uncached ? _GEN_1032 : _GEN_5677; // @[ICache.scala 169:30]
  wire  _GEN_7231 = uncached ? _GEN_1544 : _GEN_5678; // @[ICache.scala 169:30]
  wire  _GEN_7232 = uncached ? _GEN_1033 : _GEN_5679; // @[ICache.scala 169:30]
  wire  _GEN_7233 = uncached ? _GEN_1545 : _GEN_5680; // @[ICache.scala 169:30]
  wire  _GEN_7234 = uncached ? _GEN_1034 : _GEN_5681; // @[ICache.scala 169:30]
  wire  _GEN_7235 = uncached ? _GEN_1546 : _GEN_5682; // @[ICache.scala 169:30]
  wire  _GEN_7236 = uncached ? _GEN_1035 : _GEN_5683; // @[ICache.scala 169:30]
  wire  _GEN_7237 = uncached ? _GEN_1547 : _GEN_5684; // @[ICache.scala 169:30]
  wire  _GEN_7238 = uncached ? _GEN_1036 : _GEN_5685; // @[ICache.scala 169:30]
  wire  _GEN_7239 = uncached ? _GEN_1548 : _GEN_5686; // @[ICache.scala 169:30]
  wire  _GEN_7240 = uncached ? _GEN_1037 : _GEN_5687; // @[ICache.scala 169:30]
  wire  _GEN_7241 = uncached ? _GEN_1549 : _GEN_5688; // @[ICache.scala 169:30]
  wire  _GEN_7242 = uncached ? _GEN_1038 : _GEN_5689; // @[ICache.scala 169:30]
  wire  _GEN_7243 = uncached ? _GEN_1550 : _GEN_5690; // @[ICache.scala 169:30]
  wire  _GEN_7244 = uncached ? _GEN_1039 : _GEN_5691; // @[ICache.scala 169:30]
  wire  _GEN_7245 = uncached ? _GEN_1551 : _GEN_5692; // @[ICache.scala 169:30]
  wire  _GEN_7246 = uncached ? _GEN_1040 : _GEN_5693; // @[ICache.scala 169:30]
  wire  _GEN_7247 = uncached ? _GEN_1552 : _GEN_5694; // @[ICache.scala 169:30]
  wire  _GEN_7248 = uncached ? _GEN_1041 : _GEN_5695; // @[ICache.scala 169:30]
  wire  _GEN_7249 = uncached ? _GEN_1553 : _GEN_5696; // @[ICache.scala 169:30]
  wire  _GEN_7250 = uncached ? _GEN_1042 : _GEN_5697; // @[ICache.scala 169:30]
  wire  _GEN_7251 = uncached ? _GEN_1554 : _GEN_5698; // @[ICache.scala 169:30]
  wire  _GEN_7252 = uncached ? _GEN_1043 : _GEN_5699; // @[ICache.scala 169:30]
  wire  _GEN_7253 = uncached ? _GEN_1555 : _GEN_5700; // @[ICache.scala 169:30]
  wire  _GEN_7254 = uncached ? _GEN_1044 : _GEN_5701; // @[ICache.scala 169:30]
  wire  _GEN_7255 = uncached ? _GEN_1556 : _GEN_5702; // @[ICache.scala 169:30]
  wire  _GEN_7256 = uncached ? _GEN_1045 : _GEN_5703; // @[ICache.scala 169:30]
  wire  _GEN_7257 = uncached ? _GEN_1557 : _GEN_5704; // @[ICache.scala 169:30]
  wire  _GEN_7258 = uncached ? _GEN_1046 : _GEN_5705; // @[ICache.scala 169:30]
  wire  _GEN_7259 = uncached ? _GEN_1558 : _GEN_5706; // @[ICache.scala 169:30]
  wire  _GEN_7260 = uncached ? _GEN_1047 : _GEN_5707; // @[ICache.scala 169:30]
  wire  _GEN_7261 = uncached ? _GEN_1559 : _GEN_5708; // @[ICache.scala 169:30]
  wire  _GEN_7262 = uncached ? _GEN_1048 : _GEN_5709; // @[ICache.scala 169:30]
  wire  _GEN_7263 = uncached ? _GEN_1560 : _GEN_5710; // @[ICache.scala 169:30]
  wire  _GEN_7264 = uncached ? _GEN_1049 : _GEN_5711; // @[ICache.scala 169:30]
  wire  _GEN_7265 = uncached ? _GEN_1561 : _GEN_5712; // @[ICache.scala 169:30]
  wire  _GEN_7266 = uncached ? _GEN_1050 : _GEN_5713; // @[ICache.scala 169:30]
  wire  _GEN_7267 = uncached ? _GEN_1562 : _GEN_5714; // @[ICache.scala 169:30]
  wire  _GEN_7268 = uncached ? _GEN_1051 : _GEN_5715; // @[ICache.scala 169:30]
  wire  _GEN_7269 = uncached ? _GEN_1563 : _GEN_5716; // @[ICache.scala 169:30]
  wire  _GEN_7270 = uncached ? _GEN_1052 : _GEN_5717; // @[ICache.scala 169:30]
  wire  _GEN_7271 = uncached ? _GEN_1564 : _GEN_5718; // @[ICache.scala 169:30]
  wire  _GEN_7272 = uncached ? _GEN_1053 : _GEN_5719; // @[ICache.scala 169:30]
  wire  _GEN_7273 = uncached ? _GEN_1565 : _GEN_5720; // @[ICache.scala 169:30]
  wire  _GEN_7274 = uncached ? _GEN_1054 : _GEN_5721; // @[ICache.scala 169:30]
  wire  _GEN_7275 = uncached ? _GEN_1566 : _GEN_5722; // @[ICache.scala 169:30]
  wire  _GEN_7276 = uncached ? _GEN_1055 : _GEN_5723; // @[ICache.scala 169:30]
  wire  _GEN_7277 = uncached ? _GEN_1567 : _GEN_5724; // @[ICache.scala 169:30]
  wire  _GEN_7278 = uncached ? _GEN_1056 : _GEN_5725; // @[ICache.scala 169:30]
  wire  _GEN_7279 = uncached ? _GEN_1568 : _GEN_5726; // @[ICache.scala 169:30]
  wire  _GEN_7280 = uncached ? _GEN_1057 : _GEN_5727; // @[ICache.scala 169:30]
  wire  _GEN_7281 = uncached ? _GEN_1569 : _GEN_5728; // @[ICache.scala 169:30]
  wire  _GEN_7282 = uncached ? _GEN_1058 : _GEN_5729; // @[ICache.scala 169:30]
  wire  _GEN_7283 = uncached ? _GEN_1570 : _GEN_5730; // @[ICache.scala 169:30]
  wire  _GEN_7284 = uncached ? _GEN_1059 : _GEN_5731; // @[ICache.scala 169:30]
  wire  _GEN_7285 = uncached ? _GEN_1571 : _GEN_5732; // @[ICache.scala 169:30]
  wire  _GEN_7286 = uncached ? _GEN_1060 : _GEN_5733; // @[ICache.scala 169:30]
  wire  _GEN_7287 = uncached ? _GEN_1572 : _GEN_5734; // @[ICache.scala 169:30]
  wire  _GEN_7288 = uncached ? _GEN_1061 : _GEN_5735; // @[ICache.scala 169:30]
  wire  _GEN_7289 = uncached ? _GEN_1573 : _GEN_5736; // @[ICache.scala 169:30]
  wire  _GEN_7290 = uncached ? _GEN_1062 : _GEN_5737; // @[ICache.scala 169:30]
  wire  _GEN_7291 = uncached ? _GEN_1574 : _GEN_5738; // @[ICache.scala 169:30]
  wire  _GEN_7292 = uncached ? _GEN_1063 : _GEN_5739; // @[ICache.scala 169:30]
  wire  _GEN_7293 = uncached ? _GEN_1575 : _GEN_5740; // @[ICache.scala 169:30]
  wire  _GEN_7294 = uncached ? _GEN_1064 : _GEN_5741; // @[ICache.scala 169:30]
  wire  _GEN_7295 = uncached ? _GEN_1576 : _GEN_5742; // @[ICache.scala 169:30]
  wire  _GEN_7296 = uncached ? _GEN_1065 : _GEN_5743; // @[ICache.scala 169:30]
  wire  _GEN_7297 = uncached ? _GEN_1577 : _GEN_5744; // @[ICache.scala 169:30]
  wire  _GEN_7298 = uncached ? _GEN_1066 : _GEN_5745; // @[ICache.scala 169:30]
  wire  _GEN_7299 = uncached ? _GEN_1578 : _GEN_5746; // @[ICache.scala 169:30]
  wire  _GEN_7300 = uncached ? _GEN_1067 : _GEN_5747; // @[ICache.scala 169:30]
  wire  _GEN_7301 = uncached ? _GEN_1579 : _GEN_5748; // @[ICache.scala 169:30]
  wire  _GEN_7302 = uncached ? _GEN_1068 : _GEN_5749; // @[ICache.scala 169:30]
  wire  _GEN_7303 = uncached ? _GEN_1580 : _GEN_5750; // @[ICache.scala 169:30]
  wire  _GEN_7304 = uncached ? _GEN_1069 : _GEN_5751; // @[ICache.scala 169:30]
  wire  _GEN_7305 = uncached ? _GEN_1581 : _GEN_5752; // @[ICache.scala 169:30]
  wire  _GEN_7306 = uncached ? _GEN_1070 : _GEN_5753; // @[ICache.scala 169:30]
  wire  _GEN_7307 = uncached ? _GEN_1582 : _GEN_5754; // @[ICache.scala 169:30]
  wire  _GEN_7308 = uncached ? _GEN_1071 : _GEN_5755; // @[ICache.scala 169:30]
  wire  _GEN_7309 = uncached ? _GEN_1583 : _GEN_5756; // @[ICache.scala 169:30]
  wire  _GEN_7310 = uncached ? _GEN_1072 : _GEN_5757; // @[ICache.scala 169:30]
  wire  _GEN_7311 = uncached ? _GEN_1584 : _GEN_5758; // @[ICache.scala 169:30]
  wire  _GEN_7312 = uncached ? _GEN_1073 : _GEN_5759; // @[ICache.scala 169:30]
  wire  _GEN_7313 = uncached ? _GEN_1585 : _GEN_5760; // @[ICache.scala 169:30]
  wire  _GEN_7314 = uncached ? _GEN_1074 : _GEN_5761; // @[ICache.scala 169:30]
  wire  _GEN_7315 = uncached ? _GEN_1586 : _GEN_5762; // @[ICache.scala 169:30]
  wire  _GEN_7316 = uncached ? _GEN_1075 : _GEN_5763; // @[ICache.scala 169:30]
  wire  _GEN_7317 = uncached ? _GEN_1587 : _GEN_5764; // @[ICache.scala 169:30]
  wire  _GEN_7318 = uncached ? _GEN_1076 : _GEN_5765; // @[ICache.scala 169:30]
  wire  _GEN_7319 = uncached ? _GEN_1588 : _GEN_5766; // @[ICache.scala 169:30]
  wire  _GEN_7320 = uncached ? _GEN_1077 : _GEN_5767; // @[ICache.scala 169:30]
  wire  _GEN_7321 = uncached ? _GEN_1589 : _GEN_5768; // @[ICache.scala 169:30]
  wire  _GEN_7322 = uncached ? _GEN_1078 : _GEN_5769; // @[ICache.scala 169:30]
  wire  _GEN_7323 = uncached ? _GEN_1590 : _GEN_5770; // @[ICache.scala 169:30]
  wire  _GEN_7324 = uncached ? _GEN_1079 : _GEN_5771; // @[ICache.scala 169:30]
  wire  _GEN_7325 = uncached ? _GEN_1591 : _GEN_5772; // @[ICache.scala 169:30]
  wire  _GEN_7326 = uncached ? _GEN_1080 : _GEN_5773; // @[ICache.scala 169:30]
  wire  _GEN_7327 = uncached ? _GEN_1592 : _GEN_5774; // @[ICache.scala 169:30]
  wire  _GEN_7328 = uncached ? _GEN_1081 : _GEN_5775; // @[ICache.scala 169:30]
  wire  _GEN_7329 = uncached ? _GEN_1593 : _GEN_5776; // @[ICache.scala 169:30]
  wire  _GEN_7330 = uncached ? _GEN_1082 : _GEN_5777; // @[ICache.scala 169:30]
  wire  _GEN_7331 = uncached ? _GEN_1594 : _GEN_5778; // @[ICache.scala 169:30]
  wire  _GEN_7332 = uncached ? _GEN_1083 : _GEN_5779; // @[ICache.scala 169:30]
  wire  _GEN_7333 = uncached ? _GEN_1595 : _GEN_5780; // @[ICache.scala 169:30]
  wire  _GEN_7334 = uncached ? _GEN_1084 : _GEN_5781; // @[ICache.scala 169:30]
  wire  _GEN_7335 = uncached ? _GEN_1596 : _GEN_5782; // @[ICache.scala 169:30]
  wire  _GEN_7336 = uncached ? _GEN_1085 : _GEN_5783; // @[ICache.scala 169:30]
  wire  _GEN_7337 = uncached ? _GEN_1597 : _GEN_5784; // @[ICache.scala 169:30]
  wire  _GEN_7338 = uncached ? _GEN_1086 : _GEN_5785; // @[ICache.scala 169:30]
  wire  _GEN_7339 = uncached ? _GEN_1598 : _GEN_5786; // @[ICache.scala 169:30]
  wire  _GEN_7340 = uncached ? _GEN_1087 : _GEN_5787; // @[ICache.scala 169:30]
  wire  _GEN_7341 = uncached ? _GEN_1599 : _GEN_5788; // @[ICache.scala 169:30]
  wire  _GEN_7342 = uncached ? _GEN_1088 : _GEN_5789; // @[ICache.scala 169:30]
  wire  _GEN_7343 = uncached ? _GEN_1600 : _GEN_5790; // @[ICache.scala 169:30]
  wire  _GEN_7344 = uncached ? _GEN_1089 : _GEN_5791; // @[ICache.scala 169:30]
  wire  _GEN_7345 = uncached ? _GEN_1601 : _GEN_5792; // @[ICache.scala 169:30]
  wire  _GEN_7346 = uncached ? _GEN_1090 : _GEN_5793; // @[ICache.scala 169:30]
  wire  _GEN_7347 = uncached ? _GEN_1602 : _GEN_5794; // @[ICache.scala 169:30]
  wire  _GEN_7348 = uncached ? _GEN_1091 : _GEN_5795; // @[ICache.scala 169:30]
  wire  _GEN_7349 = uncached ? _GEN_1603 : _GEN_5796; // @[ICache.scala 169:30]
  wire  _GEN_7350 = uncached ? _GEN_1092 : _GEN_5797; // @[ICache.scala 169:30]
  wire  _GEN_7351 = uncached ? _GEN_1604 : _GEN_5798; // @[ICache.scala 169:30]
  wire  _GEN_7352 = uncached ? _GEN_1093 : _GEN_5799; // @[ICache.scala 169:30]
  wire  _GEN_7353 = uncached ? _GEN_1605 : _GEN_5800; // @[ICache.scala 169:30]
  wire  _GEN_7354 = uncached ? _GEN_1094 : _GEN_5801; // @[ICache.scala 169:30]
  wire  _GEN_7355 = uncached ? _GEN_1606 : _GEN_5802; // @[ICache.scala 169:30]
  wire  _GEN_7356 = uncached ? _GEN_1095 : _GEN_5803; // @[ICache.scala 169:30]
  wire  _GEN_7357 = uncached ? _GEN_1607 : _GEN_5804; // @[ICache.scala 169:30]
  wire  _GEN_7358 = uncached ? _GEN_1096 : _GEN_5805; // @[ICache.scala 169:30]
  wire  _GEN_7359 = uncached ? _GEN_1608 : _GEN_5806; // @[ICache.scala 169:30]
  wire  _GEN_7360 = uncached ? _GEN_1097 : _GEN_5807; // @[ICache.scala 169:30]
  wire  _GEN_7361 = uncached ? _GEN_1609 : _GEN_5808; // @[ICache.scala 169:30]
  wire  _GEN_7362 = uncached ? _GEN_1098 : _GEN_5809; // @[ICache.scala 169:30]
  wire  _GEN_7363 = uncached ? _GEN_1610 : _GEN_5810; // @[ICache.scala 169:30]
  wire  _GEN_7364 = uncached ? _GEN_1099 : _GEN_5811; // @[ICache.scala 169:30]
  wire  _GEN_7365 = uncached ? _GEN_1611 : _GEN_5812; // @[ICache.scala 169:30]
  wire  _GEN_7366 = uncached ? _GEN_1100 : _GEN_5813; // @[ICache.scala 169:30]
  wire  _GEN_7367 = uncached ? _GEN_1612 : _GEN_5814; // @[ICache.scala 169:30]
  wire  _GEN_7368 = uncached ? _GEN_1101 : _GEN_5815; // @[ICache.scala 169:30]
  wire  _GEN_7369 = uncached ? _GEN_1613 : _GEN_5816; // @[ICache.scala 169:30]
  wire  _GEN_7370 = uncached ? _GEN_1102 : _GEN_5817; // @[ICache.scala 169:30]
  wire  _GEN_7371 = uncached ? _GEN_1614 : _GEN_5818; // @[ICache.scala 169:30]
  wire  _GEN_7372 = uncached ? _GEN_1103 : _GEN_5819; // @[ICache.scala 169:30]
  wire  _GEN_7373 = uncached ? _GEN_1615 : _GEN_5820; // @[ICache.scala 169:30]
  wire  _GEN_7374 = uncached ? _GEN_1104 : _GEN_5821; // @[ICache.scala 169:30]
  wire  _GEN_7375 = uncached ? _GEN_1616 : _GEN_5822; // @[ICache.scala 169:30]
  wire  _GEN_7376 = uncached ? _GEN_1105 : _GEN_5823; // @[ICache.scala 169:30]
  wire  _GEN_7377 = uncached ? _GEN_1617 : _GEN_5824; // @[ICache.scala 169:30]
  wire  _GEN_7378 = uncached ? _GEN_1106 : _GEN_5825; // @[ICache.scala 169:30]
  wire  _GEN_7379 = uncached ? _GEN_1618 : _GEN_5826; // @[ICache.scala 169:30]
  wire  _GEN_7380 = uncached ? _GEN_1107 : _GEN_5827; // @[ICache.scala 169:30]
  wire  _GEN_7381 = uncached ? _GEN_1619 : _GEN_5828; // @[ICache.scala 169:30]
  wire  _GEN_7382 = uncached ? _GEN_1108 : _GEN_5829; // @[ICache.scala 169:30]
  wire  _GEN_7383 = uncached ? _GEN_1620 : _GEN_5830; // @[ICache.scala 169:30]
  wire  _GEN_7384 = uncached ? _GEN_1109 : _GEN_5831; // @[ICache.scala 169:30]
  wire  _GEN_7385 = uncached ? _GEN_1621 : _GEN_5832; // @[ICache.scala 169:30]
  wire  _GEN_7386 = uncached ? _GEN_1110 : _GEN_5833; // @[ICache.scala 169:30]
  wire  _GEN_7387 = uncached ? _GEN_1622 : _GEN_5834; // @[ICache.scala 169:30]
  wire  _GEN_7388 = uncached ? _GEN_1111 : _GEN_5835; // @[ICache.scala 169:30]
  wire  _GEN_7389 = uncached ? _GEN_1623 : _GEN_5836; // @[ICache.scala 169:30]
  wire  _GEN_7390 = uncached ? _GEN_1112 : _GEN_5837; // @[ICache.scala 169:30]
  wire  _GEN_7391 = uncached ? _GEN_1624 : _GEN_5838; // @[ICache.scala 169:30]
  wire  _GEN_7392 = uncached ? _GEN_1113 : _GEN_5839; // @[ICache.scala 169:30]
  wire  _GEN_7393 = uncached ? _GEN_1625 : _GEN_5840; // @[ICache.scala 169:30]
  wire  _GEN_7394 = uncached ? _GEN_1114 : _GEN_5841; // @[ICache.scala 169:30]
  wire  _GEN_7395 = uncached ? _GEN_1626 : _GEN_5842; // @[ICache.scala 169:30]
  wire  _GEN_7396 = uncached ? _GEN_1115 : _GEN_5843; // @[ICache.scala 169:30]
  wire  _GEN_7397 = uncached ? _GEN_1627 : _GEN_5844; // @[ICache.scala 169:30]
  wire  _GEN_7398 = uncached ? _GEN_1116 : _GEN_5845; // @[ICache.scala 169:30]
  wire  _GEN_7399 = uncached ? _GEN_1628 : _GEN_5846; // @[ICache.scala 169:30]
  wire  _GEN_7400 = uncached ? _GEN_1117 : _GEN_5847; // @[ICache.scala 169:30]
  wire  _GEN_7401 = uncached ? _GEN_1629 : _GEN_5848; // @[ICache.scala 169:30]
  wire  _GEN_7402 = uncached ? _GEN_1118 : _GEN_5849; // @[ICache.scala 169:30]
  wire  _GEN_7403 = uncached ? _GEN_1630 : _GEN_5850; // @[ICache.scala 169:30]
  wire  _GEN_7404 = uncached ? _GEN_1119 : _GEN_5851; // @[ICache.scala 169:30]
  wire  _GEN_7405 = uncached ? _GEN_1631 : _GEN_5852; // @[ICache.scala 169:30]
  wire  _GEN_7406 = uncached ? _GEN_1120 : _GEN_5853; // @[ICache.scala 169:30]
  wire  _GEN_7407 = uncached ? _GEN_1632 : _GEN_5854; // @[ICache.scala 169:30]
  wire  _GEN_7408 = uncached ? _GEN_1121 : _GEN_5855; // @[ICache.scala 169:30]
  wire  _GEN_7409 = uncached ? _GEN_1633 : _GEN_5856; // @[ICache.scala 169:30]
  wire  _GEN_7410 = uncached ? _GEN_1122 : _GEN_5857; // @[ICache.scala 169:30]
  wire  _GEN_7411 = uncached ? _GEN_1634 : _GEN_5858; // @[ICache.scala 169:30]
  wire  _GEN_7412 = uncached ? _GEN_1123 : _GEN_5859; // @[ICache.scala 169:30]
  wire  _GEN_7413 = uncached ? _GEN_1635 : _GEN_5860; // @[ICache.scala 169:30]
  wire  _GEN_7414 = uncached ? _GEN_1124 : _GEN_5861; // @[ICache.scala 169:30]
  wire  _GEN_7415 = uncached ? _GEN_1636 : _GEN_5862; // @[ICache.scala 169:30]
  wire  _GEN_7416 = uncached ? _GEN_1125 : _GEN_5863; // @[ICache.scala 169:30]
  wire  _GEN_7417 = uncached ? _GEN_1637 : _GEN_5864; // @[ICache.scala 169:30]
  wire  _GEN_7418 = uncached ? _GEN_1126 : _GEN_5865; // @[ICache.scala 169:30]
  wire  _GEN_7419 = uncached ? _GEN_1638 : _GEN_5866; // @[ICache.scala 169:30]
  wire  _GEN_7420 = uncached ? _GEN_1127 : _GEN_5867; // @[ICache.scala 169:30]
  wire  _GEN_7421 = uncached ? _GEN_1639 : _GEN_5868; // @[ICache.scala 169:30]
  wire  _GEN_7422 = uncached ? _GEN_1128 : _GEN_5869; // @[ICache.scala 169:30]
  wire  _GEN_7423 = uncached ? _GEN_1640 : _GEN_5870; // @[ICache.scala 169:30]
  wire  _GEN_7424 = uncached ? _GEN_1129 : _GEN_5871; // @[ICache.scala 169:30]
  wire  _GEN_7425 = uncached ? _GEN_1641 : _GEN_5872; // @[ICache.scala 169:30]
  wire  _GEN_7426 = uncached ? _GEN_1130 : _GEN_5873; // @[ICache.scala 169:30]
  wire  _GEN_7427 = uncached ? _GEN_1642 : _GEN_5874; // @[ICache.scala 169:30]
  wire  _GEN_7428 = uncached ? _GEN_1131 : _GEN_5875; // @[ICache.scala 169:30]
  wire  _GEN_7429 = uncached ? _GEN_1643 : _GEN_5876; // @[ICache.scala 169:30]
  wire  _GEN_7430 = uncached ? _GEN_1132 : _GEN_5877; // @[ICache.scala 169:30]
  wire  _GEN_7431 = uncached ? _GEN_1644 : _GEN_5878; // @[ICache.scala 169:30]
  wire  _GEN_7432 = uncached ? _GEN_1133 : _GEN_5879; // @[ICache.scala 169:30]
  wire  _GEN_7433 = uncached ? _GEN_1645 : _GEN_5880; // @[ICache.scala 169:30]
  wire  _GEN_7434 = uncached ? _GEN_1134 : _GEN_5881; // @[ICache.scala 169:30]
  wire  _GEN_7435 = uncached ? _GEN_1646 : _GEN_5882; // @[ICache.scala 169:30]
  wire  _GEN_7436 = uncached ? _GEN_1135 : _GEN_5883; // @[ICache.scala 169:30]
  wire  _GEN_7437 = uncached ? _GEN_1647 : _GEN_5884; // @[ICache.scala 169:30]
  wire  _GEN_7438 = uncached ? _GEN_1136 : _GEN_5885; // @[ICache.scala 169:30]
  wire  _GEN_7439 = uncached ? _GEN_1648 : _GEN_5886; // @[ICache.scala 169:30]
  wire  _GEN_7440 = uncached ? _GEN_1137 : _GEN_5887; // @[ICache.scala 169:30]
  wire  _GEN_7441 = uncached ? _GEN_1649 : _GEN_5888; // @[ICache.scala 169:30]
  wire  _GEN_7442 = uncached ? _GEN_1138 : _GEN_5889; // @[ICache.scala 169:30]
  wire  _GEN_7443 = uncached ? _GEN_1650 : _GEN_5890; // @[ICache.scala 169:30]
  wire  _GEN_7444 = uncached ? _GEN_1139 : _GEN_5891; // @[ICache.scala 169:30]
  wire  _GEN_7445 = uncached ? _GEN_1651 : _GEN_5892; // @[ICache.scala 169:30]
  wire  _GEN_7446 = uncached ? _GEN_1140 : _GEN_5893; // @[ICache.scala 169:30]
  wire  _GEN_7447 = uncached ? _GEN_1652 : _GEN_5894; // @[ICache.scala 169:30]
  wire  _GEN_7448 = uncached ? _GEN_1141 : _GEN_5895; // @[ICache.scala 169:30]
  wire  _GEN_7449 = uncached ? _GEN_1653 : _GEN_5896; // @[ICache.scala 169:30]
  wire  _GEN_7450 = uncached ? _GEN_1142 : _GEN_5897; // @[ICache.scala 169:30]
  wire  _GEN_7451 = uncached ? _GEN_1654 : _GEN_5898; // @[ICache.scala 169:30]
  wire  _GEN_7452 = uncached ? _GEN_1143 : _GEN_5899; // @[ICache.scala 169:30]
  wire  _GEN_7453 = uncached ? _GEN_1655 : _GEN_5900; // @[ICache.scala 169:30]
  wire  _GEN_7454 = uncached ? _GEN_1144 : _GEN_5901; // @[ICache.scala 169:30]
  wire  _GEN_7455 = uncached ? _GEN_1656 : _GEN_5902; // @[ICache.scala 169:30]
  wire  _GEN_7456 = uncached ? _GEN_1145 : _GEN_5903; // @[ICache.scala 169:30]
  wire  _GEN_7457 = uncached ? _GEN_1657 : _GEN_5904; // @[ICache.scala 169:30]
  wire  _GEN_7458 = uncached ? _GEN_1146 : _GEN_5905; // @[ICache.scala 169:30]
  wire  _GEN_7459 = uncached ? _GEN_1658 : _GEN_5906; // @[ICache.scala 169:30]
  wire  _GEN_7460 = uncached ? _GEN_1147 : _GEN_5907; // @[ICache.scala 169:30]
  wire  _GEN_7461 = uncached ? _GEN_1659 : _GEN_5908; // @[ICache.scala 169:30]
  wire  _GEN_7462 = uncached ? _GEN_1148 : _GEN_5909; // @[ICache.scala 169:30]
  wire  _GEN_7463 = uncached ? _GEN_1660 : _GEN_5910; // @[ICache.scala 169:30]
  wire  _GEN_7464 = uncached ? _GEN_1149 : _GEN_5911; // @[ICache.scala 169:30]
  wire  _GEN_7465 = uncached ? _GEN_1661 : _GEN_5912; // @[ICache.scala 169:30]
  wire  _GEN_7466 = uncached ? _GEN_1150 : _GEN_5913; // @[ICache.scala 169:30]
  wire  _GEN_7467 = uncached ? _GEN_1662 : _GEN_5914; // @[ICache.scala 169:30]
  wire  _GEN_7468 = uncached ? _GEN_1151 : _GEN_5915; // @[ICache.scala 169:30]
  wire  _GEN_7469 = uncached ? _GEN_1663 : _GEN_5916; // @[ICache.scala 169:30]
  wire  _GEN_7470 = uncached ? _GEN_1152 : _GEN_5917; // @[ICache.scala 169:30]
  wire  _GEN_7471 = uncached ? _GEN_1664 : _GEN_5918; // @[ICache.scala 169:30]
  wire  _GEN_7472 = uncached ? _GEN_1153 : _GEN_5919; // @[ICache.scala 169:30]
  wire  _GEN_7473 = uncached ? _GEN_1665 : _GEN_5920; // @[ICache.scala 169:30]
  wire  _GEN_7474 = uncached ? _GEN_1154 : _GEN_5921; // @[ICache.scala 169:30]
  wire  _GEN_7475 = uncached ? _GEN_1666 : _GEN_5922; // @[ICache.scala 169:30]
  wire  _GEN_7476 = uncached ? _GEN_1155 : _GEN_5923; // @[ICache.scala 169:30]
  wire  _GEN_7477 = uncached ? _GEN_1667 : _GEN_5924; // @[ICache.scala 169:30]
  wire  _GEN_7478 = uncached ? _GEN_1156 : _GEN_5925; // @[ICache.scala 169:30]
  wire  _GEN_7479 = uncached ? _GEN_1668 : _GEN_5926; // @[ICache.scala 169:30]
  wire  _GEN_7480 = uncached ? _GEN_1157 : _GEN_5927; // @[ICache.scala 169:30]
  wire  _GEN_7481 = uncached ? _GEN_1669 : _GEN_5928; // @[ICache.scala 169:30]
  wire  _GEN_7482 = uncached ? _GEN_1158 : _GEN_5929; // @[ICache.scala 169:30]
  wire  _GEN_7483 = uncached ? _GEN_1670 : _GEN_5930; // @[ICache.scala 169:30]
  wire  _GEN_7484 = uncached ? _GEN_1159 : _GEN_5931; // @[ICache.scala 169:30]
  wire  _GEN_7485 = uncached ? _GEN_1671 : _GEN_5932; // @[ICache.scala 169:30]
  wire  _GEN_7486 = uncached ? _GEN_1160 : _GEN_5933; // @[ICache.scala 169:30]
  wire  _GEN_7487 = uncached ? _GEN_1672 : _GEN_5934; // @[ICache.scala 169:30]
  wire  _GEN_7488 = uncached ? _GEN_1161 : _GEN_5935; // @[ICache.scala 169:30]
  wire  _GEN_7489 = uncached ? _GEN_1673 : _GEN_5936; // @[ICache.scala 169:30]
  wire  _GEN_7490 = uncached ? _GEN_1162 : _GEN_5937; // @[ICache.scala 169:30]
  wire  _GEN_7491 = uncached ? _GEN_1674 : _GEN_5938; // @[ICache.scala 169:30]
  wire  _GEN_7492 = uncached ? _GEN_1163 : _GEN_5939; // @[ICache.scala 169:30]
  wire  _GEN_7493 = uncached ? _GEN_1675 : _GEN_5940; // @[ICache.scala 169:30]
  wire  _GEN_7494 = uncached ? _GEN_1164 : _GEN_5941; // @[ICache.scala 169:30]
  wire  _GEN_7495 = uncached ? _GEN_1676 : _GEN_5942; // @[ICache.scala 169:30]
  wire  _GEN_7496 = uncached ? _GEN_1165 : _GEN_5943; // @[ICache.scala 169:30]
  wire  _GEN_7497 = uncached ? _GEN_1677 : _GEN_5944; // @[ICache.scala 169:30]
  wire  _GEN_7498 = uncached ? _GEN_1166 : _GEN_5945; // @[ICache.scala 169:30]
  wire  _GEN_7499 = uncached ? _GEN_1678 : _GEN_5946; // @[ICache.scala 169:30]
  wire  _GEN_7500 = uncached ? _GEN_1167 : _GEN_5947; // @[ICache.scala 169:30]
  wire  _GEN_7501 = uncached ? _GEN_1679 : _GEN_5948; // @[ICache.scala 169:30]
  wire  _GEN_7502 = uncached ? _GEN_1168 : _GEN_5949; // @[ICache.scala 169:30]
  wire  _GEN_7503 = uncached ? _GEN_1680 : _GEN_5950; // @[ICache.scala 169:30]
  wire  _GEN_7504 = uncached ? _GEN_1169 : _GEN_5951; // @[ICache.scala 169:30]
  wire  _GEN_7505 = uncached ? _GEN_1681 : _GEN_5952; // @[ICache.scala 169:30]
  wire  _GEN_7506 = uncached ? _GEN_1170 : _GEN_5953; // @[ICache.scala 169:30]
  wire  _GEN_7507 = uncached ? _GEN_1682 : _GEN_5954; // @[ICache.scala 169:30]
  wire  _GEN_7508 = uncached ? _GEN_1171 : _GEN_5955; // @[ICache.scala 169:30]
  wire  _GEN_7509 = uncached ? _GEN_1683 : _GEN_5956; // @[ICache.scala 169:30]
  wire  _GEN_7510 = uncached ? _GEN_1172 : _GEN_5957; // @[ICache.scala 169:30]
  wire  _GEN_7511 = uncached ? _GEN_1684 : _GEN_5958; // @[ICache.scala 169:30]
  wire  _GEN_7512 = uncached ? _GEN_1173 : _GEN_5959; // @[ICache.scala 169:30]
  wire  _GEN_7513 = uncached ? _GEN_1685 : _GEN_5960; // @[ICache.scala 169:30]
  wire  _GEN_7514 = uncached ? _GEN_1174 : _GEN_5961; // @[ICache.scala 169:30]
  wire  _GEN_7515 = uncached ? _GEN_1686 : _GEN_5962; // @[ICache.scala 169:30]
  wire  _GEN_7516 = uncached ? _GEN_1175 : _GEN_5963; // @[ICache.scala 169:30]
  wire  _GEN_7517 = uncached ? _GEN_1687 : _GEN_5964; // @[ICache.scala 169:30]
  wire  _GEN_7518 = uncached ? _GEN_1176 : _GEN_5965; // @[ICache.scala 169:30]
  wire  _GEN_7519 = uncached ? _GEN_1688 : _GEN_5966; // @[ICache.scala 169:30]
  wire  _GEN_7520 = uncached ? _GEN_1177 : _GEN_5967; // @[ICache.scala 169:30]
  wire  _GEN_7521 = uncached ? _GEN_1689 : _GEN_5968; // @[ICache.scala 169:30]
  wire  _GEN_7522 = uncached ? _GEN_1178 : _GEN_5969; // @[ICache.scala 169:30]
  wire  _GEN_7523 = uncached ? _GEN_1690 : _GEN_5970; // @[ICache.scala 169:30]
  wire  _GEN_7524 = uncached ? _GEN_1179 : _GEN_5971; // @[ICache.scala 169:30]
  wire  _GEN_7525 = uncached ? _GEN_1691 : _GEN_5972; // @[ICache.scala 169:30]
  wire  _GEN_7526 = uncached ? _GEN_1180 : _GEN_5973; // @[ICache.scala 169:30]
  wire  _GEN_7527 = uncached ? _GEN_1692 : _GEN_5974; // @[ICache.scala 169:30]
  wire  _GEN_7528 = uncached ? _GEN_1181 : _GEN_5975; // @[ICache.scala 169:30]
  wire  _GEN_7529 = uncached ? _GEN_1693 : _GEN_5976; // @[ICache.scala 169:30]
  wire  _GEN_7530 = uncached ? _GEN_1182 : _GEN_5977; // @[ICache.scala 169:30]
  wire  _GEN_7531 = uncached ? _GEN_1694 : _GEN_5978; // @[ICache.scala 169:30]
  wire  _GEN_7532 = uncached ? _GEN_1183 : _GEN_5979; // @[ICache.scala 169:30]
  wire  _GEN_7533 = uncached ? _GEN_1695 : _GEN_5980; // @[ICache.scala 169:30]
  wire  _GEN_7534 = uncached ? _GEN_1184 : _GEN_5981; // @[ICache.scala 169:30]
  wire  _GEN_7535 = uncached ? _GEN_1696 : _GEN_5982; // @[ICache.scala 169:30]
  wire  _GEN_7536 = uncached ? _GEN_1185 : _GEN_5983; // @[ICache.scala 169:30]
  wire  _GEN_7537 = uncached ? _GEN_1697 : _GEN_5984; // @[ICache.scala 169:30]
  wire  _GEN_7538 = uncached ? _GEN_1186 : _GEN_5985; // @[ICache.scala 169:30]
  wire  _GEN_7539 = uncached ? _GEN_1698 : _GEN_5986; // @[ICache.scala 169:30]
  wire  _GEN_7540 = uncached ? _GEN_1187 : _GEN_5987; // @[ICache.scala 169:30]
  wire  _GEN_7541 = uncached ? _GEN_1699 : _GEN_5988; // @[ICache.scala 169:30]
  wire  _GEN_7542 = uncached ? _GEN_1188 : _GEN_5989; // @[ICache.scala 169:30]
  wire  _GEN_7543 = uncached ? _GEN_1700 : _GEN_5990; // @[ICache.scala 169:30]
  wire  _GEN_7544 = uncached ? _GEN_1189 : _GEN_5991; // @[ICache.scala 169:30]
  wire  _GEN_7545 = uncached ? _GEN_1701 : _GEN_5992; // @[ICache.scala 169:30]
  wire  _GEN_7546 = uncached ? _GEN_1190 : _GEN_5993; // @[ICache.scala 169:30]
  wire  _GEN_7547 = uncached ? _GEN_1702 : _GEN_5994; // @[ICache.scala 169:30]
  wire  _GEN_7548 = uncached ? _GEN_1191 : _GEN_5995; // @[ICache.scala 169:30]
  wire  _GEN_7549 = uncached ? _GEN_1703 : _GEN_5996; // @[ICache.scala 169:30]
  wire  _GEN_7550 = uncached ? _GEN_1192 : _GEN_5997; // @[ICache.scala 169:30]
  wire  _GEN_7551 = uncached ? _GEN_1704 : _GEN_5998; // @[ICache.scala 169:30]
  wire  _GEN_7552 = uncached ? _GEN_1193 : _GEN_5999; // @[ICache.scala 169:30]
  wire  _GEN_7553 = uncached ? _GEN_1705 : _GEN_6000; // @[ICache.scala 169:30]
  wire  _GEN_7554 = uncached ? _GEN_1194 : _GEN_6001; // @[ICache.scala 169:30]
  wire  _GEN_7555 = uncached ? _GEN_1706 : _GEN_6002; // @[ICache.scala 169:30]
  wire  _GEN_7556 = uncached ? _GEN_1195 : _GEN_6003; // @[ICache.scala 169:30]
  wire  _GEN_7557 = uncached ? _GEN_1707 : _GEN_6004; // @[ICache.scala 169:30]
  wire  _GEN_7558 = uncached ? _GEN_1196 : _GEN_6005; // @[ICache.scala 169:30]
  wire  _GEN_7559 = uncached ? _GEN_1708 : _GEN_6006; // @[ICache.scala 169:30]
  wire  _GEN_7560 = uncached ? _GEN_1197 : _GEN_6007; // @[ICache.scala 169:30]
  wire  _GEN_7561 = uncached ? _GEN_1709 : _GEN_6008; // @[ICache.scala 169:30]
  wire  _GEN_7562 = uncached ? _GEN_1198 : _GEN_6009; // @[ICache.scala 169:30]
  wire  _GEN_7563 = uncached ? _GEN_1710 : _GEN_6010; // @[ICache.scala 169:30]
  wire  _GEN_7564 = uncached ? _GEN_1199 : _GEN_6011; // @[ICache.scala 169:30]
  wire  _GEN_7565 = uncached ? _GEN_1711 : _GEN_6012; // @[ICache.scala 169:30]
  wire  _GEN_7566 = uncached ? _GEN_1200 : _GEN_6013; // @[ICache.scala 169:30]
  wire  _GEN_7567 = uncached ? _GEN_1712 : _GEN_6014; // @[ICache.scala 169:30]
  wire  _GEN_7568 = uncached ? _GEN_1201 : _GEN_6015; // @[ICache.scala 169:30]
  wire  _GEN_7569 = uncached ? _GEN_1713 : _GEN_6016; // @[ICache.scala 169:30]
  wire  _GEN_7570 = uncached ? _GEN_1202 : _GEN_6017; // @[ICache.scala 169:30]
  wire  _GEN_7571 = uncached ? _GEN_1714 : _GEN_6018; // @[ICache.scala 169:30]
  wire  _GEN_7572 = uncached ? _GEN_1203 : _GEN_6019; // @[ICache.scala 169:30]
  wire  _GEN_7573 = uncached ? _GEN_1715 : _GEN_6020; // @[ICache.scala 169:30]
  wire  _GEN_7574 = uncached ? _GEN_1204 : _GEN_6021; // @[ICache.scala 169:30]
  wire  _GEN_7575 = uncached ? _GEN_1716 : _GEN_6022; // @[ICache.scala 169:30]
  wire  _GEN_7576 = uncached ? _GEN_1205 : _GEN_6023; // @[ICache.scala 169:30]
  wire  _GEN_7577 = uncached ? _GEN_1717 : _GEN_6024; // @[ICache.scala 169:30]
  wire  _GEN_7578 = uncached ? _GEN_1206 : _GEN_6025; // @[ICache.scala 169:30]
  wire  _GEN_7579 = uncached ? _GEN_1718 : _GEN_6026; // @[ICache.scala 169:30]
  wire  _GEN_7580 = uncached ? _GEN_1207 : _GEN_6027; // @[ICache.scala 169:30]
  wire  _GEN_7581 = uncached ? _GEN_1719 : _GEN_6028; // @[ICache.scala 169:30]
  wire  _GEN_7582 = uncached ? _GEN_1208 : _GEN_6029; // @[ICache.scala 169:30]
  wire  _GEN_7583 = uncached ? _GEN_1720 : _GEN_6030; // @[ICache.scala 169:30]
  wire  _GEN_7584 = uncached ? _GEN_1209 : _GEN_6031; // @[ICache.scala 169:30]
  wire  _GEN_7585 = uncached ? _GEN_1721 : _GEN_6032; // @[ICache.scala 169:30]
  wire  _GEN_7586 = uncached ? _GEN_1210 : _GEN_6033; // @[ICache.scala 169:30]
  wire  _GEN_7587 = uncached ? _GEN_1722 : _GEN_6034; // @[ICache.scala 169:30]
  wire  _GEN_7588 = uncached ? _GEN_1211 : _GEN_6035; // @[ICache.scala 169:30]
  wire  _GEN_7589 = uncached ? _GEN_1723 : _GEN_6036; // @[ICache.scala 169:30]
  wire  _GEN_7590 = uncached ? _GEN_1212 : _GEN_6037; // @[ICache.scala 169:30]
  wire  _GEN_7591 = uncached ? _GEN_1724 : _GEN_6038; // @[ICache.scala 169:30]
  wire  _GEN_7592 = uncached ? _GEN_1213 : _GEN_6039; // @[ICache.scala 169:30]
  wire  _GEN_7593 = uncached ? _GEN_1725 : _GEN_6040; // @[ICache.scala 169:30]
  wire  _GEN_7594 = uncached ? _GEN_1214 : _GEN_6041; // @[ICache.scala 169:30]
  wire  _GEN_7595 = uncached ? _GEN_1726 : _GEN_6042; // @[ICache.scala 169:30]
  wire  _GEN_7596 = uncached ? _GEN_1215 : _GEN_6043; // @[ICache.scala 169:30]
  wire  _GEN_7597 = uncached ? _GEN_1727 : _GEN_6044; // @[ICache.scala 169:30]
  wire  _GEN_7598 = uncached ? _GEN_1216 : _GEN_6045; // @[ICache.scala 169:30]
  wire  _GEN_7599 = uncached ? _GEN_1728 : _GEN_6046; // @[ICache.scala 169:30]
  wire  _GEN_7600 = uncached ? _GEN_1217 : _GEN_6047; // @[ICache.scala 169:30]
  wire  _GEN_7601 = uncached ? _GEN_1729 : _GEN_6048; // @[ICache.scala 169:30]
  wire  _GEN_7602 = uncached ? _GEN_1218 : _GEN_6049; // @[ICache.scala 169:30]
  wire  _GEN_7603 = uncached ? _GEN_1730 : _GEN_6050; // @[ICache.scala 169:30]
  wire  _GEN_7604 = uncached ? _GEN_1219 : _GEN_6051; // @[ICache.scala 169:30]
  wire  _GEN_7605 = uncached ? _GEN_1731 : _GEN_6052; // @[ICache.scala 169:30]
  wire  _GEN_7606 = uncached ? _GEN_1220 : _GEN_6053; // @[ICache.scala 169:30]
  wire  _GEN_7607 = uncached ? _GEN_1732 : _GEN_6054; // @[ICache.scala 169:30]
  wire  _GEN_7608 = uncached ? _GEN_1221 : _GEN_6055; // @[ICache.scala 169:30]
  wire  _GEN_7609 = uncached ? _GEN_1733 : _GEN_6056; // @[ICache.scala 169:30]
  wire  _GEN_7610 = uncached ? _GEN_1222 : _GEN_6057; // @[ICache.scala 169:30]
  wire  _GEN_7611 = uncached ? _GEN_1734 : _GEN_6058; // @[ICache.scala 169:30]
  wire  _GEN_7612 = uncached ? _GEN_1223 : _GEN_6059; // @[ICache.scala 169:30]
  wire  _GEN_7613 = uncached ? _GEN_1735 : _GEN_6060; // @[ICache.scala 169:30]
  wire  _GEN_7614 = uncached ? _GEN_1224 : _GEN_6061; // @[ICache.scala 169:30]
  wire  _GEN_7615 = uncached ? _GEN_1736 : _GEN_6062; // @[ICache.scala 169:30]
  wire  _GEN_7616 = uncached ? _GEN_1225 : _GEN_6063; // @[ICache.scala 169:30]
  wire  _GEN_7617 = uncached ? _GEN_1737 : _GEN_6064; // @[ICache.scala 169:30]
  wire  _GEN_7618 = uncached ? _GEN_1226 : _GEN_6065; // @[ICache.scala 169:30]
  wire  _GEN_7619 = uncached ? _GEN_1738 : _GEN_6066; // @[ICache.scala 169:30]
  wire  _GEN_7620 = uncached ? _GEN_1227 : _GEN_6067; // @[ICache.scala 169:30]
  wire  _GEN_7621 = uncached ? _GEN_1739 : _GEN_6068; // @[ICache.scala 169:30]
  wire  _GEN_7622 = uncached ? _GEN_1228 : _GEN_6069; // @[ICache.scala 169:30]
  wire  _GEN_7623 = uncached ? _GEN_1740 : _GEN_6070; // @[ICache.scala 169:30]
  wire  _GEN_7624 = uncached ? _GEN_1229 : _GEN_6071; // @[ICache.scala 169:30]
  wire  _GEN_7625 = uncached ? _GEN_1741 : _GEN_6072; // @[ICache.scala 169:30]
  wire  _GEN_7626 = uncached ? _GEN_1230 : _GEN_6073; // @[ICache.scala 169:30]
  wire  _GEN_7627 = uncached ? _GEN_1742 : _GEN_6074; // @[ICache.scala 169:30]
  wire  _GEN_7628 = uncached ? _GEN_1231 : _GEN_6075; // @[ICache.scala 169:30]
  wire  _GEN_7629 = uncached ? _GEN_1743 : _GEN_6076; // @[ICache.scala 169:30]
  wire  _GEN_7630 = uncached ? _GEN_1232 : _GEN_6077; // @[ICache.scala 169:30]
  wire  _GEN_7631 = uncached ? _GEN_1744 : _GEN_6078; // @[ICache.scala 169:30]
  wire  _GEN_7632 = uncached ? _GEN_1233 : _GEN_6079; // @[ICache.scala 169:30]
  wire  _GEN_7633 = uncached ? _GEN_1745 : _GEN_6080; // @[ICache.scala 169:30]
  wire  _GEN_7634 = uncached ? _GEN_1234 : _GEN_6081; // @[ICache.scala 169:30]
  wire  _GEN_7635 = uncached ? _GEN_1746 : _GEN_6082; // @[ICache.scala 169:30]
  wire  _GEN_7636 = uncached ? _GEN_1235 : _GEN_6083; // @[ICache.scala 169:30]
  wire  _GEN_7637 = uncached ? _GEN_1747 : _GEN_6084; // @[ICache.scala 169:30]
  wire  _GEN_7638 = uncached ? _GEN_1236 : _GEN_6085; // @[ICache.scala 169:30]
  wire  _GEN_7639 = uncached ? _GEN_1748 : _GEN_6086; // @[ICache.scala 169:30]
  wire  _GEN_7640 = uncached ? _GEN_1237 : _GEN_6087; // @[ICache.scala 169:30]
  wire  _GEN_7641 = uncached ? _GEN_1749 : _GEN_6088; // @[ICache.scala 169:30]
  wire  _GEN_7642 = uncached ? _GEN_1238 : _GEN_6089; // @[ICache.scala 169:30]
  wire  _GEN_7643 = uncached ? _GEN_1750 : _GEN_6090; // @[ICache.scala 169:30]
  wire  _GEN_7644 = uncached ? _GEN_1239 : _GEN_6091; // @[ICache.scala 169:30]
  wire  _GEN_7645 = uncached ? _GEN_1751 : _GEN_6092; // @[ICache.scala 169:30]
  wire  _GEN_7646 = uncached ? _GEN_1240 : _GEN_6093; // @[ICache.scala 169:30]
  wire  _GEN_7647 = uncached ? _GEN_1752 : _GEN_6094; // @[ICache.scala 169:30]
  wire  _GEN_7648 = uncached ? _GEN_1241 : _GEN_6095; // @[ICache.scala 169:30]
  wire  _GEN_7649 = uncached ? _GEN_1753 : _GEN_6096; // @[ICache.scala 169:30]
  wire  _GEN_7650 = uncached ? _GEN_1242 : _GEN_6097; // @[ICache.scala 169:30]
  wire  _GEN_7651 = uncached ? _GEN_1754 : _GEN_6098; // @[ICache.scala 169:30]
  wire  _GEN_7652 = uncached ? _GEN_1243 : _GEN_6099; // @[ICache.scala 169:30]
  wire  _GEN_7653 = uncached ? _GEN_1755 : _GEN_6100; // @[ICache.scala 169:30]
  wire  _GEN_7654 = uncached ? _GEN_1244 : _GEN_6101; // @[ICache.scala 169:30]
  wire  _GEN_7655 = uncached ? _GEN_1756 : _GEN_6102; // @[ICache.scala 169:30]
  wire  _GEN_7656 = uncached ? _GEN_1245 : _GEN_6103; // @[ICache.scala 169:30]
  wire  _GEN_7657 = uncached ? _GEN_1757 : _GEN_6104; // @[ICache.scala 169:30]
  wire  _GEN_7658 = uncached ? _GEN_1246 : _GEN_6105; // @[ICache.scala 169:30]
  wire  _GEN_7659 = uncached ? _GEN_1758 : _GEN_6106; // @[ICache.scala 169:30]
  wire  _GEN_7660 = uncached ? _GEN_1247 : _GEN_6107; // @[ICache.scala 169:30]
  wire  _GEN_7661 = uncached ? _GEN_1759 : _GEN_6108; // @[ICache.scala 169:30]
  wire  _GEN_7662 = uncached ? _GEN_1248 : _GEN_6109; // @[ICache.scala 169:30]
  wire  _GEN_7663 = uncached ? _GEN_1760 : _GEN_6110; // @[ICache.scala 169:30]
  wire  _GEN_7664 = uncached ? _GEN_1249 : _GEN_6111; // @[ICache.scala 169:30]
  wire  _GEN_7665 = uncached ? _GEN_1761 : _GEN_6112; // @[ICache.scala 169:30]
  wire  _GEN_7666 = uncached ? _GEN_1250 : _GEN_6113; // @[ICache.scala 169:30]
  wire  _GEN_7667 = uncached ? _GEN_1762 : _GEN_6114; // @[ICache.scala 169:30]
  wire  _GEN_7668 = uncached ? _GEN_1251 : _GEN_6115; // @[ICache.scala 169:30]
  wire  _GEN_7669 = uncached ? _GEN_1763 : _GEN_6116; // @[ICache.scala 169:30]
  wire  _GEN_7670 = uncached ? _GEN_1252 : _GEN_6117; // @[ICache.scala 169:30]
  wire  _GEN_7671 = uncached ? _GEN_1764 : _GEN_6118; // @[ICache.scala 169:30]
  wire  _GEN_7672 = uncached ? _GEN_1253 : _GEN_6119; // @[ICache.scala 169:30]
  wire  _GEN_7673 = uncached ? _GEN_1765 : _GEN_6120; // @[ICache.scala 169:30]
  wire  _GEN_7674 = uncached ? _GEN_1254 : _GEN_6121; // @[ICache.scala 169:30]
  wire  _GEN_7675 = uncached ? _GEN_1766 : _GEN_6122; // @[ICache.scala 169:30]
  wire  _GEN_7676 = uncached ? _GEN_1255 : _GEN_6123; // @[ICache.scala 169:30]
  wire  _GEN_7677 = uncached ? _GEN_1767 : _GEN_6124; // @[ICache.scala 169:30]
  wire  _GEN_7678 = uncached ? _GEN_1256 : _GEN_6125; // @[ICache.scala 169:30]
  wire  _GEN_7679 = uncached ? _GEN_1768 : _GEN_6126; // @[ICache.scala 169:30]
  wire  _GEN_7680 = uncached ? _GEN_1257 : _GEN_6127; // @[ICache.scala 169:30]
  wire  _GEN_7681 = uncached ? _GEN_1769 : _GEN_6128; // @[ICache.scala 169:30]
  wire  _GEN_7682 = uncached ? _GEN_1258 : _GEN_6129; // @[ICache.scala 169:30]
  wire  _GEN_7683 = uncached ? _GEN_1770 : _GEN_6130; // @[ICache.scala 169:30]
  wire  _GEN_7684 = uncached ? _GEN_1259 : _GEN_6131; // @[ICache.scala 169:30]
  wire  _GEN_7685 = uncached ? _GEN_1771 : _GEN_6132; // @[ICache.scala 169:30]
  wire  _GEN_7686 = uncached ? _GEN_1260 : _GEN_6133; // @[ICache.scala 169:30]
  wire  _GEN_7687 = uncached ? _GEN_1772 : _GEN_6134; // @[ICache.scala 169:30]
  wire  _GEN_7688 = uncached ? _GEN_1261 : _GEN_6135; // @[ICache.scala 169:30]
  wire  _GEN_7689 = uncached ? _GEN_1773 : _GEN_6136; // @[ICache.scala 169:30]
  wire  _GEN_7690 = uncached ? _GEN_1262 : _GEN_6137; // @[ICache.scala 169:30]
  wire  _GEN_7691 = uncached ? _GEN_1774 : _GEN_6138; // @[ICache.scala 169:30]
  wire  _GEN_7692 = uncached ? _GEN_1263 : _GEN_6139; // @[ICache.scala 169:30]
  wire  _GEN_7693 = uncached ? _GEN_1775 : _GEN_6140; // @[ICache.scala 169:30]
  wire  _GEN_7694 = uncached ? _GEN_1264 : _GEN_6141; // @[ICache.scala 169:30]
  wire  _GEN_7695 = uncached ? _GEN_1776 : _GEN_6142; // @[ICache.scala 169:30]
  wire  _GEN_7696 = uncached ? _GEN_1265 : _GEN_6143; // @[ICache.scala 169:30]
  wire  _GEN_7697 = uncached ? _GEN_1777 : _GEN_6144; // @[ICache.scala 169:30]
  wire  _GEN_7698 = uncached ? _GEN_1266 : _GEN_6145; // @[ICache.scala 169:30]
  wire  _GEN_7699 = uncached ? _GEN_1778 : _GEN_6146; // @[ICache.scala 169:30]
  wire  _GEN_7700 = uncached ? _GEN_1267 : _GEN_6147; // @[ICache.scala 169:30]
  wire  _GEN_7701 = uncached ? _GEN_1779 : _GEN_6148; // @[ICache.scala 169:30]
  wire  _GEN_7702 = uncached ? _GEN_1268 : _GEN_6149; // @[ICache.scala 169:30]
  wire  _GEN_7703 = uncached ? _GEN_1780 : _GEN_6150; // @[ICache.scala 169:30]
  wire  _GEN_7704 = uncached ? _GEN_1269 : _GEN_6151; // @[ICache.scala 169:30]
  wire  _GEN_7705 = uncached ? _GEN_1781 : _GEN_6152; // @[ICache.scala 169:30]
  wire  _GEN_7706 = uncached ? _GEN_1270 : _GEN_6153; // @[ICache.scala 169:30]
  wire  _GEN_7707 = uncached ? _GEN_1782 : _GEN_6154; // @[ICache.scala 169:30]
  wire  _GEN_7708 = uncached ? _GEN_1271 : _GEN_6155; // @[ICache.scala 169:30]
  wire  _GEN_7709 = uncached ? _GEN_1783 : _GEN_6156; // @[ICache.scala 169:30]
  wire  _GEN_7710 = uncached ? _GEN_1272 : _GEN_6157; // @[ICache.scala 169:30]
  wire  _GEN_7711 = uncached ? _GEN_1784 : _GEN_6158; // @[ICache.scala 169:30]
  wire  _GEN_7712 = uncached ? _GEN_1273 : _GEN_6159; // @[ICache.scala 169:30]
  wire  _GEN_7713 = uncached ? _GEN_1785 : _GEN_6160; // @[ICache.scala 169:30]
  wire  _GEN_7714 = uncached ? _GEN_1274 : _GEN_6161; // @[ICache.scala 169:30]
  wire  _GEN_7715 = uncached ? _GEN_1786 : _GEN_6162; // @[ICache.scala 169:30]
  wire  _GEN_7716 = uncached ? _GEN_1275 : _GEN_6163; // @[ICache.scala 169:30]
  wire  _GEN_7717 = uncached ? _GEN_1787 : _GEN_6164; // @[ICache.scala 169:30]
  wire  _GEN_7718 = uncached ? _GEN_1276 : _GEN_6165; // @[ICache.scala 169:30]
  wire  _GEN_7719 = uncached ? _GEN_1788 : _GEN_6166; // @[ICache.scala 169:30]
  wire  _GEN_7720 = uncached ? _GEN_1277 : _GEN_6167; // @[ICache.scala 169:30]
  wire  _GEN_7721 = uncached ? _GEN_1789 : _GEN_6168; // @[ICache.scala 169:30]
  wire  _GEN_7722 = uncached ? _GEN_1278 : _GEN_6169; // @[ICache.scala 169:30]
  wire  _GEN_7723 = uncached ? _GEN_1790 : _GEN_6170; // @[ICache.scala 169:30]
  wire  _GEN_7724 = uncached ? _GEN_1279 : _GEN_6171; // @[ICache.scala 169:30]
  wire  _GEN_7725 = uncached ? _GEN_1791 : _GEN_6172; // @[ICache.scala 169:30]
  wire  _GEN_7726 = uncached ? _GEN_1280 : _GEN_6173; // @[ICache.scala 169:30]
  wire  _GEN_7727 = uncached ? _GEN_1792 : _GEN_6174; // @[ICache.scala 169:30]
  wire  _GEN_7728 = uncached ? _GEN_1281 : _GEN_6175; // @[ICache.scala 169:30]
  wire  _GEN_7729 = uncached ? _GEN_1793 : _GEN_6176; // @[ICache.scala 169:30]
  wire  _GEN_7730 = uncached ? _GEN_1282 : _GEN_6177; // @[ICache.scala 169:30]
  wire  _GEN_7731 = uncached ? _GEN_1794 : _GEN_6178; // @[ICache.scala 169:30]
  wire  _GEN_7732 = uncached ? _GEN_1283 : _GEN_6179; // @[ICache.scala 169:30]
  wire  _GEN_7733 = uncached ? _GEN_1795 : _GEN_6180; // @[ICache.scala 169:30]
  wire  _GEN_7734 = uncached ? _GEN_1284 : _GEN_6181; // @[ICache.scala 169:30]
  wire  _GEN_7735 = uncached ? _GEN_1796 : _GEN_6182; // @[ICache.scala 169:30]
  wire  _GEN_7736 = uncached ? _GEN_1285 : _GEN_6183; // @[ICache.scala 169:30]
  wire  _GEN_7737 = uncached ? _GEN_1797 : _GEN_6184; // @[ICache.scala 169:30]
  wire  _GEN_7738 = uncached ? _GEN_1286 : _GEN_6185; // @[ICache.scala 169:30]
  wire  _GEN_7739 = uncached ? _GEN_1798 : _GEN_6186; // @[ICache.scala 169:30]
  wire  _GEN_7740 = uncached ? _GEN_1287 : _GEN_6187; // @[ICache.scala 169:30]
  wire  _GEN_7741 = uncached ? _GEN_1799 : _GEN_6188; // @[ICache.scala 169:30]
  wire  _GEN_7742 = uncached ? _GEN_1288 : _GEN_6189; // @[ICache.scala 169:30]
  wire  _GEN_7743 = uncached ? _GEN_1800 : _GEN_6190; // @[ICache.scala 169:30]
  wire  _GEN_7744 = uncached ? _GEN_1289 : _GEN_6191; // @[ICache.scala 169:30]
  wire  _GEN_7745 = uncached ? _GEN_1801 : _GEN_6192; // @[ICache.scala 169:30]
  wire  _GEN_7746 = uncached ? _GEN_1290 : _GEN_6193; // @[ICache.scala 169:30]
  wire  _GEN_7747 = uncached ? _GEN_1802 : _GEN_6194; // @[ICache.scala 169:30]
  wire  _GEN_7748 = uncached ? _GEN_1291 : _GEN_6195; // @[ICache.scala 169:30]
  wire  _GEN_7749 = uncached ? _GEN_1803 : _GEN_6196; // @[ICache.scala 169:30]
  wire  _GEN_7750 = uncached ? _GEN_1292 : _GEN_6197; // @[ICache.scala 169:30]
  wire  _GEN_7751 = uncached ? _GEN_1804 : _GEN_6198; // @[ICache.scala 169:30]
  wire  _GEN_7752 = uncached ? _GEN_1293 : _GEN_6199; // @[ICache.scala 169:30]
  wire  _GEN_7753 = uncached ? _GEN_1805 : _GEN_6200; // @[ICache.scala 169:30]
  wire  _GEN_7754 = uncached ? _GEN_1294 : _GEN_6201; // @[ICache.scala 169:30]
  wire  _GEN_7755 = uncached ? _GEN_1806 : _GEN_6202; // @[ICache.scala 169:30]
  wire  _GEN_7756 = uncached ? _GEN_1295 : _GEN_6203; // @[ICache.scala 169:30]
  wire  _GEN_7757 = uncached ? _GEN_1807 : _GEN_6204; // @[ICache.scala 169:30]
  wire  _GEN_7758 = uncached ? _GEN_1296 : _GEN_6205; // @[ICache.scala 169:30]
  wire  _GEN_7759 = uncached ? _GEN_1808 : _GEN_6206; // @[ICache.scala 169:30]
  wire  _GEN_7760 = uncached ? _GEN_1297 : _GEN_6207; // @[ICache.scala 169:30]
  wire  _GEN_7761 = uncached ? _GEN_1809 : _GEN_6208; // @[ICache.scala 169:30]
  wire  _GEN_7762 = uncached ? _GEN_1298 : _GEN_6209; // @[ICache.scala 169:30]
  wire  _GEN_7763 = uncached ? _GEN_1810 : _GEN_6210; // @[ICache.scala 169:30]
  wire  _GEN_7764 = uncached ? _GEN_1299 : _GEN_6211; // @[ICache.scala 169:30]
  wire  _GEN_7765 = uncached ? _GEN_1811 : _GEN_6212; // @[ICache.scala 169:30]
  wire  _GEN_7766 = uncached ? _GEN_1300 : _GEN_6213; // @[ICache.scala 169:30]
  wire  _GEN_7767 = uncached ? _GEN_1812 : _GEN_6214; // @[ICache.scala 169:30]
  wire  _GEN_7768 = uncached ? _GEN_1301 : _GEN_6215; // @[ICache.scala 169:30]
  wire  _GEN_7769 = uncached ? _GEN_1813 : _GEN_6216; // @[ICache.scala 169:30]
  wire  _GEN_7770 = uncached ? _GEN_1302 : _GEN_6217; // @[ICache.scala 169:30]
  wire  _GEN_7771 = uncached ? _GEN_1814 : _GEN_6218; // @[ICache.scala 169:30]
  wire  _GEN_7772 = uncached ? _GEN_1303 : _GEN_6219; // @[ICache.scala 169:30]
  wire  _GEN_7773 = uncached ? _GEN_1815 : _GEN_6220; // @[ICache.scala 169:30]
  wire  _GEN_7774 = uncached ? _GEN_1304 : _GEN_6221; // @[ICache.scala 169:30]
  wire  _GEN_7775 = uncached ? _GEN_1816 : _GEN_6222; // @[ICache.scala 169:30]
  wire  _GEN_7776 = uncached ? _GEN_1305 : _GEN_6223; // @[ICache.scala 169:30]
  wire  _GEN_7777 = uncached ? _GEN_1817 : _GEN_6224; // @[ICache.scala 169:30]
  wire  _GEN_7778 = uncached ? _GEN_1306 : _GEN_6225; // @[ICache.scala 169:30]
  wire  _GEN_7779 = uncached ? _GEN_1818 : _GEN_6226; // @[ICache.scala 169:30]
  wire  _GEN_7780 = uncached ? _GEN_1307 : _GEN_6227; // @[ICache.scala 169:30]
  wire  _GEN_7781 = uncached ? _GEN_1819 : _GEN_6228; // @[ICache.scala 169:30]
  wire  _GEN_7782 = uncached ? _GEN_1308 : _GEN_6229; // @[ICache.scala 169:30]
  wire  _GEN_7783 = uncached ? _GEN_1820 : _GEN_6230; // @[ICache.scala 169:30]
  wire  _GEN_7784 = uncached ? _GEN_1309 : _GEN_6231; // @[ICache.scala 169:30]
  wire  _GEN_7785 = uncached ? _GEN_1821 : _GEN_6232; // @[ICache.scala 169:30]
  wire  _GEN_7786 = uncached ? _GEN_1310 : _GEN_6233; // @[ICache.scala 169:30]
  wire  _GEN_7787 = uncached ? _GEN_1822 : _GEN_6234; // @[ICache.scala 169:30]
  wire  _GEN_7788 = uncached ? _GEN_1311 : _GEN_6235; // @[ICache.scala 169:30]
  wire  _GEN_7789 = uncached ? _GEN_1823 : _GEN_6236; // @[ICache.scala 169:30]
  wire  _GEN_7790 = uncached ? _GEN_1312 : _GEN_6237; // @[ICache.scala 169:30]
  wire  _GEN_7791 = uncached ? _GEN_1824 : _GEN_6238; // @[ICache.scala 169:30]
  wire  _GEN_7792 = uncached ? _GEN_1313 : _GEN_6239; // @[ICache.scala 169:30]
  wire  _GEN_7793 = uncached ? _GEN_1825 : _GEN_6240; // @[ICache.scala 169:30]
  wire  _GEN_7794 = uncached ? _GEN_1314 : _GEN_6241; // @[ICache.scala 169:30]
  wire  _GEN_7795 = uncached ? _GEN_1826 : _GEN_6242; // @[ICache.scala 169:30]
  wire  _GEN_7796 = uncached ? _GEN_1315 : _GEN_6243; // @[ICache.scala 169:30]
  wire  _GEN_7797 = uncached ? _GEN_1827 : _GEN_6244; // @[ICache.scala 169:30]
  wire  _GEN_7798 = uncached ? _GEN_1316 : _GEN_6245; // @[ICache.scala 169:30]
  wire  _GEN_7799 = uncached ? _GEN_1828 : _GEN_6246; // @[ICache.scala 169:30]
  wire  _GEN_7800 = uncached ? _GEN_1317 : _GEN_6247; // @[ICache.scala 169:30]
  wire  _GEN_7801 = uncached ? _GEN_1829 : _GEN_6248; // @[ICache.scala 169:30]
  wire  _GEN_7802 = uncached ? _GEN_1318 : _GEN_6249; // @[ICache.scala 169:30]
  wire  _GEN_7803 = uncached ? _GEN_1830 : _GEN_6250; // @[ICache.scala 169:30]
  wire  _GEN_7804 = uncached ? _GEN_1319 : _GEN_6251; // @[ICache.scala 169:30]
  wire  _GEN_7805 = uncached ? _GEN_1831 : _GEN_6252; // @[ICache.scala 169:30]
  wire  _GEN_7806 = uncached ? _GEN_1320 : _GEN_6253; // @[ICache.scala 169:30]
  wire  _GEN_7807 = uncached ? _GEN_1832 : _GEN_6254; // @[ICache.scala 169:30]
  wire  _GEN_7808 = uncached ? _GEN_1321 : _GEN_6255; // @[ICache.scala 169:30]
  wire  _GEN_7809 = uncached ? _GEN_1833 : _GEN_6256; // @[ICache.scala 169:30]
  wire  _GEN_7810 = uncached ? _GEN_1322 : _GEN_6257; // @[ICache.scala 169:30]
  wire  _GEN_7811 = uncached ? _GEN_1834 : _GEN_6258; // @[ICache.scala 169:30]
  wire  _GEN_7812 = uncached ? _GEN_1323 : _GEN_6259; // @[ICache.scala 169:30]
  wire  _GEN_7813 = uncached ? _GEN_1835 : _GEN_6260; // @[ICache.scala 169:30]
  wire  _GEN_7814 = uncached ? _GEN_1324 : _GEN_6261; // @[ICache.scala 169:30]
  wire  _GEN_7815 = uncached ? _GEN_1836 : _GEN_6262; // @[ICache.scala 169:30]
  wire  _GEN_7816 = uncached ? _GEN_1325 : _GEN_6263; // @[ICache.scala 169:30]
  wire  _GEN_7817 = uncached ? _GEN_1837 : _GEN_6264; // @[ICache.scala 169:30]
  wire  _GEN_7818 = uncached ? _GEN_1326 : _GEN_6265; // @[ICache.scala 169:30]
  wire  _GEN_7819 = uncached ? _GEN_1838 : _GEN_6266; // @[ICache.scala 169:30]
  wire  _GEN_7820 = uncached ? _GEN_1327 : _GEN_6267; // @[ICache.scala 169:30]
  wire  _GEN_7821 = uncached ? _GEN_1839 : _GEN_6268; // @[ICache.scala 169:30]
  wire  _GEN_7822 = uncached ? _GEN_1328 : _GEN_6269; // @[ICache.scala 169:30]
  wire  _GEN_7823 = uncached ? _GEN_1840 : _GEN_6270; // @[ICache.scala 169:30]
  wire  _GEN_7824 = uncached ? _GEN_1329 : _GEN_6271; // @[ICache.scala 169:30]
  wire  _GEN_7825 = uncached ? _GEN_1841 : _GEN_6272; // @[ICache.scala 169:30]
  wire  _GEN_7826 = uncached ? _GEN_1330 : _GEN_6273; // @[ICache.scala 169:30]
  wire  _GEN_7827 = uncached ? _GEN_1842 : _GEN_6274; // @[ICache.scala 169:30]
  wire  _GEN_7828 = uncached ? _GEN_1331 : _GEN_6275; // @[ICache.scala 169:30]
  wire  _GEN_7829 = uncached ? _GEN_1843 : _GEN_6276; // @[ICache.scala 169:30]
  wire  _GEN_7830 = uncached ? _GEN_1332 : _GEN_6277; // @[ICache.scala 169:30]
  wire  _GEN_7831 = uncached ? _GEN_1844 : _GEN_6278; // @[ICache.scala 169:30]
  wire  _GEN_7832 = uncached ? _GEN_1333 : _GEN_6279; // @[ICache.scala 169:30]
  wire  _GEN_7833 = uncached ? _GEN_1845 : _GEN_6280; // @[ICache.scala 169:30]
  wire  _GEN_7834 = uncached ? _GEN_1334 : _GEN_6281; // @[ICache.scala 169:30]
  wire  _GEN_7835 = uncached ? _GEN_1846 : _GEN_6282; // @[ICache.scala 169:30]
  wire  _GEN_7836 = uncached ? _GEN_1335 : _GEN_6283; // @[ICache.scala 169:30]
  wire  _GEN_7837 = uncached ? _GEN_1847 : _GEN_6284; // @[ICache.scala 169:30]
  wire  _GEN_7838 = uncached ? _GEN_1336 : _GEN_6285; // @[ICache.scala 169:30]
  wire  _GEN_7839 = uncached ? _GEN_1848 : _GEN_6286; // @[ICache.scala 169:30]
  wire  _GEN_7840 = uncached ? _GEN_1337 : _GEN_6287; // @[ICache.scala 169:30]
  wire  _GEN_7841 = uncached ? _GEN_1849 : _GEN_6288; // @[ICache.scala 169:30]
  wire  _GEN_7842 = uncached ? _GEN_1338 : _GEN_6289; // @[ICache.scala 169:30]
  wire  _GEN_7843 = uncached ? _GEN_1850 : _GEN_6290; // @[ICache.scala 169:30]
  wire  _GEN_7844 = uncached ? _GEN_1339 : _GEN_6291; // @[ICache.scala 169:30]
  wire  _GEN_7845 = uncached ? _GEN_1851 : _GEN_6292; // @[ICache.scala 169:30]
  wire  _GEN_7846 = uncached ? _GEN_1340 : _GEN_6293; // @[ICache.scala 169:30]
  wire  _GEN_7847 = uncached ? _GEN_1852 : _GEN_6294; // @[ICache.scala 169:30]
  wire  _GEN_7848 = uncached ? _GEN_1341 : _GEN_6295; // @[ICache.scala 169:30]
  wire  _GEN_7849 = uncached ? _GEN_1853 : _GEN_6296; // @[ICache.scala 169:30]
  wire  _GEN_7850 = uncached ? _GEN_1342 : _GEN_6297; // @[ICache.scala 169:30]
  wire  _GEN_7851 = uncached ? _GEN_1854 : _GEN_6298; // @[ICache.scala 169:30]
  wire  _GEN_7852 = uncached ? _GEN_1343 : _GEN_6299; // @[ICache.scala 169:30]
  wire  _GEN_7853 = uncached ? _GEN_1855 : _GEN_6300; // @[ICache.scala 169:30]
  wire  _GEN_7854 = uncached ? _GEN_1344 : _GEN_6301; // @[ICache.scala 169:30]
  wire  _GEN_7855 = uncached ? _GEN_1856 : _GEN_6302; // @[ICache.scala 169:30]
  wire  _GEN_7856 = uncached ? _GEN_1345 : _GEN_6303; // @[ICache.scala 169:30]
  wire  _GEN_7857 = uncached ? _GEN_1857 : _GEN_6304; // @[ICache.scala 169:30]
  wire  _GEN_7858 = uncached ? _GEN_1346 : _GEN_6305; // @[ICache.scala 169:30]
  wire  _GEN_7859 = uncached ? _GEN_1858 : _GEN_6306; // @[ICache.scala 169:30]
  wire  _GEN_7860 = uncached ? _GEN_1347 : _GEN_6307; // @[ICache.scala 169:30]
  wire  _GEN_7861 = uncached ? _GEN_1859 : _GEN_6308; // @[ICache.scala 169:30]
  wire  _GEN_7862 = uncached ? _GEN_1348 : _GEN_6309; // @[ICache.scala 169:30]
  wire  _GEN_7863 = uncached ? _GEN_1860 : _GEN_6310; // @[ICache.scala 169:30]
  wire  _GEN_7864 = uncached ? _GEN_1349 : _GEN_6311; // @[ICache.scala 169:30]
  wire  _GEN_7865 = uncached ? _GEN_1861 : _GEN_6312; // @[ICache.scala 169:30]
  wire  _GEN_7866 = uncached ? _GEN_1350 : _GEN_6313; // @[ICache.scala 169:30]
  wire  _GEN_7867 = uncached ? _GEN_1862 : _GEN_6314; // @[ICache.scala 169:30]
  wire  _GEN_7868 = uncached ? _GEN_1351 : _GEN_6315; // @[ICache.scala 169:30]
  wire  _GEN_7869 = uncached ? _GEN_1863 : _GEN_6316; // @[ICache.scala 169:30]
  wire  _GEN_7870 = uncached ? _GEN_1352 : _GEN_6317; // @[ICache.scala 169:30]
  wire  _GEN_7871 = uncached ? _GEN_1864 : _GEN_6318; // @[ICache.scala 169:30]
  wire  _GEN_7872 = uncached ? _GEN_1353 : _GEN_6319; // @[ICache.scala 169:30]
  wire  _GEN_7873 = uncached ? _GEN_1865 : _GEN_6320; // @[ICache.scala 169:30]
  wire  _GEN_7874 = uncached ? _GEN_1354 : _GEN_6321; // @[ICache.scala 169:30]
  wire  _GEN_7875 = uncached ? _GEN_1866 : _GEN_6322; // @[ICache.scala 169:30]
  wire  _GEN_7876 = uncached ? _GEN_1355 : _GEN_6323; // @[ICache.scala 169:30]
  wire  _GEN_7877 = uncached ? _GEN_1867 : _GEN_6324; // @[ICache.scala 169:30]
  wire  _GEN_7878 = uncached ? _GEN_1356 : _GEN_6325; // @[ICache.scala 169:30]
  wire  _GEN_7879 = uncached ? _GEN_1868 : _GEN_6326; // @[ICache.scala 169:30]
  wire  _GEN_7880 = uncached ? _GEN_1357 : _GEN_6327; // @[ICache.scala 169:30]
  wire  _GEN_7881 = uncached ? _GEN_1869 : _GEN_6328; // @[ICache.scala 169:30]
  wire  _GEN_7882 = uncached ? _GEN_1358 : _GEN_6329; // @[ICache.scala 169:30]
  wire  _GEN_7883 = uncached ? _GEN_1870 : _GEN_6330; // @[ICache.scala 169:30]
  wire  _GEN_7884 = uncached ? _GEN_1359 : _GEN_6331; // @[ICache.scala 169:30]
  wire  _GEN_7885 = uncached ? _GEN_1871 : _GEN_6332; // @[ICache.scala 169:30]
  wire  _GEN_7886 = uncached ? _GEN_1360 : _GEN_6333; // @[ICache.scala 169:30]
  wire  _GEN_7887 = uncached ? _GEN_1872 : _GEN_6334; // @[ICache.scala 169:30]
  wire  _GEN_7888 = uncached ? _GEN_1361 : _GEN_6335; // @[ICache.scala 169:30]
  wire  _GEN_7889 = uncached ? _GEN_1873 : _GEN_6336; // @[ICache.scala 169:30]
  wire  _GEN_7890 = uncached ? _GEN_1362 : _GEN_6337; // @[ICache.scala 169:30]
  wire  _GEN_7891 = uncached ? _GEN_1874 : _GEN_6338; // @[ICache.scala 169:30]
  wire  _GEN_7892 = uncached ? _GEN_1363 : _GEN_6339; // @[ICache.scala 169:30]
  wire  _GEN_7893 = uncached ? _GEN_1875 : _GEN_6340; // @[ICache.scala 169:30]
  wire  _GEN_7894 = uncached ? _GEN_1364 : _GEN_6341; // @[ICache.scala 169:30]
  wire  _GEN_7895 = uncached ? _GEN_1876 : _GEN_6342; // @[ICache.scala 169:30]
  wire  _GEN_7896 = uncached ? _GEN_1365 : _GEN_6343; // @[ICache.scala 169:30]
  wire  _GEN_7897 = uncached ? _GEN_1877 : _GEN_6344; // @[ICache.scala 169:30]
  wire  _GEN_7898 = uncached ? _GEN_1366 : _GEN_6345; // @[ICache.scala 169:30]
  wire  _GEN_7899 = uncached ? _GEN_1878 : _GEN_6346; // @[ICache.scala 169:30]
  wire  _GEN_7900 = uncached ? _GEN_1367 : _GEN_6347; // @[ICache.scala 169:30]
  wire  _GEN_7901 = uncached ? _GEN_1879 : _GEN_6348; // @[ICache.scala 169:30]
  wire  _GEN_7902 = uncached ? _GEN_1368 : _GEN_6349; // @[ICache.scala 169:30]
  wire  _GEN_7903 = uncached ? _GEN_1880 : _GEN_6350; // @[ICache.scala 169:30]
  wire  _GEN_7904 = uncached ? _GEN_1369 : _GEN_6351; // @[ICache.scala 169:30]
  wire  _GEN_7905 = uncached ? _GEN_1881 : _GEN_6352; // @[ICache.scala 169:30]
  wire  _GEN_7906 = uncached ? _GEN_1370 : _GEN_6353; // @[ICache.scala 169:30]
  wire  _GEN_7907 = uncached ? _GEN_1882 : _GEN_6354; // @[ICache.scala 169:30]
  wire  _GEN_7908 = uncached ? _GEN_1371 : _GEN_6355; // @[ICache.scala 169:30]
  wire  _GEN_7909 = uncached ? _GEN_1883 : _GEN_6356; // @[ICache.scala 169:30]
  wire  _GEN_7910 = uncached ? _GEN_1372 : _GEN_6357; // @[ICache.scala 169:30]
  wire  _GEN_7911 = uncached ? _GEN_1884 : _GEN_6358; // @[ICache.scala 169:30]
  wire  _GEN_7912 = uncached ? _GEN_1373 : _GEN_6359; // @[ICache.scala 169:30]
  wire  _GEN_7913 = uncached ? _GEN_1885 : _GEN_6360; // @[ICache.scala 169:30]
  wire  _GEN_7914 = uncached ? _GEN_1374 : _GEN_6361; // @[ICache.scala 169:30]
  wire  _GEN_7915 = uncached ? _GEN_1886 : _GEN_6362; // @[ICache.scala 169:30]
  wire  _GEN_7916 = uncached ? _GEN_1375 : _GEN_6363; // @[ICache.scala 169:30]
  wire  _GEN_7917 = uncached ? _GEN_1887 : _GEN_6364; // @[ICache.scala 169:30]
  wire  _GEN_7918 = uncached ? _GEN_1376 : _GEN_6365; // @[ICache.scala 169:30]
  wire  _GEN_7919 = uncached ? _GEN_1888 : _GEN_6366; // @[ICache.scala 169:30]
  wire  _GEN_7920 = uncached ? _GEN_1377 : _GEN_6367; // @[ICache.scala 169:30]
  wire  _GEN_7921 = uncached ? _GEN_1889 : _GEN_6368; // @[ICache.scala 169:30]
  wire  _GEN_7922 = uncached ? _GEN_1378 : _GEN_6369; // @[ICache.scala 169:30]
  wire  _GEN_7923 = uncached ? _GEN_1890 : _GEN_6370; // @[ICache.scala 169:30]
  wire  _GEN_7924 = uncached ? _GEN_1379 : _GEN_6371; // @[ICache.scala 169:30]
  wire  _GEN_7925 = uncached ? _GEN_1891 : _GEN_6372; // @[ICache.scala 169:30]
  wire  _GEN_7926 = uncached ? _GEN_1380 : _GEN_6373; // @[ICache.scala 169:30]
  wire  _GEN_7927 = uncached ? _GEN_1892 : _GEN_6374; // @[ICache.scala 169:30]
  wire  _GEN_7928 = uncached ? _GEN_1381 : _GEN_6375; // @[ICache.scala 169:30]
  wire  _GEN_7929 = uncached ? _GEN_1893 : _GEN_6376; // @[ICache.scala 169:30]
  wire  _GEN_7930 = uncached ? _GEN_1382 : _GEN_6377; // @[ICache.scala 169:30]
  wire  _GEN_7931 = uncached ? _GEN_1894 : _GEN_6378; // @[ICache.scala 169:30]
  wire  _GEN_7932 = uncached ? _GEN_1383 : _GEN_6379; // @[ICache.scala 169:30]
  wire  _GEN_7933 = uncached ? _GEN_1895 : _GEN_6380; // @[ICache.scala 169:30]
  wire  _GEN_7934 = uncached ? _GEN_1384 : _GEN_6381; // @[ICache.scala 169:30]
  wire  _GEN_7935 = uncached ? _GEN_1896 : _GEN_6382; // @[ICache.scala 169:30]
  wire  _GEN_7936 = uncached ? _GEN_1385 : _GEN_6383; // @[ICache.scala 169:30]
  wire  _GEN_7937 = uncached ? _GEN_1897 : _GEN_6384; // @[ICache.scala 169:30]
  wire  _GEN_7938 = uncached ? _GEN_1386 : _GEN_6385; // @[ICache.scala 169:30]
  wire  _GEN_7939 = uncached ? _GEN_1898 : _GEN_6386; // @[ICache.scala 169:30]
  wire  _GEN_7940 = uncached ? _GEN_1387 : _GEN_6387; // @[ICache.scala 169:30]
  wire  _GEN_7941 = uncached ? _GEN_1899 : _GEN_6388; // @[ICache.scala 169:30]
  wire  _GEN_7942 = uncached ? _GEN_1388 : _GEN_6389; // @[ICache.scala 169:30]
  wire  _GEN_7943 = uncached ? _GEN_1900 : _GEN_6390; // @[ICache.scala 169:30]
  wire  _GEN_7944 = uncached ? _GEN_1389 : _GEN_6391; // @[ICache.scala 169:30]
  wire  _GEN_7945 = uncached ? _GEN_1901 : _GEN_6392; // @[ICache.scala 169:30]
  wire  _GEN_7946 = uncached ? _GEN_1390 : _GEN_6393; // @[ICache.scala 169:30]
  wire  _GEN_7947 = uncached ? _GEN_1902 : _GEN_6394; // @[ICache.scala 169:30]
  wire  _GEN_7948 = uncached ? _GEN_1391 : _GEN_6395; // @[ICache.scala 169:30]
  wire  _GEN_7949 = uncached ? _GEN_1903 : _GEN_6396; // @[ICache.scala 169:30]
  wire  _GEN_7950 = uncached ? _GEN_1392 : _GEN_6397; // @[ICache.scala 169:30]
  wire  _GEN_7951 = uncached ? _GEN_1904 : _GEN_6398; // @[ICache.scala 169:30]
  wire  _GEN_7952 = uncached ? _GEN_1393 : _GEN_6399; // @[ICache.scala 169:30]
  wire  _GEN_7953 = uncached ? _GEN_1905 : _GEN_6400; // @[ICache.scala 169:30]
  wire  _GEN_7954 = uncached ? _GEN_1394 : _GEN_6401; // @[ICache.scala 169:30]
  wire  _GEN_7955 = uncached ? _GEN_1906 : _GEN_6402; // @[ICache.scala 169:30]
  wire  _GEN_7956 = uncached ? _GEN_1395 : _GEN_6403; // @[ICache.scala 169:30]
  wire  _GEN_7957 = uncached ? _GEN_1907 : _GEN_6404; // @[ICache.scala 169:30]
  wire  _GEN_7958 = uncached ? _GEN_1396 : _GEN_6405; // @[ICache.scala 169:30]
  wire  _GEN_7959 = uncached ? _GEN_1908 : _GEN_6406; // @[ICache.scala 169:30]
  wire  _GEN_7960 = uncached ? _GEN_1397 : _GEN_6407; // @[ICache.scala 169:30]
  wire  _GEN_7961 = uncached ? _GEN_1909 : _GEN_6408; // @[ICache.scala 169:30]
  wire  _GEN_7962 = uncached ? _GEN_1398 : _GEN_6409; // @[ICache.scala 169:30]
  wire  _GEN_7963 = uncached ? _GEN_1910 : _GEN_6410; // @[ICache.scala 169:30]
  wire  _GEN_7964 = uncached ? _GEN_1399 : _GEN_6411; // @[ICache.scala 169:30]
  wire  _GEN_7965 = uncached ? _GEN_1911 : _GEN_6412; // @[ICache.scala 169:30]
  wire  _GEN_7966 = uncached ? _GEN_1400 : _GEN_6413; // @[ICache.scala 169:30]
  wire  _GEN_7967 = uncached ? _GEN_1912 : _GEN_6414; // @[ICache.scala 169:30]
  wire  _GEN_7968 = uncached ? _GEN_1401 : _GEN_6415; // @[ICache.scala 169:30]
  wire  _GEN_7969 = uncached ? _GEN_1913 : _GEN_6416; // @[ICache.scala 169:30]
  wire  _GEN_7970 = uncached ? _GEN_1402 : _GEN_6417; // @[ICache.scala 169:30]
  wire  _GEN_7971 = uncached ? _GEN_1914 : _GEN_6418; // @[ICache.scala 169:30]
  wire  _GEN_7972 = uncached ? _GEN_1403 : _GEN_6419; // @[ICache.scala 169:30]
  wire  _GEN_7973 = uncached ? _GEN_1915 : _GEN_6420; // @[ICache.scala 169:30]
  wire  _GEN_7974 = uncached ? _GEN_1404 : _GEN_6421; // @[ICache.scala 169:30]
  wire  _GEN_7975 = uncached ? _GEN_1916 : _GEN_6422; // @[ICache.scala 169:30]
  wire  _GEN_7976 = uncached ? _GEN_1405 : _GEN_6423; // @[ICache.scala 169:30]
  wire  _GEN_7977 = uncached ? _GEN_1917 : _GEN_6424; // @[ICache.scala 169:30]
  wire  _GEN_7978 = uncached ? _GEN_1406 : _GEN_6425; // @[ICache.scala 169:30]
  wire  _GEN_7979 = uncached ? _GEN_1918 : _GEN_6426; // @[ICache.scala 169:30]
  wire  _GEN_7980 = uncached ? _GEN_1407 : _GEN_6427; // @[ICache.scala 169:30]
  wire  _GEN_7981 = uncached ? _GEN_1919 : _GEN_6428; // @[ICache.scala 169:30]
  wire  _GEN_7982 = uncached ? _GEN_1408 : _GEN_6429; // @[ICache.scala 169:30]
  wire  _GEN_7983 = uncached ? _GEN_1920 : _GEN_6430; // @[ICache.scala 169:30]
  wire  _GEN_7984 = uncached ? _GEN_1409 : _GEN_6431; // @[ICache.scala 169:30]
  wire  _GEN_7985 = uncached ? _GEN_1921 : _GEN_6432; // @[ICache.scala 169:30]
  wire  _GEN_7986 = uncached ? _GEN_1410 : _GEN_6433; // @[ICache.scala 169:30]
  wire  _GEN_7987 = uncached ? _GEN_1922 : _GEN_6434; // @[ICache.scala 169:30]
  wire  _GEN_7988 = uncached ? _GEN_1411 : _GEN_6435; // @[ICache.scala 169:30]
  wire  _GEN_7989 = uncached ? _GEN_1923 : _GEN_6436; // @[ICache.scala 169:30]
  wire  _GEN_7990 = uncached ? _GEN_1412 : _GEN_6437; // @[ICache.scala 169:30]
  wire  _GEN_7991 = uncached ? _GEN_1924 : _GEN_6438; // @[ICache.scala 169:30]
  wire  _GEN_7992 = uncached ? _GEN_1413 : _GEN_6439; // @[ICache.scala 169:30]
  wire  _GEN_7993 = uncached ? _GEN_1925 : _GEN_6440; // @[ICache.scala 169:30]
  wire  _GEN_7994 = uncached ? _GEN_1414 : _GEN_6441; // @[ICache.scala 169:30]
  wire  _GEN_7995 = uncached ? _GEN_1926 : _GEN_6442; // @[ICache.scala 169:30]
  wire  _GEN_7996 = uncached ? _GEN_1415 : _GEN_6443; // @[ICache.scala 169:30]
  wire  _GEN_7997 = uncached ? _GEN_1927 : _GEN_6444; // @[ICache.scala 169:30]
  wire  _GEN_7998 = uncached ? _GEN_1416 : _GEN_6445; // @[ICache.scala 169:30]
  wire  _GEN_7999 = uncached ? _GEN_1928 : _GEN_6446; // @[ICache.scala 169:30]
  wire  _GEN_8000 = uncached ? _GEN_1417 : _GEN_6447; // @[ICache.scala 169:30]
  wire  _GEN_8001 = uncached ? _GEN_1929 : _GEN_6448; // @[ICache.scala 169:30]
  wire  _GEN_8002 = uncached ? _GEN_1418 : _GEN_6449; // @[ICache.scala 169:30]
  wire  _GEN_8003 = uncached ? _GEN_1930 : _GEN_6450; // @[ICache.scala 169:30]
  wire  _GEN_8004 = uncached ? _GEN_1419 : _GEN_6451; // @[ICache.scala 169:30]
  wire  _GEN_8005 = uncached ? _GEN_1931 : _GEN_6452; // @[ICache.scala 169:30]
  wire  _GEN_8006 = uncached ? _GEN_1420 : _GEN_6453; // @[ICache.scala 169:30]
  wire  _GEN_8007 = uncached ? _GEN_1932 : _GEN_6454; // @[ICache.scala 169:30]
  wire  _GEN_8008 = uncached ? _GEN_1421 : _GEN_6455; // @[ICache.scala 169:30]
  wire  _GEN_8009 = uncached ? _GEN_1933 : _GEN_6456; // @[ICache.scala 169:30]
  wire  _GEN_8010 = uncached ? _GEN_1422 : _GEN_6457; // @[ICache.scala 169:30]
  wire  _GEN_8011 = uncached ? _GEN_1934 : _GEN_6458; // @[ICache.scala 169:30]
  wire  _GEN_8012 = uncached ? _GEN_1423 : _GEN_6459; // @[ICache.scala 169:30]
  wire  _GEN_8013 = uncached ? _GEN_1935 : _GEN_6460; // @[ICache.scala 169:30]
  wire  _GEN_8014 = uncached ? _GEN_1424 : _GEN_6461; // @[ICache.scala 169:30]
  wire  _GEN_8015 = uncached ? _GEN_1936 : _GEN_6462; // @[ICache.scala 169:30]
  wire  _GEN_8016 = uncached ? _GEN_1425 : _GEN_6463; // @[ICache.scala 169:30]
  wire  _GEN_8017 = uncached ? _GEN_1937 : _GEN_6464; // @[ICache.scala 169:30]
  wire  _GEN_8018 = uncached ? _GEN_1426 : _GEN_6465; // @[ICache.scala 169:30]
  wire  _GEN_8019 = uncached ? _GEN_1938 : _GEN_6466; // @[ICache.scala 169:30]
  wire  _GEN_8020 = uncached ? _GEN_1427 : _GEN_6467; // @[ICache.scala 169:30]
  wire  _GEN_8021 = uncached ? _GEN_1939 : _GEN_6468; // @[ICache.scala 169:30]
  wire  _GEN_8022 = uncached ? _GEN_1428 : _GEN_6469; // @[ICache.scala 169:30]
  wire  _GEN_8023 = uncached ? _GEN_1940 : _GEN_6470; // @[ICache.scala 169:30]
  wire  _GEN_8024 = uncached ? _GEN_1429 : _GEN_6471; // @[ICache.scala 169:30]
  wire  _GEN_8025 = uncached ? _GEN_1941 : _GEN_6472; // @[ICache.scala 169:30]
  wire  _GEN_8026 = uncached ? _GEN_1430 : _GEN_6473; // @[ICache.scala 169:30]
  wire  _GEN_8027 = uncached ? _GEN_1942 : _GEN_6474; // @[ICache.scala 169:30]
  wire  _GEN_8028 = uncached ? _GEN_1431 : _GEN_6475; // @[ICache.scala 169:30]
  wire  _GEN_8029 = uncached ? _GEN_1943 : _GEN_6476; // @[ICache.scala 169:30]
  wire  _GEN_8030 = uncached ? _GEN_1432 : _GEN_6477; // @[ICache.scala 169:30]
  wire  _GEN_8031 = uncached ? _GEN_1944 : _GEN_6478; // @[ICache.scala 169:30]
  wire  _GEN_8032 = uncached ? _GEN_1433 : _GEN_6479; // @[ICache.scala 169:30]
  wire  _GEN_8033 = uncached ? _GEN_1945 : _GEN_6480; // @[ICache.scala 169:30]
  wire  _GEN_8034 = uncached ? _GEN_1434 : _GEN_6481; // @[ICache.scala 169:30]
  wire  _GEN_8035 = uncached ? _GEN_1946 : _GEN_6482; // @[ICache.scala 169:30]
  wire  _GEN_8036 = uncached ? _GEN_1435 : _GEN_6483; // @[ICache.scala 169:30]
  wire  _GEN_8037 = uncached ? _GEN_1947 : _GEN_6484; // @[ICache.scala 169:30]
  wire  _GEN_8038 = uncached ? _GEN_1436 : _GEN_6485; // @[ICache.scala 169:30]
  wire  _GEN_8039 = uncached ? _GEN_1948 : _GEN_6486; // @[ICache.scala 169:30]
  wire  _GEN_8040 = uncached ? _GEN_1437 : _GEN_6487; // @[ICache.scala 169:30]
  wire  _GEN_8041 = uncached ? _GEN_1949 : _GEN_6488; // @[ICache.scala 169:30]
  wire  _GEN_8042 = uncached ? _GEN_1438 : _GEN_6489; // @[ICache.scala 169:30]
  wire  _GEN_8043 = uncached ? _GEN_1950 : _GEN_6490; // @[ICache.scala 169:30]
  wire  _GEN_8044 = uncached ? _GEN_1439 : _GEN_6491; // @[ICache.scala 169:30]
  wire  _GEN_8045 = uncached ? _GEN_1951 : _GEN_6492; // @[ICache.scala 169:30]
  wire  _GEN_8046 = uncached ? _GEN_1440 : _GEN_6493; // @[ICache.scala 169:30]
  wire  _GEN_8047 = uncached ? _GEN_1952 : _GEN_6494; // @[ICache.scala 169:30]
  wire  _GEN_8048 = uncached ? _GEN_1441 : _GEN_6495; // @[ICache.scala 169:30]
  wire  _GEN_8049 = uncached ? _GEN_1953 : _GEN_6496; // @[ICache.scala 169:30]
  wire  _GEN_8050 = uncached ? _GEN_1442 : _GEN_6497; // @[ICache.scala 169:30]
  wire  _GEN_8051 = uncached ? _GEN_1954 : _GEN_6498; // @[ICache.scala 169:30]
  wire  _GEN_8052 = uncached ? _GEN_1443 : _GEN_6499; // @[ICache.scala 169:30]
  wire  _GEN_8053 = uncached ? _GEN_1955 : _GEN_6500; // @[ICache.scala 169:30]
  wire  _GEN_8054 = uncached ? _GEN_1444 : _GEN_6501; // @[ICache.scala 169:30]
  wire  _GEN_8055 = uncached ? _GEN_1956 : _GEN_6502; // @[ICache.scala 169:30]
  wire  _GEN_8056 = uncached ? _GEN_1445 : _GEN_6503; // @[ICache.scala 169:30]
  wire  _GEN_8057 = uncached ? _GEN_1957 : _GEN_6504; // @[ICache.scala 169:30]
  wire  _GEN_8058 = uncached ? _GEN_1446 : _GEN_6505; // @[ICache.scala 169:30]
  wire  _GEN_8059 = uncached ? _GEN_1958 : _GEN_6506; // @[ICache.scala 169:30]
  wire  _GEN_8060 = uncached ? _GEN_1447 : _GEN_6507; // @[ICache.scala 169:30]
  wire  _GEN_8061 = uncached ? _GEN_1959 : _GEN_6508; // @[ICache.scala 169:30]
  wire  _GEN_8062 = uncached ? _GEN_1448 : _GEN_6509; // @[ICache.scala 169:30]
  wire  _GEN_8063 = uncached ? _GEN_1960 : _GEN_6510; // @[ICache.scala 169:30]
  wire  _GEN_8064 = uncached ? _GEN_1449 : _GEN_6511; // @[ICache.scala 169:30]
  wire  _GEN_8065 = uncached ? _GEN_1961 : _GEN_6512; // @[ICache.scala 169:30]
  wire  _GEN_8066 = uncached ? _GEN_1450 : _GEN_6513; // @[ICache.scala 169:30]
  wire  _GEN_8067 = uncached ? _GEN_1962 : _GEN_6514; // @[ICache.scala 169:30]
  wire  _GEN_8068 = uncached ? _GEN_1451 : _GEN_6515; // @[ICache.scala 169:30]
  wire  _GEN_8069 = uncached ? _GEN_1963 : _GEN_6516; // @[ICache.scala 169:30]
  wire  _GEN_8070 = uncached ? _GEN_1452 : _GEN_6517; // @[ICache.scala 169:30]
  wire  _GEN_8071 = uncached ? _GEN_1964 : _GEN_6518; // @[ICache.scala 169:30]
  wire  _GEN_8072 = uncached ? _GEN_1453 : _GEN_6519; // @[ICache.scala 169:30]
  wire  _GEN_8073 = uncached ? _GEN_1965 : _GEN_6520; // @[ICache.scala 169:30]
  wire  _GEN_8074 = uncached ? _GEN_1454 : _GEN_6521; // @[ICache.scala 169:30]
  wire  _GEN_8075 = uncached ? _GEN_1966 : _GEN_6522; // @[ICache.scala 169:30]
  wire  _GEN_8076 = uncached ? _GEN_1455 : _GEN_6523; // @[ICache.scala 169:30]
  wire  _GEN_8077 = uncached ? _GEN_1967 : _GEN_6524; // @[ICache.scala 169:30]
  wire  _GEN_8078 = uncached ? _GEN_1456 : _GEN_6525; // @[ICache.scala 169:30]
  wire  _GEN_8079 = uncached ? _GEN_1968 : _GEN_6526; // @[ICache.scala 169:30]
  wire  _GEN_8080 = uncached ? _GEN_1457 : _GEN_6527; // @[ICache.scala 169:30]
  wire  _GEN_8081 = uncached ? _GEN_1969 : _GEN_6528; // @[ICache.scala 169:30]
  wire  _GEN_8082 = uncached ? _GEN_1458 : _GEN_6529; // @[ICache.scala 169:30]
  wire  _GEN_8083 = uncached ? _GEN_1970 : _GEN_6530; // @[ICache.scala 169:30]
  wire  _GEN_8084 = uncached ? _GEN_1459 : _GEN_6531; // @[ICache.scala 169:30]
  wire  _GEN_8085 = uncached ? _GEN_1971 : _GEN_6532; // @[ICache.scala 169:30]
  wire  _GEN_8086 = uncached ? _GEN_1460 : _GEN_6533; // @[ICache.scala 169:30]
  wire  _GEN_8087 = uncached ? _GEN_1972 : _GEN_6534; // @[ICache.scala 169:30]
  wire  _GEN_8088 = uncached ? _GEN_1461 : _GEN_6535; // @[ICache.scala 169:30]
  wire  _GEN_8089 = uncached ? _GEN_1973 : _GEN_6536; // @[ICache.scala 169:30]
  wire  _GEN_8090 = uncached ? _GEN_1462 : _GEN_6537; // @[ICache.scala 169:30]
  wire  _GEN_8091 = uncached ? _GEN_1974 : _GEN_6538; // @[ICache.scala 169:30]
  wire  _GEN_8092 = uncached ? _GEN_1463 : _GEN_6539; // @[ICache.scala 169:30]
  wire  _GEN_8093 = uncached ? _GEN_1975 : _GEN_6540; // @[ICache.scala 169:30]
  wire  _GEN_8094 = uncached ? _GEN_1464 : _GEN_6541; // @[ICache.scala 169:30]
  wire  _GEN_8095 = uncached ? _GEN_1976 : _GEN_6542; // @[ICache.scala 169:30]
  wire  _GEN_8096 = uncached ? _GEN_1465 : _GEN_6543; // @[ICache.scala 169:30]
  wire  _GEN_8097 = uncached ? _GEN_1977 : _GEN_6544; // @[ICache.scala 169:30]
  wire  _GEN_8098 = uncached ? _GEN_1466 : _GEN_6545; // @[ICache.scala 169:30]
  wire  _GEN_8099 = uncached ? _GEN_1978 : _GEN_6546; // @[ICache.scala 169:30]
  wire  _GEN_8100 = uncached ? _GEN_1467 : _GEN_6547; // @[ICache.scala 169:30]
  wire  _GEN_8101 = uncached ? _GEN_1979 : _GEN_6548; // @[ICache.scala 169:30]
  wire  _GEN_8102 = uncached ? _GEN_1468 : _GEN_6549; // @[ICache.scala 169:30]
  wire  _GEN_8103 = uncached ? _GEN_1980 : _GEN_6550; // @[ICache.scala 169:30]
  wire  _GEN_8104 = uncached ? _GEN_1469 : _GEN_6551; // @[ICache.scala 169:30]
  wire  _GEN_8105 = uncached ? _GEN_1981 : _GEN_6552; // @[ICache.scala 169:30]
  wire  _GEN_8106 = uncached ? _GEN_1470 : _GEN_6553; // @[ICache.scala 169:30]
  wire  _GEN_8107 = uncached ? _GEN_1982 : _GEN_6554; // @[ICache.scala 169:30]
  wire  _GEN_8108 = uncached ? _GEN_1471 : _GEN_6555; // @[ICache.scala 169:30]
  wire  _GEN_8109 = uncached ? _GEN_1983 : _GEN_6556; // @[ICache.scala 169:30]
  wire  _GEN_8110 = uncached ? _GEN_1472 : _GEN_6557; // @[ICache.scala 169:30]
  wire  _GEN_8111 = uncached ? _GEN_1984 : _GEN_6558; // @[ICache.scala 169:30]
  wire  _GEN_8112 = uncached ? _GEN_1473 : _GEN_6559; // @[ICache.scala 169:30]
  wire  _GEN_8113 = uncached ? _GEN_1985 : _GEN_6560; // @[ICache.scala 169:30]
  wire  _GEN_8114 = uncached ? _GEN_1474 : _GEN_6561; // @[ICache.scala 169:30]
  wire  _GEN_8115 = uncached ? _GEN_1986 : _GEN_6562; // @[ICache.scala 169:30]
  wire  _GEN_8116 = uncached ? _GEN_1475 : _GEN_6563; // @[ICache.scala 169:30]
  wire  _GEN_8117 = uncached ? _GEN_1987 : _GEN_6564; // @[ICache.scala 169:30]
  wire  _GEN_8118 = uncached ? _GEN_1476 : _GEN_6565; // @[ICache.scala 169:30]
  wire  _GEN_8119 = uncached ? _GEN_1988 : _GEN_6566; // @[ICache.scala 169:30]
  wire  _GEN_8120 = uncached ? _GEN_1477 : _GEN_6567; // @[ICache.scala 169:30]
  wire  _GEN_8121 = uncached ? _GEN_1989 : _GEN_6568; // @[ICache.scala 169:30]
  wire  _GEN_8122 = uncached ? _GEN_1478 : _GEN_6569; // @[ICache.scala 169:30]
  wire  _GEN_8123 = uncached ? _GEN_1990 : _GEN_6570; // @[ICache.scala 169:30]
  wire  _GEN_8124 = uncached ? _GEN_1479 : _GEN_6571; // @[ICache.scala 169:30]
  wire  _GEN_8125 = uncached ? _GEN_1991 : _GEN_6572; // @[ICache.scala 169:30]
  wire  _GEN_8126 = uncached ? _GEN_1480 : _GEN_6573; // @[ICache.scala 169:30]
  wire  _GEN_8127 = uncached ? _GEN_1992 : _GEN_6574; // @[ICache.scala 169:30]
  wire  _GEN_8128 = uncached ? _GEN_1481 : _GEN_6575; // @[ICache.scala 169:30]
  wire  _GEN_8129 = uncached ? _GEN_1993 : _GEN_6576; // @[ICache.scala 169:30]
  wire  _GEN_8130 = uncached ? _GEN_1482 : _GEN_6577; // @[ICache.scala 169:30]
  wire  _GEN_8131 = uncached ? _GEN_1994 : _GEN_6578; // @[ICache.scala 169:30]
  wire  _GEN_8132 = uncached ? _GEN_1483 : _GEN_6579; // @[ICache.scala 169:30]
  wire  _GEN_8133 = uncached ? _GEN_1995 : _GEN_6580; // @[ICache.scala 169:30]
  wire  _GEN_8134 = uncached ? _GEN_1484 : _GEN_6581; // @[ICache.scala 169:30]
  wire  _GEN_8135 = uncached ? _GEN_1996 : _GEN_6582; // @[ICache.scala 169:30]
  wire  _GEN_8136 = uncached ? _GEN_1485 : _GEN_6583; // @[ICache.scala 169:30]
  wire  _GEN_8137 = uncached ? _GEN_1997 : _GEN_6584; // @[ICache.scala 169:30]
  wire  _GEN_8138 = uncached ? _GEN_1486 : _GEN_6585; // @[ICache.scala 169:30]
  wire  _GEN_8139 = uncached ? _GEN_1998 : _GEN_6586; // @[ICache.scala 169:30]
  wire  _GEN_8140 = uncached ? _GEN_1487 : _GEN_6587; // @[ICache.scala 169:30]
  wire  _GEN_8141 = uncached ? _GEN_1999 : _GEN_6588; // @[ICache.scala 169:30]
  wire  _GEN_8142 = uncached ? _GEN_1488 : _GEN_6589; // @[ICache.scala 169:30]
  wire  _GEN_8143 = uncached ? _GEN_2000 : _GEN_6590; // @[ICache.scala 169:30]
  wire  _GEN_8144 = uncached ? _GEN_1489 : _GEN_6591; // @[ICache.scala 169:30]
  wire  _GEN_8145 = uncached ? _GEN_2001 : _GEN_6592; // @[ICache.scala 169:30]
  wire  _GEN_8146 = uncached ? _GEN_1490 : _GEN_6593; // @[ICache.scala 169:30]
  wire  _GEN_8147 = uncached ? _GEN_2002 : _GEN_6594; // @[ICache.scala 169:30]
  wire  _GEN_8148 = uncached ? _GEN_1491 : _GEN_6595; // @[ICache.scala 169:30]
  wire  _GEN_8149 = uncached ? _GEN_2003 : _GEN_6596; // @[ICache.scala 169:30]
  wire  _GEN_8150 = uncached ? _GEN_1492 : _GEN_6597; // @[ICache.scala 169:30]
  wire  _GEN_8151 = uncached ? _GEN_2004 : _GEN_6598; // @[ICache.scala 169:30]
  wire  _GEN_8152 = uncached ? _GEN_1493 : _GEN_6599; // @[ICache.scala 169:30]
  wire  _GEN_8153 = uncached ? _GEN_2005 : _GEN_6600; // @[ICache.scala 169:30]
  wire  _GEN_8154 = uncached ? _GEN_1494 : _GEN_6601; // @[ICache.scala 169:30]
  wire  _GEN_8155 = uncached ? _GEN_2006 : _GEN_6602; // @[ICache.scala 169:30]
  wire  _GEN_8156 = uncached ? _GEN_1495 : _GEN_6603; // @[ICache.scala 169:30]
  wire  _GEN_8157 = uncached ? _GEN_2007 : _GEN_6604; // @[ICache.scala 169:30]
  wire  _GEN_8158 = uncached ? _GEN_1496 : _GEN_6605; // @[ICache.scala 169:30]
  wire  _GEN_8159 = uncached ? _GEN_2008 : _GEN_6606; // @[ICache.scala 169:30]
  wire  _GEN_8160 = uncached ? _GEN_1497 : _GEN_6607; // @[ICache.scala 169:30]
  wire  _GEN_8161 = uncached ? _GEN_2009 : _GEN_6608; // @[ICache.scala 169:30]
  wire  _GEN_8162 = uncached ? _GEN_1498 : _GEN_6609; // @[ICache.scala 169:30]
  wire  _GEN_8163 = uncached ? _GEN_2010 : _GEN_6610; // @[ICache.scala 169:30]
  wire  _GEN_8164 = uncached ? _GEN_1499 : _GEN_6611; // @[ICache.scala 169:30]
  wire  _GEN_8165 = uncached ? _GEN_2011 : _GEN_6612; // @[ICache.scala 169:30]
  wire  _GEN_8166 = uncached ? _GEN_1500 : _GEN_6613; // @[ICache.scala 169:30]
  wire  _GEN_8167 = uncached ? _GEN_2012 : _GEN_6614; // @[ICache.scala 169:30]
  wire  _GEN_8168 = uncached ? _GEN_1501 : _GEN_6615; // @[ICache.scala 169:30]
  wire  _GEN_8169 = uncached ? _GEN_2013 : _GEN_6616; // @[ICache.scala 169:30]
  wire  _GEN_8170 = uncached ? _GEN_1502 : _GEN_6617; // @[ICache.scala 169:30]
  wire  _GEN_8171 = uncached ? _GEN_2014 : _GEN_6618; // @[ICache.scala 169:30]
  wire  _GEN_8172 = uncached ? _GEN_1503 : _GEN_6619; // @[ICache.scala 169:30]
  wire  _GEN_8173 = uncached ? _GEN_2015 : _GEN_6620; // @[ICache.scala 169:30]
  wire  _GEN_8174 = uncached ? _GEN_1504 : _GEN_6621; // @[ICache.scala 169:30]
  wire  _GEN_8175 = uncached ? _GEN_2016 : _GEN_6622; // @[ICache.scala 169:30]
  wire  _GEN_8176 = uncached ? _GEN_1505 : _GEN_6623; // @[ICache.scala 169:30]
  wire  _GEN_8177 = uncached ? _GEN_2017 : _GEN_6624; // @[ICache.scala 169:30]
  wire  _GEN_8178 = uncached ? _GEN_1506 : _GEN_6625; // @[ICache.scala 169:30]
  wire  _GEN_8179 = uncached ? _GEN_2018 : _GEN_6626; // @[ICache.scala 169:30]
  wire  _GEN_8180 = uncached ? _GEN_1507 : _GEN_6627; // @[ICache.scala 169:30]
  wire  _GEN_8181 = uncached ? _GEN_2019 : _GEN_6628; // @[ICache.scala 169:30]
  wire  _GEN_8182 = uncached ? _GEN_1508 : _GEN_6629; // @[ICache.scala 169:30]
  wire  _GEN_8183 = uncached ? _GEN_2020 : _GEN_6630; // @[ICache.scala 169:30]
  wire  _GEN_8184 = uncached ? _GEN_1509 : _GEN_6631; // @[ICache.scala 169:30]
  wire  _GEN_8185 = uncached ? _GEN_2021 : _GEN_6632; // @[ICache.scala 169:30]
  wire  _GEN_8186 = uncached ? _GEN_1510 : _GEN_6633; // @[ICache.scala 169:30]
  wire  _GEN_8187 = uncached ? _GEN_2022 : _GEN_6634; // @[ICache.scala 169:30]
  wire  _GEN_8188 = uncached ? _GEN_1511 : _GEN_6635; // @[ICache.scala 169:30]
  wire  _GEN_8189 = uncached ? _GEN_2023 : _GEN_6636; // @[ICache.scala 169:30]
  wire  _GEN_8190 = uncached ? _GEN_1512 : _GEN_6637; // @[ICache.scala 169:30]
  wire  _GEN_8191 = uncached ? _GEN_2024 : _GEN_6638; // @[ICache.scala 169:30]
  wire  _GEN_8192 = uncached ? _GEN_1513 : _GEN_6639; // @[ICache.scala 169:30]
  wire  _GEN_8193 = uncached ? _GEN_2025 : _GEN_6640; // @[ICache.scala 169:30]
  wire  _GEN_8194 = uncached ? _GEN_1514 : _GEN_6641; // @[ICache.scala 169:30]
  wire  _GEN_8195 = uncached ? _GEN_2026 : _GEN_6642; // @[ICache.scala 169:30]
  wire  _GEN_8196 = uncached ? _GEN_1515 : _GEN_6643; // @[ICache.scala 169:30]
  wire  _GEN_8197 = uncached ? _GEN_2027 : _GEN_6644; // @[ICache.scala 169:30]
  wire  _GEN_8198 = uncached ? _GEN_1516 : _GEN_6645; // @[ICache.scala 169:30]
  wire  _GEN_8199 = uncached ? _GEN_2028 : _GEN_6646; // @[ICache.scala 169:30]
  wire  _GEN_8200 = uncached ? _GEN_1517 : _GEN_6647; // @[ICache.scala 169:30]
  wire  _GEN_8201 = uncached ? _GEN_2029 : _GEN_6648; // @[ICache.scala 169:30]
  wire  _GEN_8202 = uncached ? _GEN_1518 : _GEN_6649; // @[ICache.scala 169:30]
  wire  _GEN_8203 = uncached ? _GEN_2030 : _GEN_6650; // @[ICache.scala 169:30]
  wire  _GEN_8204 = uncached ? _GEN_1519 : _GEN_6651; // @[ICache.scala 169:30]
  wire  _GEN_8205 = uncached ? _GEN_2031 : _GEN_6652; // @[ICache.scala 169:30]
  wire  _GEN_8206 = uncached ? _GEN_1520 : _GEN_6653; // @[ICache.scala 169:30]
  wire  _GEN_8207 = uncached ? _GEN_2032 : _GEN_6654; // @[ICache.scala 169:30]
  wire  _GEN_8208 = uncached ? _GEN_1521 : _GEN_6655; // @[ICache.scala 169:30]
  wire  _GEN_8209 = uncached ? _GEN_2033 : _GEN_6656; // @[ICache.scala 169:30]
  wire  _GEN_8210 = uncached ? _GEN_1522 : _GEN_6657; // @[ICache.scala 169:30]
  wire  _GEN_8211 = uncached ? _GEN_2034 : _GEN_6658; // @[ICache.scala 169:30]
  wire  _GEN_8212 = uncached ? _GEN_1523 : _GEN_6659; // @[ICache.scala 169:30]
  wire  _GEN_8213 = uncached ? _GEN_2035 : _GEN_6660; // @[ICache.scala 169:30]
  wire  _GEN_8214 = uncached ? _GEN_1524 : _GEN_6661; // @[ICache.scala 169:30]
  wire  _GEN_8215 = uncached ? _GEN_2036 : _GEN_6662; // @[ICache.scala 169:30]
  wire  _GEN_8216 = uncached ? _GEN_1525 : _GEN_6663; // @[ICache.scala 169:30]
  wire  _GEN_8217 = uncached ? _GEN_2037 : _GEN_6664; // @[ICache.scala 169:30]
  wire  _GEN_8218 = uncached ? _GEN_1526 : _GEN_6665; // @[ICache.scala 169:30]
  wire  _GEN_8219 = uncached ? _GEN_2038 : _GEN_6666; // @[ICache.scala 169:30]
  wire  _GEN_8220 = uncached ? _GEN_1527 : _GEN_6667; // @[ICache.scala 169:30]
  wire  _GEN_8221 = uncached ? _GEN_2039 : _GEN_6668; // @[ICache.scala 169:30]
  wire  _GEN_8222 = uncached ? _GEN_1528 : _GEN_6669; // @[ICache.scala 169:30]
  wire  _GEN_8223 = uncached ? _GEN_2040 : _GEN_6670; // @[ICache.scala 169:30]
  wire  _GEN_8224 = uncached ? _GEN_1529 : _GEN_6671; // @[ICache.scala 169:30]
  wire  _GEN_8225 = uncached ? _GEN_2041 : _GEN_6672; // @[ICache.scala 169:30]
  wire  _GEN_8226 = uncached ? _GEN_1530 : _GEN_6673; // @[ICache.scala 169:30]
  wire  _GEN_8227 = uncached ? _GEN_2042 : _GEN_6674; // @[ICache.scala 169:30]
  wire  _GEN_8228 = uncached ? _GEN_1531 : _GEN_6675; // @[ICache.scala 169:30]
  wire  _GEN_8229 = uncached ? _GEN_2043 : _GEN_6676; // @[ICache.scala 169:30]
  wire  _GEN_8230 = uncached ? _GEN_1532 : _GEN_6677; // @[ICache.scala 169:30]
  wire  _GEN_8231 = uncached ? _GEN_2044 : _GEN_6678; // @[ICache.scala 169:30]
  wire  _GEN_8232 = uncached ? _GEN_1533 : _GEN_6679; // @[ICache.scala 169:30]
  wire  _GEN_8233 = uncached ? _GEN_2045 : _GEN_6680; // @[ICache.scala 169:30]
  wire  _GEN_8234 = uncached ? _GEN_1534 : _GEN_6681; // @[ICache.scala 169:30]
  wire  _GEN_8235 = uncached ? _GEN_2046 : _GEN_6682; // @[ICache.scala 169:30]
  wire  _GEN_8236 = uncached ? _GEN_1535 : _GEN_6683; // @[ICache.scala 169:30]
  wire  _GEN_8237 = uncached ? _GEN_2047 : _GEN_6684; // @[ICache.scala 169:30]
  wire  _GEN_8238 = uncached ? _GEN_1536 : _GEN_6685; // @[ICache.scala 169:30]
  wire  _GEN_8239 = uncached ? _GEN_2048 : _GEN_6686; // @[ICache.scala 169:30]
  wire  _GEN_8240 = uncached ? _GEN_1537 : _GEN_6687; // @[ICache.scala 169:30]
  wire  _GEN_8241 = uncached ? _GEN_2049 : _GEN_6688; // @[ICache.scala 169:30]
  wire  _GEN_8242 = uncached ? _GEN_1538 : _GEN_6689; // @[ICache.scala 169:30]
  wire  _GEN_8243 = uncached ? _GEN_2050 : _GEN_6690; // @[ICache.scala 169:30]
  wire [4:0] _GEN_8244 = uncached ? axi_cnt_value : _GEN_6691; // @[ICache.scala 169:30 Counter.scala 61:40]
  wire  _GEN_8245 = uncached ? lru_0 : _GEN_6692; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8246 = uncached ? lru_1 : _GEN_6693; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8247 = uncached ? lru_2 : _GEN_6694; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8248 = uncached ? lru_3 : _GEN_6695; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8249 = uncached ? lru_4 : _GEN_6696; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8250 = uncached ? lru_5 : _GEN_6697; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8251 = uncached ? lru_6 : _GEN_6698; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8252 = uncached ? lru_7 : _GEN_6699; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8253 = uncached ? lru_8 : _GEN_6700; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8254 = uncached ? lru_9 : _GEN_6701; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8255 = uncached ? lru_10 : _GEN_6702; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8256 = uncached ? lru_11 : _GEN_6703; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8257 = uncached ? lru_12 : _GEN_6704; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8258 = uncached ? lru_13 : _GEN_6705; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8259 = uncached ? lru_14 : _GEN_6706; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8260 = uncached ? lru_15 : _GEN_6707; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8261 = uncached ? lru_16 : _GEN_6708; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8262 = uncached ? lru_17 : _GEN_6709; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8263 = uncached ? lru_18 : _GEN_6710; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8264 = uncached ? lru_19 : _GEN_6711; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8265 = uncached ? lru_20 : _GEN_6712; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8266 = uncached ? lru_21 : _GEN_6713; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8267 = uncached ? lru_22 : _GEN_6714; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8268 = uncached ? lru_23 : _GEN_6715; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8269 = uncached ? lru_24 : _GEN_6716; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8270 = uncached ? lru_25 : _GEN_6717; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8271 = uncached ? lru_26 : _GEN_6718; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8272 = uncached ? lru_27 : _GEN_6719; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8273 = uncached ? lru_28 : _GEN_6720; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8274 = uncached ? lru_29 : _GEN_6721; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8275 = uncached ? lru_30 : _GEN_6722; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8276 = uncached ? lru_31 : _GEN_6723; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8277 = uncached ? lru_32 : _GEN_6724; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8278 = uncached ? lru_33 : _GEN_6725; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8279 = uncached ? lru_34 : _GEN_6726; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8280 = uncached ? lru_35 : _GEN_6727; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8281 = uncached ? lru_36 : _GEN_6728; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8282 = uncached ? lru_37 : _GEN_6729; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8283 = uncached ? lru_38 : _GEN_6730; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8284 = uncached ? lru_39 : _GEN_6731; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8285 = uncached ? lru_40 : _GEN_6732; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8286 = uncached ? lru_41 : _GEN_6733; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8287 = uncached ? lru_42 : _GEN_6734; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8288 = uncached ? lru_43 : _GEN_6735; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8289 = uncached ? lru_44 : _GEN_6736; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8290 = uncached ? lru_45 : _GEN_6737; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8291 = uncached ? lru_46 : _GEN_6738; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8292 = uncached ? lru_47 : _GEN_6739; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8293 = uncached ? lru_48 : _GEN_6740; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8294 = uncached ? lru_49 : _GEN_6741; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8295 = uncached ? lru_50 : _GEN_6742; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8296 = uncached ? lru_51 : _GEN_6743; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8297 = uncached ? lru_52 : _GEN_6744; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8298 = uncached ? lru_53 : _GEN_6745; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8299 = uncached ? lru_54 : _GEN_6746; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8300 = uncached ? lru_55 : _GEN_6747; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8301 = uncached ? lru_56 : _GEN_6748; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8302 = uncached ? lru_57 : _GEN_6749; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8303 = uncached ? lru_58 : _GEN_6750; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8304 = uncached ? lru_59 : _GEN_6751; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8305 = uncached ? lru_60 : _GEN_6752; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8306 = uncached ? lru_61 : _GEN_6753; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8307 = uncached ? lru_62 : _GEN_6754; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8308 = uncached ? lru_63 : _GEN_6755; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8309 = uncached ? lru_64 : _GEN_6756; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8310 = uncached ? lru_65 : _GEN_6757; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8311 = uncached ? lru_66 : _GEN_6758; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8312 = uncached ? lru_67 : _GEN_6759; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8313 = uncached ? lru_68 : _GEN_6760; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8314 = uncached ? lru_69 : _GEN_6761; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8315 = uncached ? lru_70 : _GEN_6762; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8316 = uncached ? lru_71 : _GEN_6763; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8317 = uncached ? lru_72 : _GEN_6764; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8318 = uncached ? lru_73 : _GEN_6765; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8319 = uncached ? lru_74 : _GEN_6766; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8320 = uncached ? lru_75 : _GEN_6767; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8321 = uncached ? lru_76 : _GEN_6768; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8322 = uncached ? lru_77 : _GEN_6769; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8323 = uncached ? lru_78 : _GEN_6770; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8324 = uncached ? lru_79 : _GEN_6771; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8325 = uncached ? lru_80 : _GEN_6772; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8326 = uncached ? lru_81 : _GEN_6773; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8327 = uncached ? lru_82 : _GEN_6774; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8328 = uncached ? lru_83 : _GEN_6775; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8329 = uncached ? lru_84 : _GEN_6776; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8330 = uncached ? lru_85 : _GEN_6777; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8331 = uncached ? lru_86 : _GEN_6778; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8332 = uncached ? lru_87 : _GEN_6779; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8333 = uncached ? lru_88 : _GEN_6780; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8334 = uncached ? lru_89 : _GEN_6781; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8335 = uncached ? lru_90 : _GEN_6782; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8336 = uncached ? lru_91 : _GEN_6783; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8337 = uncached ? lru_92 : _GEN_6784; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8338 = uncached ? lru_93 : _GEN_6785; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8339 = uncached ? lru_94 : _GEN_6786; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8340 = uncached ? lru_95 : _GEN_6787; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8341 = uncached ? lru_96 : _GEN_6788; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8342 = uncached ? lru_97 : _GEN_6789; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8343 = uncached ? lru_98 : _GEN_6790; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8344 = uncached ? lru_99 : _GEN_6791; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8345 = uncached ? lru_100 : _GEN_6792; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8346 = uncached ? lru_101 : _GEN_6793; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8347 = uncached ? lru_102 : _GEN_6794; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8348 = uncached ? lru_103 : _GEN_6795; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8349 = uncached ? lru_104 : _GEN_6796; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8350 = uncached ? lru_105 : _GEN_6797; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8351 = uncached ? lru_106 : _GEN_6798; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8352 = uncached ? lru_107 : _GEN_6799; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8353 = uncached ? lru_108 : _GEN_6800; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8354 = uncached ? lru_109 : _GEN_6801; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8355 = uncached ? lru_110 : _GEN_6802; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8356 = uncached ? lru_111 : _GEN_6803; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8357 = uncached ? lru_112 : _GEN_6804; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8358 = uncached ? lru_113 : _GEN_6805; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8359 = uncached ? lru_114 : _GEN_6806; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8360 = uncached ? lru_115 : _GEN_6807; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8361 = uncached ? lru_116 : _GEN_6808; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8362 = uncached ? lru_117 : _GEN_6809; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8363 = uncached ? lru_118 : _GEN_6810; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8364 = uncached ? lru_119 : _GEN_6811; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8365 = uncached ? lru_120 : _GEN_6812; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8366 = uncached ? lru_121 : _GEN_6813; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8367 = uncached ? lru_122 : _GEN_6814; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8368 = uncached ? lru_123 : _GEN_6815; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8369 = uncached ? lru_124 : _GEN_6816; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8370 = uncached ? lru_125 : _GEN_6817; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8371 = uncached ? lru_126 : _GEN_6818; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8372 = uncached ? lru_127 : _GEN_6819; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8373 = uncached ? lru_128 : _GEN_6820; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8374 = uncached ? lru_129 : _GEN_6821; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8375 = uncached ? lru_130 : _GEN_6822; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8376 = uncached ? lru_131 : _GEN_6823; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8377 = uncached ? lru_132 : _GEN_6824; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8378 = uncached ? lru_133 : _GEN_6825; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8379 = uncached ? lru_134 : _GEN_6826; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8380 = uncached ? lru_135 : _GEN_6827; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8381 = uncached ? lru_136 : _GEN_6828; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8382 = uncached ? lru_137 : _GEN_6829; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8383 = uncached ? lru_138 : _GEN_6830; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8384 = uncached ? lru_139 : _GEN_6831; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8385 = uncached ? lru_140 : _GEN_6832; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8386 = uncached ? lru_141 : _GEN_6833; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8387 = uncached ? lru_142 : _GEN_6834; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8388 = uncached ? lru_143 : _GEN_6835; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8389 = uncached ? lru_144 : _GEN_6836; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8390 = uncached ? lru_145 : _GEN_6837; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8391 = uncached ? lru_146 : _GEN_6838; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8392 = uncached ? lru_147 : _GEN_6839; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8393 = uncached ? lru_148 : _GEN_6840; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8394 = uncached ? lru_149 : _GEN_6841; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8395 = uncached ? lru_150 : _GEN_6842; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8396 = uncached ? lru_151 : _GEN_6843; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8397 = uncached ? lru_152 : _GEN_6844; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8398 = uncached ? lru_153 : _GEN_6845; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8399 = uncached ? lru_154 : _GEN_6846; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8400 = uncached ? lru_155 : _GEN_6847; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8401 = uncached ? lru_156 : _GEN_6848; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8402 = uncached ? lru_157 : _GEN_6849; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8403 = uncached ? lru_158 : _GEN_6850; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8404 = uncached ? lru_159 : _GEN_6851; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8405 = uncached ? lru_160 : _GEN_6852; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8406 = uncached ? lru_161 : _GEN_6853; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8407 = uncached ? lru_162 : _GEN_6854; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8408 = uncached ? lru_163 : _GEN_6855; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8409 = uncached ? lru_164 : _GEN_6856; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8410 = uncached ? lru_165 : _GEN_6857; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8411 = uncached ? lru_166 : _GEN_6858; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8412 = uncached ? lru_167 : _GEN_6859; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8413 = uncached ? lru_168 : _GEN_6860; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8414 = uncached ? lru_169 : _GEN_6861; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8415 = uncached ? lru_170 : _GEN_6862; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8416 = uncached ? lru_171 : _GEN_6863; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8417 = uncached ? lru_172 : _GEN_6864; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8418 = uncached ? lru_173 : _GEN_6865; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8419 = uncached ? lru_174 : _GEN_6866; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8420 = uncached ? lru_175 : _GEN_6867; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8421 = uncached ? lru_176 : _GEN_6868; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8422 = uncached ? lru_177 : _GEN_6869; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8423 = uncached ? lru_178 : _GEN_6870; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8424 = uncached ? lru_179 : _GEN_6871; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8425 = uncached ? lru_180 : _GEN_6872; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8426 = uncached ? lru_181 : _GEN_6873; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8427 = uncached ? lru_182 : _GEN_6874; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8428 = uncached ? lru_183 : _GEN_6875; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8429 = uncached ? lru_184 : _GEN_6876; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8430 = uncached ? lru_185 : _GEN_6877; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8431 = uncached ? lru_186 : _GEN_6878; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8432 = uncached ? lru_187 : _GEN_6879; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8433 = uncached ? lru_188 : _GEN_6880; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8434 = uncached ? lru_189 : _GEN_6881; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8435 = uncached ? lru_190 : _GEN_6882; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8436 = uncached ? lru_191 : _GEN_6883; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8437 = uncached ? lru_192 : _GEN_6884; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8438 = uncached ? lru_193 : _GEN_6885; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8439 = uncached ? lru_194 : _GEN_6886; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8440 = uncached ? lru_195 : _GEN_6887; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8441 = uncached ? lru_196 : _GEN_6888; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8442 = uncached ? lru_197 : _GEN_6889; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8443 = uncached ? lru_198 : _GEN_6890; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8444 = uncached ? lru_199 : _GEN_6891; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8445 = uncached ? lru_200 : _GEN_6892; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8446 = uncached ? lru_201 : _GEN_6893; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8447 = uncached ? lru_202 : _GEN_6894; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8448 = uncached ? lru_203 : _GEN_6895; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8449 = uncached ? lru_204 : _GEN_6896; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8450 = uncached ? lru_205 : _GEN_6897; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8451 = uncached ? lru_206 : _GEN_6898; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8452 = uncached ? lru_207 : _GEN_6899; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8453 = uncached ? lru_208 : _GEN_6900; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8454 = uncached ? lru_209 : _GEN_6901; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8455 = uncached ? lru_210 : _GEN_6902; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8456 = uncached ? lru_211 : _GEN_6903; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8457 = uncached ? lru_212 : _GEN_6904; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8458 = uncached ? lru_213 : _GEN_6905; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8459 = uncached ? lru_214 : _GEN_6906; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8460 = uncached ? lru_215 : _GEN_6907; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8461 = uncached ? lru_216 : _GEN_6908; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8462 = uncached ? lru_217 : _GEN_6909; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8463 = uncached ? lru_218 : _GEN_6910; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8464 = uncached ? lru_219 : _GEN_6911; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8465 = uncached ? lru_220 : _GEN_6912; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8466 = uncached ? lru_221 : _GEN_6913; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8467 = uncached ? lru_222 : _GEN_6914; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8468 = uncached ? lru_223 : _GEN_6915; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8469 = uncached ? lru_224 : _GEN_6916; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8470 = uncached ? lru_225 : _GEN_6917; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8471 = uncached ? lru_226 : _GEN_6918; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8472 = uncached ? lru_227 : _GEN_6919; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8473 = uncached ? lru_228 : _GEN_6920; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8474 = uncached ? lru_229 : _GEN_6921; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8475 = uncached ? lru_230 : _GEN_6922; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8476 = uncached ? lru_231 : _GEN_6923; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8477 = uncached ? lru_232 : _GEN_6924; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8478 = uncached ? lru_233 : _GEN_6925; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8479 = uncached ? lru_234 : _GEN_6926; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8480 = uncached ? lru_235 : _GEN_6927; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8481 = uncached ? lru_236 : _GEN_6928; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8482 = uncached ? lru_237 : _GEN_6929; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8483 = uncached ? lru_238 : _GEN_6930; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8484 = uncached ? lru_239 : _GEN_6931; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8485 = uncached ? lru_240 : _GEN_6932; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8486 = uncached ? lru_241 : _GEN_6933; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8487 = uncached ? lru_242 : _GEN_6934; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8488 = uncached ? lru_243 : _GEN_6935; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8489 = uncached ? lru_244 : _GEN_6936; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8490 = uncached ? lru_245 : _GEN_6937; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8491 = uncached ? lru_246 : _GEN_6938; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8492 = uncached ? lru_247 : _GEN_6939; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8493 = uncached ? lru_248 : _GEN_6940; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8494 = uncached ? lru_249 : _GEN_6941; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8495 = uncached ? lru_250 : _GEN_6942; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8496 = uncached ? lru_251 : _GEN_6943; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8497 = uncached ? lru_252 : _GEN_6944; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8498 = uncached ? lru_253 : _GEN_6945; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8499 = uncached ? lru_254 : _GEN_6946; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8500 = uncached ? lru_255 : _GEN_6947; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8501 = uncached ? lru_256 : _GEN_6948; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8502 = uncached ? lru_257 : _GEN_6949; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8503 = uncached ? lru_258 : _GEN_6950; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8504 = uncached ? lru_259 : _GEN_6951; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8505 = uncached ? lru_260 : _GEN_6952; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8506 = uncached ? lru_261 : _GEN_6953; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8507 = uncached ? lru_262 : _GEN_6954; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8508 = uncached ? lru_263 : _GEN_6955; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8509 = uncached ? lru_264 : _GEN_6956; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8510 = uncached ? lru_265 : _GEN_6957; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8511 = uncached ? lru_266 : _GEN_6958; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8512 = uncached ? lru_267 : _GEN_6959; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8513 = uncached ? lru_268 : _GEN_6960; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8514 = uncached ? lru_269 : _GEN_6961; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8515 = uncached ? lru_270 : _GEN_6962; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8516 = uncached ? lru_271 : _GEN_6963; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8517 = uncached ? lru_272 : _GEN_6964; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8518 = uncached ? lru_273 : _GEN_6965; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8519 = uncached ? lru_274 : _GEN_6966; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8520 = uncached ? lru_275 : _GEN_6967; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8521 = uncached ? lru_276 : _GEN_6968; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8522 = uncached ? lru_277 : _GEN_6969; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8523 = uncached ? lru_278 : _GEN_6970; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8524 = uncached ? lru_279 : _GEN_6971; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8525 = uncached ? lru_280 : _GEN_6972; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8526 = uncached ? lru_281 : _GEN_6973; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8527 = uncached ? lru_282 : _GEN_6974; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8528 = uncached ? lru_283 : _GEN_6975; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8529 = uncached ? lru_284 : _GEN_6976; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8530 = uncached ? lru_285 : _GEN_6977; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8531 = uncached ? lru_286 : _GEN_6978; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8532 = uncached ? lru_287 : _GEN_6979; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8533 = uncached ? lru_288 : _GEN_6980; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8534 = uncached ? lru_289 : _GEN_6981; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8535 = uncached ? lru_290 : _GEN_6982; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8536 = uncached ? lru_291 : _GEN_6983; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8537 = uncached ? lru_292 : _GEN_6984; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8538 = uncached ? lru_293 : _GEN_6985; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8539 = uncached ? lru_294 : _GEN_6986; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8540 = uncached ? lru_295 : _GEN_6987; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8541 = uncached ? lru_296 : _GEN_6988; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8542 = uncached ? lru_297 : _GEN_6989; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8543 = uncached ? lru_298 : _GEN_6990; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8544 = uncached ? lru_299 : _GEN_6991; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8545 = uncached ? lru_300 : _GEN_6992; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8546 = uncached ? lru_301 : _GEN_6993; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8547 = uncached ? lru_302 : _GEN_6994; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8548 = uncached ? lru_303 : _GEN_6995; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8549 = uncached ? lru_304 : _GEN_6996; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8550 = uncached ? lru_305 : _GEN_6997; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8551 = uncached ? lru_306 : _GEN_6998; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8552 = uncached ? lru_307 : _GEN_6999; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8553 = uncached ? lru_308 : _GEN_7000; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8554 = uncached ? lru_309 : _GEN_7001; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8555 = uncached ? lru_310 : _GEN_7002; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8556 = uncached ? lru_311 : _GEN_7003; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8557 = uncached ? lru_312 : _GEN_7004; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8558 = uncached ? lru_313 : _GEN_7005; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8559 = uncached ? lru_314 : _GEN_7006; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8560 = uncached ? lru_315 : _GEN_7007; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8561 = uncached ? lru_316 : _GEN_7008; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8562 = uncached ? lru_317 : _GEN_7009; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8563 = uncached ? lru_318 : _GEN_7010; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8564 = uncached ? lru_319 : _GEN_7011; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8565 = uncached ? lru_320 : _GEN_7012; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8566 = uncached ? lru_321 : _GEN_7013; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8567 = uncached ? lru_322 : _GEN_7014; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8568 = uncached ? lru_323 : _GEN_7015; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8569 = uncached ? lru_324 : _GEN_7016; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8570 = uncached ? lru_325 : _GEN_7017; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8571 = uncached ? lru_326 : _GEN_7018; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8572 = uncached ? lru_327 : _GEN_7019; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8573 = uncached ? lru_328 : _GEN_7020; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8574 = uncached ? lru_329 : _GEN_7021; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8575 = uncached ? lru_330 : _GEN_7022; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8576 = uncached ? lru_331 : _GEN_7023; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8577 = uncached ? lru_332 : _GEN_7024; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8578 = uncached ? lru_333 : _GEN_7025; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8579 = uncached ? lru_334 : _GEN_7026; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8580 = uncached ? lru_335 : _GEN_7027; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8581 = uncached ? lru_336 : _GEN_7028; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8582 = uncached ? lru_337 : _GEN_7029; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8583 = uncached ? lru_338 : _GEN_7030; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8584 = uncached ? lru_339 : _GEN_7031; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8585 = uncached ? lru_340 : _GEN_7032; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8586 = uncached ? lru_341 : _GEN_7033; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8587 = uncached ? lru_342 : _GEN_7034; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8588 = uncached ? lru_343 : _GEN_7035; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8589 = uncached ? lru_344 : _GEN_7036; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8590 = uncached ? lru_345 : _GEN_7037; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8591 = uncached ? lru_346 : _GEN_7038; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8592 = uncached ? lru_347 : _GEN_7039; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8593 = uncached ? lru_348 : _GEN_7040; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8594 = uncached ? lru_349 : _GEN_7041; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8595 = uncached ? lru_350 : _GEN_7042; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8596 = uncached ? lru_351 : _GEN_7043; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8597 = uncached ? lru_352 : _GEN_7044; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8598 = uncached ? lru_353 : _GEN_7045; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8599 = uncached ? lru_354 : _GEN_7046; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8600 = uncached ? lru_355 : _GEN_7047; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8601 = uncached ? lru_356 : _GEN_7048; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8602 = uncached ? lru_357 : _GEN_7049; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8603 = uncached ? lru_358 : _GEN_7050; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8604 = uncached ? lru_359 : _GEN_7051; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8605 = uncached ? lru_360 : _GEN_7052; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8606 = uncached ? lru_361 : _GEN_7053; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8607 = uncached ? lru_362 : _GEN_7054; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8608 = uncached ? lru_363 : _GEN_7055; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8609 = uncached ? lru_364 : _GEN_7056; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8610 = uncached ? lru_365 : _GEN_7057; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8611 = uncached ? lru_366 : _GEN_7058; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8612 = uncached ? lru_367 : _GEN_7059; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8613 = uncached ? lru_368 : _GEN_7060; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8614 = uncached ? lru_369 : _GEN_7061; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8615 = uncached ? lru_370 : _GEN_7062; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8616 = uncached ? lru_371 : _GEN_7063; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8617 = uncached ? lru_372 : _GEN_7064; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8618 = uncached ? lru_373 : _GEN_7065; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8619 = uncached ? lru_374 : _GEN_7066; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8620 = uncached ? lru_375 : _GEN_7067; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8621 = uncached ? lru_376 : _GEN_7068; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8622 = uncached ? lru_377 : _GEN_7069; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8623 = uncached ? lru_378 : _GEN_7070; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8624 = uncached ? lru_379 : _GEN_7071; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8625 = uncached ? lru_380 : _GEN_7072; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8626 = uncached ? lru_381 : _GEN_7073; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8627 = uncached ? lru_382 : _GEN_7074; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8628 = uncached ? lru_383 : _GEN_7075; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8629 = uncached ? lru_384 : _GEN_7076; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8630 = uncached ? lru_385 : _GEN_7077; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8631 = uncached ? lru_386 : _GEN_7078; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8632 = uncached ? lru_387 : _GEN_7079; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8633 = uncached ? lru_388 : _GEN_7080; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8634 = uncached ? lru_389 : _GEN_7081; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8635 = uncached ? lru_390 : _GEN_7082; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8636 = uncached ? lru_391 : _GEN_7083; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8637 = uncached ? lru_392 : _GEN_7084; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8638 = uncached ? lru_393 : _GEN_7085; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8639 = uncached ? lru_394 : _GEN_7086; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8640 = uncached ? lru_395 : _GEN_7087; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8641 = uncached ? lru_396 : _GEN_7088; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8642 = uncached ? lru_397 : _GEN_7089; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8643 = uncached ? lru_398 : _GEN_7090; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8644 = uncached ? lru_399 : _GEN_7091; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8645 = uncached ? lru_400 : _GEN_7092; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8646 = uncached ? lru_401 : _GEN_7093; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8647 = uncached ? lru_402 : _GEN_7094; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8648 = uncached ? lru_403 : _GEN_7095; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8649 = uncached ? lru_404 : _GEN_7096; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8650 = uncached ? lru_405 : _GEN_7097; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8651 = uncached ? lru_406 : _GEN_7098; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8652 = uncached ? lru_407 : _GEN_7099; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8653 = uncached ? lru_408 : _GEN_7100; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8654 = uncached ? lru_409 : _GEN_7101; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8655 = uncached ? lru_410 : _GEN_7102; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8656 = uncached ? lru_411 : _GEN_7103; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8657 = uncached ? lru_412 : _GEN_7104; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8658 = uncached ? lru_413 : _GEN_7105; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8659 = uncached ? lru_414 : _GEN_7106; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8660 = uncached ? lru_415 : _GEN_7107; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8661 = uncached ? lru_416 : _GEN_7108; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8662 = uncached ? lru_417 : _GEN_7109; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8663 = uncached ? lru_418 : _GEN_7110; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8664 = uncached ? lru_419 : _GEN_7111; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8665 = uncached ? lru_420 : _GEN_7112; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8666 = uncached ? lru_421 : _GEN_7113; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8667 = uncached ? lru_422 : _GEN_7114; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8668 = uncached ? lru_423 : _GEN_7115; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8669 = uncached ? lru_424 : _GEN_7116; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8670 = uncached ? lru_425 : _GEN_7117; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8671 = uncached ? lru_426 : _GEN_7118; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8672 = uncached ? lru_427 : _GEN_7119; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8673 = uncached ? lru_428 : _GEN_7120; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8674 = uncached ? lru_429 : _GEN_7121; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8675 = uncached ? lru_430 : _GEN_7122; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8676 = uncached ? lru_431 : _GEN_7123; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8677 = uncached ? lru_432 : _GEN_7124; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8678 = uncached ? lru_433 : _GEN_7125; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8679 = uncached ? lru_434 : _GEN_7126; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8680 = uncached ? lru_435 : _GEN_7127; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8681 = uncached ? lru_436 : _GEN_7128; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8682 = uncached ? lru_437 : _GEN_7129; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8683 = uncached ? lru_438 : _GEN_7130; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8684 = uncached ? lru_439 : _GEN_7131; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8685 = uncached ? lru_440 : _GEN_7132; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8686 = uncached ? lru_441 : _GEN_7133; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8687 = uncached ? lru_442 : _GEN_7134; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8688 = uncached ? lru_443 : _GEN_7135; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8689 = uncached ? lru_444 : _GEN_7136; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8690 = uncached ? lru_445 : _GEN_7137; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8691 = uncached ? lru_446 : _GEN_7138; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8692 = uncached ? lru_447 : _GEN_7139; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8693 = uncached ? lru_448 : _GEN_7140; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8694 = uncached ? lru_449 : _GEN_7141; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8695 = uncached ? lru_450 : _GEN_7142; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8696 = uncached ? lru_451 : _GEN_7143; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8697 = uncached ? lru_452 : _GEN_7144; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8698 = uncached ? lru_453 : _GEN_7145; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8699 = uncached ? lru_454 : _GEN_7146; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8700 = uncached ? lru_455 : _GEN_7147; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8701 = uncached ? lru_456 : _GEN_7148; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8702 = uncached ? lru_457 : _GEN_7149; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8703 = uncached ? lru_458 : _GEN_7150; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8704 = uncached ? lru_459 : _GEN_7151; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8705 = uncached ? lru_460 : _GEN_7152; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8706 = uncached ? lru_461 : _GEN_7153; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8707 = uncached ? lru_462 : _GEN_7154; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8708 = uncached ? lru_463 : _GEN_7155; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8709 = uncached ? lru_464 : _GEN_7156; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8710 = uncached ? lru_465 : _GEN_7157; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8711 = uncached ? lru_466 : _GEN_7158; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8712 = uncached ? lru_467 : _GEN_7159; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8713 = uncached ? lru_468 : _GEN_7160; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8714 = uncached ? lru_469 : _GEN_7161; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8715 = uncached ? lru_470 : _GEN_7162; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8716 = uncached ? lru_471 : _GEN_7163; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8717 = uncached ? lru_472 : _GEN_7164; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8718 = uncached ? lru_473 : _GEN_7165; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8719 = uncached ? lru_474 : _GEN_7166; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8720 = uncached ? lru_475 : _GEN_7167; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8721 = uncached ? lru_476 : _GEN_7168; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8722 = uncached ? lru_477 : _GEN_7169; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8723 = uncached ? lru_478 : _GEN_7170; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8724 = uncached ? lru_479 : _GEN_7171; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8725 = uncached ? lru_480 : _GEN_7172; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8726 = uncached ? lru_481 : _GEN_7173; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8727 = uncached ? lru_482 : _GEN_7174; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8728 = uncached ? lru_483 : _GEN_7175; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8729 = uncached ? lru_484 : _GEN_7176; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8730 = uncached ? lru_485 : _GEN_7177; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8731 = uncached ? lru_486 : _GEN_7178; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8732 = uncached ? lru_487 : _GEN_7179; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8733 = uncached ? lru_488 : _GEN_7180; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8734 = uncached ? lru_489 : _GEN_7181; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8735 = uncached ? lru_490 : _GEN_7182; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8736 = uncached ? lru_491 : _GEN_7183; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8737 = uncached ? lru_492 : _GEN_7184; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8738 = uncached ? lru_493 : _GEN_7185; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8739 = uncached ? lru_494 : _GEN_7186; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8740 = uncached ? lru_495 : _GEN_7187; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8741 = uncached ? lru_496 : _GEN_7188; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8742 = uncached ? lru_497 : _GEN_7189; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8743 = uncached ? lru_498 : _GEN_7190; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8744 = uncached ? lru_499 : _GEN_7191; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8745 = uncached ? lru_500 : _GEN_7192; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8746 = uncached ? lru_501 : _GEN_7193; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8747 = uncached ? lru_502 : _GEN_7194; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8748 = uncached ? lru_503 : _GEN_7195; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8749 = uncached ? lru_504 : _GEN_7196; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8750 = uncached ? lru_505 : _GEN_7197; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8751 = uncached ? lru_506 : _GEN_7198; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8752 = uncached ? lru_507 : _GEN_7199; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8753 = uncached ? lru_508 : _GEN_7200; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8754 = uncached ? lru_509 : _GEN_7201; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8755 = uncached ? lru_510 : _GEN_7202; // @[ICache.scala 169:30 68:20]
  wire  _GEN_8756 = uncached ? lru_511 : _GEN_7203; // @[ICache.scala 169:30 68:20]
  wire [31:0] _GEN_8757 = uncached ? saved_1_inst : _GEN_7204; // @[ICache.scala 113:22 169:30]
  wire  _GEN_8758 = uncached ? saved_0_valid : _GEN_7205; // @[ICache.scala 113:22 169:30]
  wire  _GEN_8759 = uncached ? saved_1_valid : _GEN_7206; // @[ICache.scala 113:22 169:30]
  wire [19:0] _GEN_11867 = inst_vpn[12] ? io_cpu_tlb2_entry_pfn_1 : io_cpu_tlb2_entry_pfn_0; // @[ICache.scala 204:{22,22}]
  wire  _GEN_11869 = inst_vpn[12] ? io_cpu_tlb2_entry_c_1 : io_cpu_tlb2_entry_c_0; // @[ICache.scala 205:{22,22}]
  wire  _GEN_11874 = io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_v_1 | ~inst_vpn[12] & io_cpu_tlb2_entry_v_0)
     | _GEN_2; // @[ICache.scala 201:118 206:22]
  wire  _GEN_11878 = io_axi_ar_ready ? 1'h0 : arvalid; // @[ICache.scala 216:31 217:19 150:24]
  wire  _GEN_11879 = io_axi_ar_ready | rready; // @[ICache.scala 216:31 218:19 155:23]
  wire  _T_21 = io_axi_r_ready & io_axi_r_valid; // @[Decoupled.scala 52:35]
  wire [2:0] _GEN_11880 = _T_21 ? 3'h4 : state; // @[ICache.scala 220:33 221:24 39:81]
  wire [31:0] _GEN_11881 = _T_21 ? io_axi_r_bits_data : saved_0_inst; // @[ICache.scala 113:22 220:33 222:24]
  wire  _GEN_11882 = _T_21 | saved_0_valid; // @[ICache.scala 113:22 220:33 223:24]
  wire  _GEN_11883 = _T_21 ? 1'h0 : rready; // @[ICache.scala 155:23 220:33 224:24]
  wire  _GEN_11884 = io_axi_ar_valid ? _GEN_11878 : arvalid; // @[ICache.scala 150:24 215:29]
  wire  _GEN_11885 = io_axi_ar_valid ? _GEN_11879 : _GEN_11883; // @[ICache.scala 215:29]
  wire [2:0] _GEN_11886 = io_axi_ar_valid ? state : _GEN_11880; // @[ICache.scala 215:29 39:81]
  wire [31:0] _GEN_11887 = io_axi_ar_valid ? saved_0_inst : _GEN_11881; // @[ICache.scala 113:22 215:29]
  wire  _GEN_11888 = io_axi_ar_valid ? saved_0_valid : _GEN_11882; // @[ICache.scala 113:22 215:29]
  wire [4:0] _value_T_1 = axi_cnt_value + 5'h1; // @[Counter.scala 77:24]
  wire [3:0] _GEN_11890 = _GEN_3591 ? data_wstrb_1_0 : data_wstrb_0_0; // @[ICache.scala 236:{39,39}]
  wire [3:0] _data_wstrb_0_T = ~_GEN_11890; // @[ICache.scala 236:39]
  wire [3:0] _GEN_11891 = ~_GEN_3591 ? _data_wstrb_0_T : data_wstrb_0_0; // @[ICache.scala 236:{36,36} 61:27]
  wire [3:0] _GEN_11892 = _GEN_3591 ? _data_wstrb_0_T : data_wstrb_1_0; // @[ICache.scala 236:{36,36} 61:27]
  wire [3:0] _GEN_11894 = _GEN_3591 ? data_wstrb_1_1 : data_wstrb_0_1; // @[ICache.scala 237:{39,39}]
  wire [3:0] _data_wstrb_1_T = ~_GEN_11894; // @[ICache.scala 237:39]
  wire [3:0] _GEN_11895 = ~_GEN_3591 ? _data_wstrb_1_T : data_wstrb_0_1; // @[ICache.scala 237:{36,36} 61:27]
  wire [3:0] _GEN_11896 = _GEN_3591 ? _data_wstrb_1_T : data_wstrb_1_1; // @[ICache.scala 237:{36,36} 61:27]
  wire [3:0] _GEN_11897 = ~_GEN_3591 ? 4'h0 : data_wstrb_0_0; // @[ICache.scala 240:{33,33} 61:27]
  wire [3:0] _GEN_11898 = _GEN_3591 ? 4'h0 : data_wstrb_1_0; // @[ICache.scala 240:{33,33} 61:27]
  wire  _GEN_11901 = ~_GEN_3591 ? 1'h0 : tag_wstrb_0; // @[ICache.scala 241:{33,33} 64:26]
  wire  _GEN_11902 = _GEN_3591 ? 1'h0 : tag_wstrb_1; // @[ICache.scala 241:{33,33} 64:26]
  wire [4:0] _GEN_11903 = ~io_axi_r_bits_last ? _value_T_1 : axi_cnt_value; // @[ICache.scala 234:35 Counter.scala 77:15 61:40]
  wire [3:0] _GEN_11904 = ~io_axi_r_bits_last ? _GEN_11891 : _GEN_11897; // @[ICache.scala 234:35]
  wire [3:0] _GEN_11905 = ~io_axi_r_bits_last ? _GEN_11892 : _GEN_11898; // @[ICache.scala 234:35]
  wire [3:0] _GEN_11906 = ~io_axi_r_bits_last ? _GEN_11895 : _GEN_3594; // @[ICache.scala 234:35]
  wire [3:0] _GEN_11907 = ~io_axi_r_bits_last ? _GEN_11896 : _GEN_3595; // @[ICache.scala 234:35]
  wire  _GEN_11908 = ~io_axi_r_bits_last & rready; // @[ICache.scala 155:23 234:35 239:33]
  wire  _GEN_11909 = ~io_axi_r_bits_last ? tag_wstrb_0 : _GEN_11901; // @[ICache.scala 234:35 64:26]
  wire  _GEN_11910 = ~io_axi_r_bits_last ? tag_wstrb_1 : _GEN_11902; // @[ICache.scala 234:35 64:26]
  wire [2:0] _GEN_11911 = ~io_axi_r_ready ? 3'h0 : state; // @[ICache.scala 243:35 244:15 39:81]
  wire [4:0] _GEN_11912 = _T_21 ? _GEN_11903 : axi_cnt_value; // @[ICache.scala 233:33 Counter.scala 61:40]
  wire [3:0] _GEN_11913 = _T_21 ? _GEN_11904 : data_wstrb_0_0; // @[ICache.scala 233:33 61:27]
  wire [3:0] _GEN_11914 = _T_21 ? _GEN_11905 : data_wstrb_1_0; // @[ICache.scala 233:33 61:27]
  wire [3:0] _GEN_11915 = _T_21 ? _GEN_11906 : data_wstrb_0_1; // @[ICache.scala 233:33 61:27]
  wire [3:0] _GEN_11916 = _T_21 ? _GEN_11907 : data_wstrb_1_1; // @[ICache.scala 233:33 61:27]
  wire  _GEN_11917 = _T_21 ? _GEN_11908 : rready; // @[ICache.scala 155:23 233:33]
  wire  _GEN_11918 = _T_21 ? _GEN_11909 : tag_wstrb_0; // @[ICache.scala 233:33 64:26]
  wire  _GEN_11919 = _T_21 ? _GEN_11910 : tag_wstrb_1; // @[ICache.scala 233:33 64:26]
  wire [2:0] _GEN_11920 = _T_21 ? state : _GEN_11911; // @[ICache.scala 233:33 39:81]
  wire  _GEN_11921 = io_axi_ar_valid ? _GEN_11879 : _GEN_11917; // @[ICache.scala 228:29]
  wire [4:0] _GEN_11922 = io_axi_ar_valid ? axi_cnt_value : _GEN_11912; // @[ICache.scala 228:29 Counter.scala 61:40]
  wire [3:0] _GEN_11923 = io_axi_ar_valid ? data_wstrb_0_0 : _GEN_11913; // @[ICache.scala 228:29 61:27]
  wire [3:0] _GEN_11924 = io_axi_ar_valid ? data_wstrb_1_0 : _GEN_11914; // @[ICache.scala 228:29 61:27]
  wire [3:0] _GEN_11925 = io_axi_ar_valid ? data_wstrb_0_1 : _GEN_11915; // @[ICache.scala 228:29 61:27]
  wire [3:0] _GEN_11926 = io_axi_ar_valid ? data_wstrb_1_1 : _GEN_11916; // @[ICache.scala 228:29 61:27]
  wire  _GEN_11927 = io_axi_ar_valid ? tag_wstrb_0 : _GEN_11918; // @[ICache.scala 228:29 64:26]
  wire  _GEN_11928 = io_axi_ar_valid ? tag_wstrb_1 : _GEN_11919; // @[ICache.scala 228:29 64:26]
  wire [2:0] _GEN_11929 = io_axi_ar_valid ? state : _GEN_11920; // @[ICache.scala 228:29 39:81]
  wire [2:0] _GEN_11930 = _T_2 & _T ? 3'h0 : state; // @[ICache.scala 248:55 249:24 39:81]
  wire  _GEN_11931 = _T_2 & _T ? 1'h0 : tlb1_invalid; // @[ICache.scala 248:55 250:24 159:29]
  wire  _GEN_11932 = _T_2 & _T ? 1'h0 : saved_0_valid; // @[ICache.scala 113:22 248:55 251:24]
  wire  _GEN_11933 = _T_2 & _T ? 1'h0 : saved_1_valid; // @[ICache.scala 113:22 248:55 252:24]
  wire [2:0] _GEN_11934 = 3'h4 == state ? _GEN_11930 : state; // @[ICache.scala 164:17 39:81]
  wire  _GEN_11935 = 3'h4 == state ? _GEN_11931 : tlb1_invalid; // @[ICache.scala 164:17 159:29]
  wire  _GEN_11936 = 3'h4 == state ? _GEN_11932 : saved_0_valid; // @[ICache.scala 164:17 113:22]
  wire  _GEN_11937 = 3'h4 == state ? _GEN_11933 : saved_1_valid; // @[ICache.scala 164:17 113:22]
  wire  _GEN_11938 = 3'h3 == state ? _GEN_11884 : arvalid; // @[ICache.scala 164:17 150:24]
  wire  _GEN_11939 = 3'h3 == state ? _GEN_11921 : rready; // @[ICache.scala 164:17 155:23]
  wire [4:0] _GEN_11940 = 3'h3 == state ? _GEN_11922 : axi_cnt_value; // @[ICache.scala 164:17 Counter.scala 61:40]
  wire [3:0] _GEN_11941 = 3'h3 == state ? _GEN_11923 : data_wstrb_0_0; // @[ICache.scala 164:17 61:27]
  wire [3:0] _GEN_11942 = 3'h3 == state ? _GEN_11924 : data_wstrb_1_0; // @[ICache.scala 164:17 61:27]
  wire [3:0] _GEN_11943 = 3'h3 == state ? _GEN_11925 : data_wstrb_0_1; // @[ICache.scala 164:17 61:27]
  wire [3:0] _GEN_11944 = 3'h3 == state ? _GEN_11926 : data_wstrb_1_1; // @[ICache.scala 164:17 61:27]
  wire  _GEN_11945 = 3'h3 == state ? _GEN_11927 : tag_wstrb_0; // @[ICache.scala 164:17 64:26]
  wire  _GEN_11946 = 3'h3 == state ? _GEN_11928 : tag_wstrb_1; // @[ICache.scala 164:17 64:26]
  wire [2:0] _GEN_11947 = 3'h3 == state ? _GEN_11929 : _GEN_11934; // @[ICache.scala 164:17]
  wire  _GEN_11948 = 3'h3 == state ? tlb1_invalid : _GEN_11935; // @[ICache.scala 164:17 159:29]
  wire  _GEN_11949 = 3'h3 == state ? saved_0_valid : _GEN_11936; // @[ICache.scala 164:17 113:22]
  wire  _GEN_11950 = 3'h3 == state ? saved_1_valid : _GEN_11937; // @[ICache.scala 164:17 113:22]
  SimpleDualPortRam bank ( // @[ICache.scala 122:22]
    .clock(bank_clock),
    .reset(bank_reset),
    .io_raddr(bank_io_raddr),
    .io_rdata(bank_io_rdata),
    .io_waddr(bank_io_waddr),
    .io_wen(bank_io_wen),
    .io_wstrb(bank_io_wstrb),
    .io_wdata(bank_io_wdata)
  );
  SimpleDualPortRam_1 tag_bram ( // @[ICache.scala 132:26]
    .clock(tag_bram_clock),
    .reset(tag_bram_reset),
    .io_raddr(tag_bram_io_raddr),
    .io_rdata(tag_bram_io_rdata),
    .io_waddr(tag_bram_io_waddr),
    .io_wen(tag_bram_io_wen),
    .io_wstrb(tag_bram_io_wstrb),
    .io_wdata(tag_bram_io_wdata)
  );
  SimpleDualPortRam bank_1 ( // @[ICache.scala 122:22]
    .clock(bank_1_clock),
    .reset(bank_1_reset),
    .io_raddr(bank_1_io_raddr),
    .io_rdata(bank_1_io_rdata),
    .io_waddr(bank_1_io_waddr),
    .io_wen(bank_1_io_wen),
    .io_wstrb(bank_1_io_wstrb),
    .io_wdata(bank_1_io_wdata)
  );
  SimpleDualPortRam_1 tag_bram_1 ( // @[ICache.scala 132:26]
    .clock(tag_bram_1_clock),
    .reset(tag_bram_1_reset),
    .io_raddr(tag_bram_1_io_raddr),
    .io_rdata(tag_bram_1_io_rdata),
    .io_waddr(tag_bram_1_io_waddr),
    .io_wen(tag_bram_1_io_wen),
    .io_wstrb(tag_bram_1_io_wstrb),
    .io_wdata(tag_bram_1_io_wdata)
  );
  SimpleDualPortRam bank_2 ( // @[ICache.scala 122:22]
    .clock(bank_2_clock),
    .reset(bank_2_reset),
    .io_raddr(bank_2_io_raddr),
    .io_rdata(bank_2_io_rdata),
    .io_waddr(bank_2_io_waddr),
    .io_wen(bank_2_io_wen),
    .io_wstrb(bank_2_io_wstrb),
    .io_wdata(bank_2_io_wdata)
  );
  SimpleDualPortRam_1 tag_bram_2 ( // @[ICache.scala 132:26]
    .clock(tag_bram_2_clock),
    .reset(tag_bram_2_reset),
    .io_raddr(tag_bram_2_io_raddr),
    .io_rdata(tag_bram_2_io_rdata),
    .io_waddr(tag_bram_2_io_waddr),
    .io_wen(tag_bram_2_io_wen),
    .io_wstrb(tag_bram_2_io_wstrb),
    .io_wdata(tag_bram_2_io_wdata)
  );
  SimpleDualPortRam bank_3 ( // @[ICache.scala 122:22]
    .clock(bank_3_clock),
    .reset(bank_3_reset),
    .io_raddr(bank_3_io_raddr),
    .io_rdata(bank_3_io_rdata),
    .io_waddr(bank_3_io_waddr),
    .io_wen(bank_3_io_wen),
    .io_wstrb(bank_3_io_wstrb),
    .io_wdata(bank_3_io_wdata)
  );
  SimpleDualPortRam_1 tag_bram_3 ( // @[ICache.scala 132:26]
    .clock(tag_bram_3_clock),
    .reset(tag_bram_3_reset),
    .io_raddr(tag_bram_3_io_raddr),
    .io_rdata(tag_bram_3_io_rdata),
    .io_waddr(tag_bram_3_io_waddr),
    .io_wen(tag_bram_3_io_wen),
    .io_wstrb(tag_bram_3_io_wstrb),
    .io_wdata(tag_bram_3_io_wdata)
  );
  assign io_cpu_inst_0 = _should_next_addr_T ? inst_0 : saved_0_inst; // @[ICache.scala 143:32]
  assign io_cpu_inst_1 = _should_next_addr_T ? inst_1 : saved_1_inst; // @[ICache.scala 143:32]
  assign io_cpu_inst_valid_0 = _io_cpu_inst_valid_0_T_4 & io_cpu_req; // @[ICache.scala 142:82]
  assign io_cpu_inst_valid_1 = _io_cpu_inst_valid_1_T_4 & io_cpu_req; // @[ICache.scala 142:82]
  assign io_cpu_icache_stall = _should_next_addr_T ? ~cache_hit_available & io_cpu_req : state != 3'h4; // @[ICache.scala 147:29]
  assign io_cpu_tlb1_invalid = tlb1_invalid; // @[ICache.scala 160:23]
  assign io_cpu_tlb2_vpn = io_cpu_tlb2_vpn_r[18:0]; // @[ICache.scala 162:19]
  assign io_axi_ar_valid = arvalid; // @[ICache.scala 152:11]
  assign io_axi_ar_bits_addr = ar_addr; // @[ICache.scala 151:6]
  assign io_axi_ar_bits_len = ar_len; // @[ICache.scala 151:6]
  assign io_axi_ar_bits_size = ar_size; // @[ICache.scala 151:6]
  assign io_axi_r_ready = rready; // @[ICache.scala 157:10]
  assign bank_clock = clock;
  assign bank_reset = reset;
  assign bank_io_raddr = _GEN_1[11:3]; // @[ICache.scala 60:49]
  assign bank_io_waddr = {rset,axi_cnt_value[3:1]}; // @[Cat.scala 33:92]
  assign bank_io_wen = |data_wstrb_0_0; // @[ICache.scala 127:39]
  assign bank_io_wstrb = data_wstrb_0_0; // @[ICache.scala 130:19]
  assign bank_io_wdata = ~axi_cnt_value[0] ? io_axi_r_bits_data : 32'h0; // @[ICache.scala 129:25]
  assign tag_bram_clock = clock;
  assign tag_bram_reset = reset;
  assign tag_bram_io_raddr = _GEN_1[11:6]; // @[ICache.scala 63:48]
  assign tag_bram_io_waddr = rset; // @[ICache.scala 138:23]
  assign tag_bram_io_wen = |tag_wstrb_0; // @[ICache.scala 137:39]
  assign tag_bram_io_wstrb = tag_wstrb_0; // @[ICache.scala 140:23]
  assign tag_bram_io_wdata = tag_wdata; // @[ICache.scala 139:23]
  assign bank_1_clock = clock;
  assign bank_1_reset = reset;
  assign bank_1_io_raddr = _GEN_1[11:3]; // @[ICache.scala 60:49]
  assign bank_1_io_waddr = {rset,axi_cnt_value[3:1]}; // @[Cat.scala 33:92]
  assign bank_1_io_wen = |data_wstrb_0_1; // @[ICache.scala 127:39]
  assign bank_1_io_wstrb = data_wstrb_0_1; // @[ICache.scala 130:19]
  assign bank_1_io_wdata = axi_cnt_value[0] ? io_axi_r_bits_data : 32'h0; // @[ICache.scala 129:25]
  assign tag_bram_1_clock = clock;
  assign tag_bram_1_reset = reset;
  assign tag_bram_1_io_raddr = _GEN_1[11:6]; // @[ICache.scala 63:48]
  assign tag_bram_1_io_waddr = rset; // @[ICache.scala 138:23]
  assign tag_bram_1_io_wen = |tag_wstrb_0; // @[ICache.scala 137:39]
  assign tag_bram_1_io_wstrb = tag_wstrb_0; // @[ICache.scala 140:23]
  assign tag_bram_1_io_wdata = tag_wdata; // @[ICache.scala 139:23]
  assign bank_2_clock = clock;
  assign bank_2_reset = reset;
  assign bank_2_io_raddr = _GEN_1[11:3]; // @[ICache.scala 60:49]
  assign bank_2_io_waddr = {rset,axi_cnt_value[3:1]}; // @[Cat.scala 33:92]
  assign bank_2_io_wen = |data_wstrb_1_0; // @[ICache.scala 127:39]
  assign bank_2_io_wstrb = data_wstrb_1_0; // @[ICache.scala 130:19]
  assign bank_2_io_wdata = ~axi_cnt_value[0] ? io_axi_r_bits_data : 32'h0; // @[ICache.scala 129:25]
  assign tag_bram_2_clock = clock;
  assign tag_bram_2_reset = reset;
  assign tag_bram_2_io_raddr = _GEN_1[11:6]; // @[ICache.scala 63:48]
  assign tag_bram_2_io_waddr = rset; // @[ICache.scala 138:23]
  assign tag_bram_2_io_wen = |tag_wstrb_1; // @[ICache.scala 137:39]
  assign tag_bram_2_io_wstrb = tag_wstrb_1; // @[ICache.scala 140:23]
  assign tag_bram_2_io_wdata = tag_wdata; // @[ICache.scala 139:23]
  assign bank_3_clock = clock;
  assign bank_3_reset = reset;
  assign bank_3_io_raddr = _GEN_1[11:3]; // @[ICache.scala 60:49]
  assign bank_3_io_waddr = {rset,axi_cnt_value[3:1]}; // @[Cat.scala 33:92]
  assign bank_3_io_wen = |data_wstrb_1_1; // @[ICache.scala 127:39]
  assign bank_3_io_wstrb = data_wstrb_1_1; // @[ICache.scala 130:19]
  assign bank_3_io_wdata = axi_cnt_value[0] ? io_axi_r_bits_data : 32'h0; // @[ICache.scala 129:25]
  assign tag_bram_3_clock = clock;
  assign tag_bram_3_reset = reset;
  assign tag_bram_3_io_raddr = _GEN_1[11:6]; // @[ICache.scala 63:48]
  assign tag_bram_3_io_waddr = rset; // @[ICache.scala 138:23]
  assign tag_bram_3_io_wen = |tag_wstrb_1; // @[ICache.scala 137:39]
  assign tag_bram_3_io_wstrb = tag_wstrb_1; // @[ICache.scala 140:23]
  assign tag_bram_3_io_wdata = tag_wdata; // @[ICache.scala 139:23]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 39:81]
      state <= 3'h0; // @[ICache.scala 39:81]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          state <= 3'h1; // @[ICache.scala 168:17]
        end else begin
          state <= _GEN_7207;
        end
      end
    end else if (3'h1 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_v_1 | ~inst_vpn[12] & io_cpu_tlb2_entry_v_0)) begin // @[ICache.scala 201:118]
        state <= 3'h0; // @[ICache.scala 202:22]
      end else begin
        state <= 3'h4; // @[ICache.scala 208:24]
      end
    end else if (3'h2 == state) begin // @[ICache.scala 164:17]
      state <= _GEN_11886;
    end else begin
      state <= _GEN_11947;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_0_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_0_0 <= _GEN_1027;
        end else begin
          valid_0_0 <= _GEN_7220;
        end
      end else begin
        valid_0_0 <= _GEN_1027;
      end
    end else begin
      valid_0_0 <= _GEN_1027;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_0_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_0_1 <= _GEN_1539;
        end else begin
          valid_0_1 <= _GEN_7221;
        end
      end else begin
        valid_0_1 <= _GEN_1539;
      end
    end else begin
      valid_0_1 <= _GEN_1539;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_1_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_1_0 <= _GEN_1028;
        end else begin
          valid_1_0 <= _GEN_7222;
        end
      end else begin
        valid_1_0 <= _GEN_1028;
      end
    end else begin
      valid_1_0 <= _GEN_1028;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_1_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_1_1 <= _GEN_1540;
        end else begin
          valid_1_1 <= _GEN_7223;
        end
      end else begin
        valid_1_1 <= _GEN_1540;
      end
    end else begin
      valid_1_1 <= _GEN_1540;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_2_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_2_0 <= _GEN_1029;
        end else begin
          valid_2_0 <= _GEN_7224;
        end
      end else begin
        valid_2_0 <= _GEN_1029;
      end
    end else begin
      valid_2_0 <= _GEN_1029;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_2_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_2_1 <= _GEN_1541;
        end else begin
          valid_2_1 <= _GEN_7225;
        end
      end else begin
        valid_2_1 <= _GEN_1541;
      end
    end else begin
      valid_2_1 <= _GEN_1541;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_3_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_3_0 <= _GEN_1030;
        end else begin
          valid_3_0 <= _GEN_7226;
        end
      end else begin
        valid_3_0 <= _GEN_1030;
      end
    end else begin
      valid_3_0 <= _GEN_1030;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_3_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_3_1 <= _GEN_1542;
        end else begin
          valid_3_1 <= _GEN_7227;
        end
      end else begin
        valid_3_1 <= _GEN_1542;
      end
    end else begin
      valid_3_1 <= _GEN_1542;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_4_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_4_0 <= _GEN_1031;
        end else begin
          valid_4_0 <= _GEN_7228;
        end
      end else begin
        valid_4_0 <= _GEN_1031;
      end
    end else begin
      valid_4_0 <= _GEN_1031;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_4_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_4_1 <= _GEN_1543;
        end else begin
          valid_4_1 <= _GEN_7229;
        end
      end else begin
        valid_4_1 <= _GEN_1543;
      end
    end else begin
      valid_4_1 <= _GEN_1543;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_5_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_5_0 <= _GEN_1032;
        end else begin
          valid_5_0 <= _GEN_7230;
        end
      end else begin
        valid_5_0 <= _GEN_1032;
      end
    end else begin
      valid_5_0 <= _GEN_1032;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_5_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_5_1 <= _GEN_1544;
        end else begin
          valid_5_1 <= _GEN_7231;
        end
      end else begin
        valid_5_1 <= _GEN_1544;
      end
    end else begin
      valid_5_1 <= _GEN_1544;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_6_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_6_0 <= _GEN_1033;
        end else begin
          valid_6_0 <= _GEN_7232;
        end
      end else begin
        valid_6_0 <= _GEN_1033;
      end
    end else begin
      valid_6_0 <= _GEN_1033;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_6_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_6_1 <= _GEN_1545;
        end else begin
          valid_6_1 <= _GEN_7233;
        end
      end else begin
        valid_6_1 <= _GEN_1545;
      end
    end else begin
      valid_6_1 <= _GEN_1545;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_7_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_7_0 <= _GEN_1034;
        end else begin
          valid_7_0 <= _GEN_7234;
        end
      end else begin
        valid_7_0 <= _GEN_1034;
      end
    end else begin
      valid_7_0 <= _GEN_1034;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_7_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_7_1 <= _GEN_1546;
        end else begin
          valid_7_1 <= _GEN_7235;
        end
      end else begin
        valid_7_1 <= _GEN_1546;
      end
    end else begin
      valid_7_1 <= _GEN_1546;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_8_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_8_0 <= _GEN_1035;
        end else begin
          valid_8_0 <= _GEN_7236;
        end
      end else begin
        valid_8_0 <= _GEN_1035;
      end
    end else begin
      valid_8_0 <= _GEN_1035;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_8_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_8_1 <= _GEN_1547;
        end else begin
          valid_8_1 <= _GEN_7237;
        end
      end else begin
        valid_8_1 <= _GEN_1547;
      end
    end else begin
      valid_8_1 <= _GEN_1547;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_9_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_9_0 <= _GEN_1036;
        end else begin
          valid_9_0 <= _GEN_7238;
        end
      end else begin
        valid_9_0 <= _GEN_1036;
      end
    end else begin
      valid_9_0 <= _GEN_1036;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_9_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_9_1 <= _GEN_1548;
        end else begin
          valid_9_1 <= _GEN_7239;
        end
      end else begin
        valid_9_1 <= _GEN_1548;
      end
    end else begin
      valid_9_1 <= _GEN_1548;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_10_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_10_0 <= _GEN_1037;
        end else begin
          valid_10_0 <= _GEN_7240;
        end
      end else begin
        valid_10_0 <= _GEN_1037;
      end
    end else begin
      valid_10_0 <= _GEN_1037;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_10_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_10_1 <= _GEN_1549;
        end else begin
          valid_10_1 <= _GEN_7241;
        end
      end else begin
        valid_10_1 <= _GEN_1549;
      end
    end else begin
      valid_10_1 <= _GEN_1549;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_11_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_11_0 <= _GEN_1038;
        end else begin
          valid_11_0 <= _GEN_7242;
        end
      end else begin
        valid_11_0 <= _GEN_1038;
      end
    end else begin
      valid_11_0 <= _GEN_1038;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_11_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_11_1 <= _GEN_1550;
        end else begin
          valid_11_1 <= _GEN_7243;
        end
      end else begin
        valid_11_1 <= _GEN_1550;
      end
    end else begin
      valid_11_1 <= _GEN_1550;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_12_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_12_0 <= _GEN_1039;
        end else begin
          valid_12_0 <= _GEN_7244;
        end
      end else begin
        valid_12_0 <= _GEN_1039;
      end
    end else begin
      valid_12_0 <= _GEN_1039;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_12_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_12_1 <= _GEN_1551;
        end else begin
          valid_12_1 <= _GEN_7245;
        end
      end else begin
        valid_12_1 <= _GEN_1551;
      end
    end else begin
      valid_12_1 <= _GEN_1551;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_13_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_13_0 <= _GEN_1040;
        end else begin
          valid_13_0 <= _GEN_7246;
        end
      end else begin
        valid_13_0 <= _GEN_1040;
      end
    end else begin
      valid_13_0 <= _GEN_1040;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_13_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_13_1 <= _GEN_1552;
        end else begin
          valid_13_1 <= _GEN_7247;
        end
      end else begin
        valid_13_1 <= _GEN_1552;
      end
    end else begin
      valid_13_1 <= _GEN_1552;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_14_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_14_0 <= _GEN_1041;
        end else begin
          valid_14_0 <= _GEN_7248;
        end
      end else begin
        valid_14_0 <= _GEN_1041;
      end
    end else begin
      valid_14_0 <= _GEN_1041;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_14_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_14_1 <= _GEN_1553;
        end else begin
          valid_14_1 <= _GEN_7249;
        end
      end else begin
        valid_14_1 <= _GEN_1553;
      end
    end else begin
      valid_14_1 <= _GEN_1553;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_15_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_15_0 <= _GEN_1042;
        end else begin
          valid_15_0 <= _GEN_7250;
        end
      end else begin
        valid_15_0 <= _GEN_1042;
      end
    end else begin
      valid_15_0 <= _GEN_1042;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_15_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_15_1 <= _GEN_1554;
        end else begin
          valid_15_1 <= _GEN_7251;
        end
      end else begin
        valid_15_1 <= _GEN_1554;
      end
    end else begin
      valid_15_1 <= _GEN_1554;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_16_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_16_0 <= _GEN_1043;
        end else begin
          valid_16_0 <= _GEN_7252;
        end
      end else begin
        valid_16_0 <= _GEN_1043;
      end
    end else begin
      valid_16_0 <= _GEN_1043;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_16_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_16_1 <= _GEN_1555;
        end else begin
          valid_16_1 <= _GEN_7253;
        end
      end else begin
        valid_16_1 <= _GEN_1555;
      end
    end else begin
      valid_16_1 <= _GEN_1555;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_17_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_17_0 <= _GEN_1044;
        end else begin
          valid_17_0 <= _GEN_7254;
        end
      end else begin
        valid_17_0 <= _GEN_1044;
      end
    end else begin
      valid_17_0 <= _GEN_1044;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_17_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_17_1 <= _GEN_1556;
        end else begin
          valid_17_1 <= _GEN_7255;
        end
      end else begin
        valid_17_1 <= _GEN_1556;
      end
    end else begin
      valid_17_1 <= _GEN_1556;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_18_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_18_0 <= _GEN_1045;
        end else begin
          valid_18_0 <= _GEN_7256;
        end
      end else begin
        valid_18_0 <= _GEN_1045;
      end
    end else begin
      valid_18_0 <= _GEN_1045;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_18_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_18_1 <= _GEN_1557;
        end else begin
          valid_18_1 <= _GEN_7257;
        end
      end else begin
        valid_18_1 <= _GEN_1557;
      end
    end else begin
      valid_18_1 <= _GEN_1557;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_19_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_19_0 <= _GEN_1046;
        end else begin
          valid_19_0 <= _GEN_7258;
        end
      end else begin
        valid_19_0 <= _GEN_1046;
      end
    end else begin
      valid_19_0 <= _GEN_1046;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_19_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_19_1 <= _GEN_1558;
        end else begin
          valid_19_1 <= _GEN_7259;
        end
      end else begin
        valid_19_1 <= _GEN_1558;
      end
    end else begin
      valid_19_1 <= _GEN_1558;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_20_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_20_0 <= _GEN_1047;
        end else begin
          valid_20_0 <= _GEN_7260;
        end
      end else begin
        valid_20_0 <= _GEN_1047;
      end
    end else begin
      valid_20_0 <= _GEN_1047;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_20_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_20_1 <= _GEN_1559;
        end else begin
          valid_20_1 <= _GEN_7261;
        end
      end else begin
        valid_20_1 <= _GEN_1559;
      end
    end else begin
      valid_20_1 <= _GEN_1559;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_21_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_21_0 <= _GEN_1048;
        end else begin
          valid_21_0 <= _GEN_7262;
        end
      end else begin
        valid_21_0 <= _GEN_1048;
      end
    end else begin
      valid_21_0 <= _GEN_1048;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_21_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_21_1 <= _GEN_1560;
        end else begin
          valid_21_1 <= _GEN_7263;
        end
      end else begin
        valid_21_1 <= _GEN_1560;
      end
    end else begin
      valid_21_1 <= _GEN_1560;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_22_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_22_0 <= _GEN_1049;
        end else begin
          valid_22_0 <= _GEN_7264;
        end
      end else begin
        valid_22_0 <= _GEN_1049;
      end
    end else begin
      valid_22_0 <= _GEN_1049;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_22_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_22_1 <= _GEN_1561;
        end else begin
          valid_22_1 <= _GEN_7265;
        end
      end else begin
        valid_22_1 <= _GEN_1561;
      end
    end else begin
      valid_22_1 <= _GEN_1561;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_23_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_23_0 <= _GEN_1050;
        end else begin
          valid_23_0 <= _GEN_7266;
        end
      end else begin
        valid_23_0 <= _GEN_1050;
      end
    end else begin
      valid_23_0 <= _GEN_1050;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_23_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_23_1 <= _GEN_1562;
        end else begin
          valid_23_1 <= _GEN_7267;
        end
      end else begin
        valid_23_1 <= _GEN_1562;
      end
    end else begin
      valid_23_1 <= _GEN_1562;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_24_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_24_0 <= _GEN_1051;
        end else begin
          valid_24_0 <= _GEN_7268;
        end
      end else begin
        valid_24_0 <= _GEN_1051;
      end
    end else begin
      valid_24_0 <= _GEN_1051;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_24_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_24_1 <= _GEN_1563;
        end else begin
          valid_24_1 <= _GEN_7269;
        end
      end else begin
        valid_24_1 <= _GEN_1563;
      end
    end else begin
      valid_24_1 <= _GEN_1563;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_25_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_25_0 <= _GEN_1052;
        end else begin
          valid_25_0 <= _GEN_7270;
        end
      end else begin
        valid_25_0 <= _GEN_1052;
      end
    end else begin
      valid_25_0 <= _GEN_1052;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_25_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_25_1 <= _GEN_1564;
        end else begin
          valid_25_1 <= _GEN_7271;
        end
      end else begin
        valid_25_1 <= _GEN_1564;
      end
    end else begin
      valid_25_1 <= _GEN_1564;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_26_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_26_0 <= _GEN_1053;
        end else begin
          valid_26_0 <= _GEN_7272;
        end
      end else begin
        valid_26_0 <= _GEN_1053;
      end
    end else begin
      valid_26_0 <= _GEN_1053;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_26_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_26_1 <= _GEN_1565;
        end else begin
          valid_26_1 <= _GEN_7273;
        end
      end else begin
        valid_26_1 <= _GEN_1565;
      end
    end else begin
      valid_26_1 <= _GEN_1565;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_27_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_27_0 <= _GEN_1054;
        end else begin
          valid_27_0 <= _GEN_7274;
        end
      end else begin
        valid_27_0 <= _GEN_1054;
      end
    end else begin
      valid_27_0 <= _GEN_1054;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_27_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_27_1 <= _GEN_1566;
        end else begin
          valid_27_1 <= _GEN_7275;
        end
      end else begin
        valid_27_1 <= _GEN_1566;
      end
    end else begin
      valid_27_1 <= _GEN_1566;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_28_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_28_0 <= _GEN_1055;
        end else begin
          valid_28_0 <= _GEN_7276;
        end
      end else begin
        valid_28_0 <= _GEN_1055;
      end
    end else begin
      valid_28_0 <= _GEN_1055;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_28_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_28_1 <= _GEN_1567;
        end else begin
          valid_28_1 <= _GEN_7277;
        end
      end else begin
        valid_28_1 <= _GEN_1567;
      end
    end else begin
      valid_28_1 <= _GEN_1567;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_29_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_29_0 <= _GEN_1056;
        end else begin
          valid_29_0 <= _GEN_7278;
        end
      end else begin
        valid_29_0 <= _GEN_1056;
      end
    end else begin
      valid_29_0 <= _GEN_1056;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_29_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_29_1 <= _GEN_1568;
        end else begin
          valid_29_1 <= _GEN_7279;
        end
      end else begin
        valid_29_1 <= _GEN_1568;
      end
    end else begin
      valid_29_1 <= _GEN_1568;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_30_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_30_0 <= _GEN_1057;
        end else begin
          valid_30_0 <= _GEN_7280;
        end
      end else begin
        valid_30_0 <= _GEN_1057;
      end
    end else begin
      valid_30_0 <= _GEN_1057;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_30_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_30_1 <= _GEN_1569;
        end else begin
          valid_30_1 <= _GEN_7281;
        end
      end else begin
        valid_30_1 <= _GEN_1569;
      end
    end else begin
      valid_30_1 <= _GEN_1569;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_31_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_31_0 <= _GEN_1058;
        end else begin
          valid_31_0 <= _GEN_7282;
        end
      end else begin
        valid_31_0 <= _GEN_1058;
      end
    end else begin
      valid_31_0 <= _GEN_1058;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_31_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_31_1 <= _GEN_1570;
        end else begin
          valid_31_1 <= _GEN_7283;
        end
      end else begin
        valid_31_1 <= _GEN_1570;
      end
    end else begin
      valid_31_1 <= _GEN_1570;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_32_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_32_0 <= _GEN_1059;
        end else begin
          valid_32_0 <= _GEN_7284;
        end
      end else begin
        valid_32_0 <= _GEN_1059;
      end
    end else begin
      valid_32_0 <= _GEN_1059;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_32_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_32_1 <= _GEN_1571;
        end else begin
          valid_32_1 <= _GEN_7285;
        end
      end else begin
        valid_32_1 <= _GEN_1571;
      end
    end else begin
      valid_32_1 <= _GEN_1571;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_33_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_33_0 <= _GEN_1060;
        end else begin
          valid_33_0 <= _GEN_7286;
        end
      end else begin
        valid_33_0 <= _GEN_1060;
      end
    end else begin
      valid_33_0 <= _GEN_1060;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_33_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_33_1 <= _GEN_1572;
        end else begin
          valid_33_1 <= _GEN_7287;
        end
      end else begin
        valid_33_1 <= _GEN_1572;
      end
    end else begin
      valid_33_1 <= _GEN_1572;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_34_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_34_0 <= _GEN_1061;
        end else begin
          valid_34_0 <= _GEN_7288;
        end
      end else begin
        valid_34_0 <= _GEN_1061;
      end
    end else begin
      valid_34_0 <= _GEN_1061;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_34_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_34_1 <= _GEN_1573;
        end else begin
          valid_34_1 <= _GEN_7289;
        end
      end else begin
        valid_34_1 <= _GEN_1573;
      end
    end else begin
      valid_34_1 <= _GEN_1573;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_35_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_35_0 <= _GEN_1062;
        end else begin
          valid_35_0 <= _GEN_7290;
        end
      end else begin
        valid_35_0 <= _GEN_1062;
      end
    end else begin
      valid_35_0 <= _GEN_1062;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_35_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_35_1 <= _GEN_1574;
        end else begin
          valid_35_1 <= _GEN_7291;
        end
      end else begin
        valid_35_1 <= _GEN_1574;
      end
    end else begin
      valid_35_1 <= _GEN_1574;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_36_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_36_0 <= _GEN_1063;
        end else begin
          valid_36_0 <= _GEN_7292;
        end
      end else begin
        valid_36_0 <= _GEN_1063;
      end
    end else begin
      valid_36_0 <= _GEN_1063;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_36_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_36_1 <= _GEN_1575;
        end else begin
          valid_36_1 <= _GEN_7293;
        end
      end else begin
        valid_36_1 <= _GEN_1575;
      end
    end else begin
      valid_36_1 <= _GEN_1575;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_37_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_37_0 <= _GEN_1064;
        end else begin
          valid_37_0 <= _GEN_7294;
        end
      end else begin
        valid_37_0 <= _GEN_1064;
      end
    end else begin
      valid_37_0 <= _GEN_1064;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_37_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_37_1 <= _GEN_1576;
        end else begin
          valid_37_1 <= _GEN_7295;
        end
      end else begin
        valid_37_1 <= _GEN_1576;
      end
    end else begin
      valid_37_1 <= _GEN_1576;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_38_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_38_0 <= _GEN_1065;
        end else begin
          valid_38_0 <= _GEN_7296;
        end
      end else begin
        valid_38_0 <= _GEN_1065;
      end
    end else begin
      valid_38_0 <= _GEN_1065;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_38_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_38_1 <= _GEN_1577;
        end else begin
          valid_38_1 <= _GEN_7297;
        end
      end else begin
        valid_38_1 <= _GEN_1577;
      end
    end else begin
      valid_38_1 <= _GEN_1577;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_39_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_39_0 <= _GEN_1066;
        end else begin
          valid_39_0 <= _GEN_7298;
        end
      end else begin
        valid_39_0 <= _GEN_1066;
      end
    end else begin
      valid_39_0 <= _GEN_1066;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_39_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_39_1 <= _GEN_1578;
        end else begin
          valid_39_1 <= _GEN_7299;
        end
      end else begin
        valid_39_1 <= _GEN_1578;
      end
    end else begin
      valid_39_1 <= _GEN_1578;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_40_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_40_0 <= _GEN_1067;
        end else begin
          valid_40_0 <= _GEN_7300;
        end
      end else begin
        valid_40_0 <= _GEN_1067;
      end
    end else begin
      valid_40_0 <= _GEN_1067;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_40_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_40_1 <= _GEN_1579;
        end else begin
          valid_40_1 <= _GEN_7301;
        end
      end else begin
        valid_40_1 <= _GEN_1579;
      end
    end else begin
      valid_40_1 <= _GEN_1579;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_41_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_41_0 <= _GEN_1068;
        end else begin
          valid_41_0 <= _GEN_7302;
        end
      end else begin
        valid_41_0 <= _GEN_1068;
      end
    end else begin
      valid_41_0 <= _GEN_1068;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_41_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_41_1 <= _GEN_1580;
        end else begin
          valid_41_1 <= _GEN_7303;
        end
      end else begin
        valid_41_1 <= _GEN_1580;
      end
    end else begin
      valid_41_1 <= _GEN_1580;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_42_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_42_0 <= _GEN_1069;
        end else begin
          valid_42_0 <= _GEN_7304;
        end
      end else begin
        valid_42_0 <= _GEN_1069;
      end
    end else begin
      valid_42_0 <= _GEN_1069;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_42_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_42_1 <= _GEN_1581;
        end else begin
          valid_42_1 <= _GEN_7305;
        end
      end else begin
        valid_42_1 <= _GEN_1581;
      end
    end else begin
      valid_42_1 <= _GEN_1581;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_43_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_43_0 <= _GEN_1070;
        end else begin
          valid_43_0 <= _GEN_7306;
        end
      end else begin
        valid_43_0 <= _GEN_1070;
      end
    end else begin
      valid_43_0 <= _GEN_1070;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_43_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_43_1 <= _GEN_1582;
        end else begin
          valid_43_1 <= _GEN_7307;
        end
      end else begin
        valid_43_1 <= _GEN_1582;
      end
    end else begin
      valid_43_1 <= _GEN_1582;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_44_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_44_0 <= _GEN_1071;
        end else begin
          valid_44_0 <= _GEN_7308;
        end
      end else begin
        valid_44_0 <= _GEN_1071;
      end
    end else begin
      valid_44_0 <= _GEN_1071;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_44_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_44_1 <= _GEN_1583;
        end else begin
          valid_44_1 <= _GEN_7309;
        end
      end else begin
        valid_44_1 <= _GEN_1583;
      end
    end else begin
      valid_44_1 <= _GEN_1583;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_45_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_45_0 <= _GEN_1072;
        end else begin
          valid_45_0 <= _GEN_7310;
        end
      end else begin
        valid_45_0 <= _GEN_1072;
      end
    end else begin
      valid_45_0 <= _GEN_1072;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_45_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_45_1 <= _GEN_1584;
        end else begin
          valid_45_1 <= _GEN_7311;
        end
      end else begin
        valid_45_1 <= _GEN_1584;
      end
    end else begin
      valid_45_1 <= _GEN_1584;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_46_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_46_0 <= _GEN_1073;
        end else begin
          valid_46_0 <= _GEN_7312;
        end
      end else begin
        valid_46_0 <= _GEN_1073;
      end
    end else begin
      valid_46_0 <= _GEN_1073;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_46_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_46_1 <= _GEN_1585;
        end else begin
          valid_46_1 <= _GEN_7313;
        end
      end else begin
        valid_46_1 <= _GEN_1585;
      end
    end else begin
      valid_46_1 <= _GEN_1585;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_47_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_47_0 <= _GEN_1074;
        end else begin
          valid_47_0 <= _GEN_7314;
        end
      end else begin
        valid_47_0 <= _GEN_1074;
      end
    end else begin
      valid_47_0 <= _GEN_1074;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_47_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_47_1 <= _GEN_1586;
        end else begin
          valid_47_1 <= _GEN_7315;
        end
      end else begin
        valid_47_1 <= _GEN_1586;
      end
    end else begin
      valid_47_1 <= _GEN_1586;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_48_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_48_0 <= _GEN_1075;
        end else begin
          valid_48_0 <= _GEN_7316;
        end
      end else begin
        valid_48_0 <= _GEN_1075;
      end
    end else begin
      valid_48_0 <= _GEN_1075;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_48_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_48_1 <= _GEN_1587;
        end else begin
          valid_48_1 <= _GEN_7317;
        end
      end else begin
        valid_48_1 <= _GEN_1587;
      end
    end else begin
      valid_48_1 <= _GEN_1587;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_49_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_49_0 <= _GEN_1076;
        end else begin
          valid_49_0 <= _GEN_7318;
        end
      end else begin
        valid_49_0 <= _GEN_1076;
      end
    end else begin
      valid_49_0 <= _GEN_1076;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_49_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_49_1 <= _GEN_1588;
        end else begin
          valid_49_1 <= _GEN_7319;
        end
      end else begin
        valid_49_1 <= _GEN_1588;
      end
    end else begin
      valid_49_1 <= _GEN_1588;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_50_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_50_0 <= _GEN_1077;
        end else begin
          valid_50_0 <= _GEN_7320;
        end
      end else begin
        valid_50_0 <= _GEN_1077;
      end
    end else begin
      valid_50_0 <= _GEN_1077;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_50_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_50_1 <= _GEN_1589;
        end else begin
          valid_50_1 <= _GEN_7321;
        end
      end else begin
        valid_50_1 <= _GEN_1589;
      end
    end else begin
      valid_50_1 <= _GEN_1589;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_51_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_51_0 <= _GEN_1078;
        end else begin
          valid_51_0 <= _GEN_7322;
        end
      end else begin
        valid_51_0 <= _GEN_1078;
      end
    end else begin
      valid_51_0 <= _GEN_1078;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_51_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_51_1 <= _GEN_1590;
        end else begin
          valid_51_1 <= _GEN_7323;
        end
      end else begin
        valid_51_1 <= _GEN_1590;
      end
    end else begin
      valid_51_1 <= _GEN_1590;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_52_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_52_0 <= _GEN_1079;
        end else begin
          valid_52_0 <= _GEN_7324;
        end
      end else begin
        valid_52_0 <= _GEN_1079;
      end
    end else begin
      valid_52_0 <= _GEN_1079;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_52_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_52_1 <= _GEN_1591;
        end else begin
          valid_52_1 <= _GEN_7325;
        end
      end else begin
        valid_52_1 <= _GEN_1591;
      end
    end else begin
      valid_52_1 <= _GEN_1591;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_53_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_53_0 <= _GEN_1080;
        end else begin
          valid_53_0 <= _GEN_7326;
        end
      end else begin
        valid_53_0 <= _GEN_1080;
      end
    end else begin
      valid_53_0 <= _GEN_1080;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_53_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_53_1 <= _GEN_1592;
        end else begin
          valid_53_1 <= _GEN_7327;
        end
      end else begin
        valid_53_1 <= _GEN_1592;
      end
    end else begin
      valid_53_1 <= _GEN_1592;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_54_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_54_0 <= _GEN_1081;
        end else begin
          valid_54_0 <= _GEN_7328;
        end
      end else begin
        valid_54_0 <= _GEN_1081;
      end
    end else begin
      valid_54_0 <= _GEN_1081;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_54_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_54_1 <= _GEN_1593;
        end else begin
          valid_54_1 <= _GEN_7329;
        end
      end else begin
        valid_54_1 <= _GEN_1593;
      end
    end else begin
      valid_54_1 <= _GEN_1593;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_55_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_55_0 <= _GEN_1082;
        end else begin
          valid_55_0 <= _GEN_7330;
        end
      end else begin
        valid_55_0 <= _GEN_1082;
      end
    end else begin
      valid_55_0 <= _GEN_1082;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_55_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_55_1 <= _GEN_1594;
        end else begin
          valid_55_1 <= _GEN_7331;
        end
      end else begin
        valid_55_1 <= _GEN_1594;
      end
    end else begin
      valid_55_1 <= _GEN_1594;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_56_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_56_0 <= _GEN_1083;
        end else begin
          valid_56_0 <= _GEN_7332;
        end
      end else begin
        valid_56_0 <= _GEN_1083;
      end
    end else begin
      valid_56_0 <= _GEN_1083;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_56_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_56_1 <= _GEN_1595;
        end else begin
          valid_56_1 <= _GEN_7333;
        end
      end else begin
        valid_56_1 <= _GEN_1595;
      end
    end else begin
      valid_56_1 <= _GEN_1595;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_57_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_57_0 <= _GEN_1084;
        end else begin
          valid_57_0 <= _GEN_7334;
        end
      end else begin
        valid_57_0 <= _GEN_1084;
      end
    end else begin
      valid_57_0 <= _GEN_1084;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_57_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_57_1 <= _GEN_1596;
        end else begin
          valid_57_1 <= _GEN_7335;
        end
      end else begin
        valid_57_1 <= _GEN_1596;
      end
    end else begin
      valid_57_1 <= _GEN_1596;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_58_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_58_0 <= _GEN_1085;
        end else begin
          valid_58_0 <= _GEN_7336;
        end
      end else begin
        valid_58_0 <= _GEN_1085;
      end
    end else begin
      valid_58_0 <= _GEN_1085;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_58_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_58_1 <= _GEN_1597;
        end else begin
          valid_58_1 <= _GEN_7337;
        end
      end else begin
        valid_58_1 <= _GEN_1597;
      end
    end else begin
      valid_58_1 <= _GEN_1597;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_59_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_59_0 <= _GEN_1086;
        end else begin
          valid_59_0 <= _GEN_7338;
        end
      end else begin
        valid_59_0 <= _GEN_1086;
      end
    end else begin
      valid_59_0 <= _GEN_1086;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_59_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_59_1 <= _GEN_1598;
        end else begin
          valid_59_1 <= _GEN_7339;
        end
      end else begin
        valid_59_1 <= _GEN_1598;
      end
    end else begin
      valid_59_1 <= _GEN_1598;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_60_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_60_0 <= _GEN_1087;
        end else begin
          valid_60_0 <= _GEN_7340;
        end
      end else begin
        valid_60_0 <= _GEN_1087;
      end
    end else begin
      valid_60_0 <= _GEN_1087;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_60_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_60_1 <= _GEN_1599;
        end else begin
          valid_60_1 <= _GEN_7341;
        end
      end else begin
        valid_60_1 <= _GEN_1599;
      end
    end else begin
      valid_60_1 <= _GEN_1599;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_61_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_61_0 <= _GEN_1088;
        end else begin
          valid_61_0 <= _GEN_7342;
        end
      end else begin
        valid_61_0 <= _GEN_1088;
      end
    end else begin
      valid_61_0 <= _GEN_1088;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_61_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_61_1 <= _GEN_1600;
        end else begin
          valid_61_1 <= _GEN_7343;
        end
      end else begin
        valid_61_1 <= _GEN_1600;
      end
    end else begin
      valid_61_1 <= _GEN_1600;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_62_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_62_0 <= _GEN_1089;
        end else begin
          valid_62_0 <= _GEN_7344;
        end
      end else begin
        valid_62_0 <= _GEN_1089;
      end
    end else begin
      valid_62_0 <= _GEN_1089;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_62_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_62_1 <= _GEN_1601;
        end else begin
          valid_62_1 <= _GEN_7345;
        end
      end else begin
        valid_62_1 <= _GEN_1601;
      end
    end else begin
      valid_62_1 <= _GEN_1601;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_63_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_63_0 <= _GEN_1090;
        end else begin
          valid_63_0 <= _GEN_7346;
        end
      end else begin
        valid_63_0 <= _GEN_1090;
      end
    end else begin
      valid_63_0 <= _GEN_1090;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_63_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_63_1 <= _GEN_1602;
        end else begin
          valid_63_1 <= _GEN_7347;
        end
      end else begin
        valid_63_1 <= _GEN_1602;
      end
    end else begin
      valid_63_1 <= _GEN_1602;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_64_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_64_0 <= _GEN_1091;
        end else begin
          valid_64_0 <= _GEN_7348;
        end
      end else begin
        valid_64_0 <= _GEN_1091;
      end
    end else begin
      valid_64_0 <= _GEN_1091;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_64_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_64_1 <= _GEN_1603;
        end else begin
          valid_64_1 <= _GEN_7349;
        end
      end else begin
        valid_64_1 <= _GEN_1603;
      end
    end else begin
      valid_64_1 <= _GEN_1603;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_65_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_65_0 <= _GEN_1092;
        end else begin
          valid_65_0 <= _GEN_7350;
        end
      end else begin
        valid_65_0 <= _GEN_1092;
      end
    end else begin
      valid_65_0 <= _GEN_1092;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_65_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_65_1 <= _GEN_1604;
        end else begin
          valid_65_1 <= _GEN_7351;
        end
      end else begin
        valid_65_1 <= _GEN_1604;
      end
    end else begin
      valid_65_1 <= _GEN_1604;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_66_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_66_0 <= _GEN_1093;
        end else begin
          valid_66_0 <= _GEN_7352;
        end
      end else begin
        valid_66_0 <= _GEN_1093;
      end
    end else begin
      valid_66_0 <= _GEN_1093;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_66_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_66_1 <= _GEN_1605;
        end else begin
          valid_66_1 <= _GEN_7353;
        end
      end else begin
        valid_66_1 <= _GEN_1605;
      end
    end else begin
      valid_66_1 <= _GEN_1605;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_67_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_67_0 <= _GEN_1094;
        end else begin
          valid_67_0 <= _GEN_7354;
        end
      end else begin
        valid_67_0 <= _GEN_1094;
      end
    end else begin
      valid_67_0 <= _GEN_1094;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_67_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_67_1 <= _GEN_1606;
        end else begin
          valid_67_1 <= _GEN_7355;
        end
      end else begin
        valid_67_1 <= _GEN_1606;
      end
    end else begin
      valid_67_1 <= _GEN_1606;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_68_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_68_0 <= _GEN_1095;
        end else begin
          valid_68_0 <= _GEN_7356;
        end
      end else begin
        valid_68_0 <= _GEN_1095;
      end
    end else begin
      valid_68_0 <= _GEN_1095;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_68_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_68_1 <= _GEN_1607;
        end else begin
          valid_68_1 <= _GEN_7357;
        end
      end else begin
        valid_68_1 <= _GEN_1607;
      end
    end else begin
      valid_68_1 <= _GEN_1607;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_69_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_69_0 <= _GEN_1096;
        end else begin
          valid_69_0 <= _GEN_7358;
        end
      end else begin
        valid_69_0 <= _GEN_1096;
      end
    end else begin
      valid_69_0 <= _GEN_1096;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_69_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_69_1 <= _GEN_1608;
        end else begin
          valid_69_1 <= _GEN_7359;
        end
      end else begin
        valid_69_1 <= _GEN_1608;
      end
    end else begin
      valid_69_1 <= _GEN_1608;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_70_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_70_0 <= _GEN_1097;
        end else begin
          valid_70_0 <= _GEN_7360;
        end
      end else begin
        valid_70_0 <= _GEN_1097;
      end
    end else begin
      valid_70_0 <= _GEN_1097;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_70_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_70_1 <= _GEN_1609;
        end else begin
          valid_70_1 <= _GEN_7361;
        end
      end else begin
        valid_70_1 <= _GEN_1609;
      end
    end else begin
      valid_70_1 <= _GEN_1609;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_71_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_71_0 <= _GEN_1098;
        end else begin
          valid_71_0 <= _GEN_7362;
        end
      end else begin
        valid_71_0 <= _GEN_1098;
      end
    end else begin
      valid_71_0 <= _GEN_1098;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_71_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_71_1 <= _GEN_1610;
        end else begin
          valid_71_1 <= _GEN_7363;
        end
      end else begin
        valid_71_1 <= _GEN_1610;
      end
    end else begin
      valid_71_1 <= _GEN_1610;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_72_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_72_0 <= _GEN_1099;
        end else begin
          valid_72_0 <= _GEN_7364;
        end
      end else begin
        valid_72_0 <= _GEN_1099;
      end
    end else begin
      valid_72_0 <= _GEN_1099;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_72_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_72_1 <= _GEN_1611;
        end else begin
          valid_72_1 <= _GEN_7365;
        end
      end else begin
        valid_72_1 <= _GEN_1611;
      end
    end else begin
      valid_72_1 <= _GEN_1611;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_73_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_73_0 <= _GEN_1100;
        end else begin
          valid_73_0 <= _GEN_7366;
        end
      end else begin
        valid_73_0 <= _GEN_1100;
      end
    end else begin
      valid_73_0 <= _GEN_1100;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_73_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_73_1 <= _GEN_1612;
        end else begin
          valid_73_1 <= _GEN_7367;
        end
      end else begin
        valid_73_1 <= _GEN_1612;
      end
    end else begin
      valid_73_1 <= _GEN_1612;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_74_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_74_0 <= _GEN_1101;
        end else begin
          valid_74_0 <= _GEN_7368;
        end
      end else begin
        valid_74_0 <= _GEN_1101;
      end
    end else begin
      valid_74_0 <= _GEN_1101;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_74_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_74_1 <= _GEN_1613;
        end else begin
          valid_74_1 <= _GEN_7369;
        end
      end else begin
        valid_74_1 <= _GEN_1613;
      end
    end else begin
      valid_74_1 <= _GEN_1613;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_75_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_75_0 <= _GEN_1102;
        end else begin
          valid_75_0 <= _GEN_7370;
        end
      end else begin
        valid_75_0 <= _GEN_1102;
      end
    end else begin
      valid_75_0 <= _GEN_1102;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_75_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_75_1 <= _GEN_1614;
        end else begin
          valid_75_1 <= _GEN_7371;
        end
      end else begin
        valid_75_1 <= _GEN_1614;
      end
    end else begin
      valid_75_1 <= _GEN_1614;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_76_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_76_0 <= _GEN_1103;
        end else begin
          valid_76_0 <= _GEN_7372;
        end
      end else begin
        valid_76_0 <= _GEN_1103;
      end
    end else begin
      valid_76_0 <= _GEN_1103;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_76_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_76_1 <= _GEN_1615;
        end else begin
          valid_76_1 <= _GEN_7373;
        end
      end else begin
        valid_76_1 <= _GEN_1615;
      end
    end else begin
      valid_76_1 <= _GEN_1615;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_77_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_77_0 <= _GEN_1104;
        end else begin
          valid_77_0 <= _GEN_7374;
        end
      end else begin
        valid_77_0 <= _GEN_1104;
      end
    end else begin
      valid_77_0 <= _GEN_1104;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_77_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_77_1 <= _GEN_1616;
        end else begin
          valid_77_1 <= _GEN_7375;
        end
      end else begin
        valid_77_1 <= _GEN_1616;
      end
    end else begin
      valid_77_1 <= _GEN_1616;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_78_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_78_0 <= _GEN_1105;
        end else begin
          valid_78_0 <= _GEN_7376;
        end
      end else begin
        valid_78_0 <= _GEN_1105;
      end
    end else begin
      valid_78_0 <= _GEN_1105;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_78_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_78_1 <= _GEN_1617;
        end else begin
          valid_78_1 <= _GEN_7377;
        end
      end else begin
        valid_78_1 <= _GEN_1617;
      end
    end else begin
      valid_78_1 <= _GEN_1617;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_79_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_79_0 <= _GEN_1106;
        end else begin
          valid_79_0 <= _GEN_7378;
        end
      end else begin
        valid_79_0 <= _GEN_1106;
      end
    end else begin
      valid_79_0 <= _GEN_1106;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_79_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_79_1 <= _GEN_1618;
        end else begin
          valid_79_1 <= _GEN_7379;
        end
      end else begin
        valid_79_1 <= _GEN_1618;
      end
    end else begin
      valid_79_1 <= _GEN_1618;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_80_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_80_0 <= _GEN_1107;
        end else begin
          valid_80_0 <= _GEN_7380;
        end
      end else begin
        valid_80_0 <= _GEN_1107;
      end
    end else begin
      valid_80_0 <= _GEN_1107;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_80_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_80_1 <= _GEN_1619;
        end else begin
          valid_80_1 <= _GEN_7381;
        end
      end else begin
        valid_80_1 <= _GEN_1619;
      end
    end else begin
      valid_80_1 <= _GEN_1619;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_81_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_81_0 <= _GEN_1108;
        end else begin
          valid_81_0 <= _GEN_7382;
        end
      end else begin
        valid_81_0 <= _GEN_1108;
      end
    end else begin
      valid_81_0 <= _GEN_1108;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_81_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_81_1 <= _GEN_1620;
        end else begin
          valid_81_1 <= _GEN_7383;
        end
      end else begin
        valid_81_1 <= _GEN_1620;
      end
    end else begin
      valid_81_1 <= _GEN_1620;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_82_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_82_0 <= _GEN_1109;
        end else begin
          valid_82_0 <= _GEN_7384;
        end
      end else begin
        valid_82_0 <= _GEN_1109;
      end
    end else begin
      valid_82_0 <= _GEN_1109;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_82_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_82_1 <= _GEN_1621;
        end else begin
          valid_82_1 <= _GEN_7385;
        end
      end else begin
        valid_82_1 <= _GEN_1621;
      end
    end else begin
      valid_82_1 <= _GEN_1621;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_83_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_83_0 <= _GEN_1110;
        end else begin
          valid_83_0 <= _GEN_7386;
        end
      end else begin
        valid_83_0 <= _GEN_1110;
      end
    end else begin
      valid_83_0 <= _GEN_1110;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_83_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_83_1 <= _GEN_1622;
        end else begin
          valid_83_1 <= _GEN_7387;
        end
      end else begin
        valid_83_1 <= _GEN_1622;
      end
    end else begin
      valid_83_1 <= _GEN_1622;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_84_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_84_0 <= _GEN_1111;
        end else begin
          valid_84_0 <= _GEN_7388;
        end
      end else begin
        valid_84_0 <= _GEN_1111;
      end
    end else begin
      valid_84_0 <= _GEN_1111;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_84_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_84_1 <= _GEN_1623;
        end else begin
          valid_84_1 <= _GEN_7389;
        end
      end else begin
        valid_84_1 <= _GEN_1623;
      end
    end else begin
      valid_84_1 <= _GEN_1623;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_85_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_85_0 <= _GEN_1112;
        end else begin
          valid_85_0 <= _GEN_7390;
        end
      end else begin
        valid_85_0 <= _GEN_1112;
      end
    end else begin
      valid_85_0 <= _GEN_1112;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_85_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_85_1 <= _GEN_1624;
        end else begin
          valid_85_1 <= _GEN_7391;
        end
      end else begin
        valid_85_1 <= _GEN_1624;
      end
    end else begin
      valid_85_1 <= _GEN_1624;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_86_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_86_0 <= _GEN_1113;
        end else begin
          valid_86_0 <= _GEN_7392;
        end
      end else begin
        valid_86_0 <= _GEN_1113;
      end
    end else begin
      valid_86_0 <= _GEN_1113;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_86_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_86_1 <= _GEN_1625;
        end else begin
          valid_86_1 <= _GEN_7393;
        end
      end else begin
        valid_86_1 <= _GEN_1625;
      end
    end else begin
      valid_86_1 <= _GEN_1625;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_87_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_87_0 <= _GEN_1114;
        end else begin
          valid_87_0 <= _GEN_7394;
        end
      end else begin
        valid_87_0 <= _GEN_1114;
      end
    end else begin
      valid_87_0 <= _GEN_1114;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_87_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_87_1 <= _GEN_1626;
        end else begin
          valid_87_1 <= _GEN_7395;
        end
      end else begin
        valid_87_1 <= _GEN_1626;
      end
    end else begin
      valid_87_1 <= _GEN_1626;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_88_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_88_0 <= _GEN_1115;
        end else begin
          valid_88_0 <= _GEN_7396;
        end
      end else begin
        valid_88_0 <= _GEN_1115;
      end
    end else begin
      valid_88_0 <= _GEN_1115;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_88_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_88_1 <= _GEN_1627;
        end else begin
          valid_88_1 <= _GEN_7397;
        end
      end else begin
        valid_88_1 <= _GEN_1627;
      end
    end else begin
      valid_88_1 <= _GEN_1627;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_89_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_89_0 <= _GEN_1116;
        end else begin
          valid_89_0 <= _GEN_7398;
        end
      end else begin
        valid_89_0 <= _GEN_1116;
      end
    end else begin
      valid_89_0 <= _GEN_1116;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_89_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_89_1 <= _GEN_1628;
        end else begin
          valid_89_1 <= _GEN_7399;
        end
      end else begin
        valid_89_1 <= _GEN_1628;
      end
    end else begin
      valid_89_1 <= _GEN_1628;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_90_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_90_0 <= _GEN_1117;
        end else begin
          valid_90_0 <= _GEN_7400;
        end
      end else begin
        valid_90_0 <= _GEN_1117;
      end
    end else begin
      valid_90_0 <= _GEN_1117;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_90_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_90_1 <= _GEN_1629;
        end else begin
          valid_90_1 <= _GEN_7401;
        end
      end else begin
        valid_90_1 <= _GEN_1629;
      end
    end else begin
      valid_90_1 <= _GEN_1629;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_91_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_91_0 <= _GEN_1118;
        end else begin
          valid_91_0 <= _GEN_7402;
        end
      end else begin
        valid_91_0 <= _GEN_1118;
      end
    end else begin
      valid_91_0 <= _GEN_1118;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_91_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_91_1 <= _GEN_1630;
        end else begin
          valid_91_1 <= _GEN_7403;
        end
      end else begin
        valid_91_1 <= _GEN_1630;
      end
    end else begin
      valid_91_1 <= _GEN_1630;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_92_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_92_0 <= _GEN_1119;
        end else begin
          valid_92_0 <= _GEN_7404;
        end
      end else begin
        valid_92_0 <= _GEN_1119;
      end
    end else begin
      valid_92_0 <= _GEN_1119;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_92_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_92_1 <= _GEN_1631;
        end else begin
          valid_92_1 <= _GEN_7405;
        end
      end else begin
        valid_92_1 <= _GEN_1631;
      end
    end else begin
      valid_92_1 <= _GEN_1631;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_93_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_93_0 <= _GEN_1120;
        end else begin
          valid_93_0 <= _GEN_7406;
        end
      end else begin
        valid_93_0 <= _GEN_1120;
      end
    end else begin
      valid_93_0 <= _GEN_1120;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_93_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_93_1 <= _GEN_1632;
        end else begin
          valid_93_1 <= _GEN_7407;
        end
      end else begin
        valid_93_1 <= _GEN_1632;
      end
    end else begin
      valid_93_1 <= _GEN_1632;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_94_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_94_0 <= _GEN_1121;
        end else begin
          valid_94_0 <= _GEN_7408;
        end
      end else begin
        valid_94_0 <= _GEN_1121;
      end
    end else begin
      valid_94_0 <= _GEN_1121;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_94_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_94_1 <= _GEN_1633;
        end else begin
          valid_94_1 <= _GEN_7409;
        end
      end else begin
        valid_94_1 <= _GEN_1633;
      end
    end else begin
      valid_94_1 <= _GEN_1633;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_95_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_95_0 <= _GEN_1122;
        end else begin
          valid_95_0 <= _GEN_7410;
        end
      end else begin
        valid_95_0 <= _GEN_1122;
      end
    end else begin
      valid_95_0 <= _GEN_1122;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_95_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_95_1 <= _GEN_1634;
        end else begin
          valid_95_1 <= _GEN_7411;
        end
      end else begin
        valid_95_1 <= _GEN_1634;
      end
    end else begin
      valid_95_1 <= _GEN_1634;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_96_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_96_0 <= _GEN_1123;
        end else begin
          valid_96_0 <= _GEN_7412;
        end
      end else begin
        valid_96_0 <= _GEN_1123;
      end
    end else begin
      valid_96_0 <= _GEN_1123;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_96_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_96_1 <= _GEN_1635;
        end else begin
          valid_96_1 <= _GEN_7413;
        end
      end else begin
        valid_96_1 <= _GEN_1635;
      end
    end else begin
      valid_96_1 <= _GEN_1635;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_97_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_97_0 <= _GEN_1124;
        end else begin
          valid_97_0 <= _GEN_7414;
        end
      end else begin
        valid_97_0 <= _GEN_1124;
      end
    end else begin
      valid_97_0 <= _GEN_1124;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_97_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_97_1 <= _GEN_1636;
        end else begin
          valid_97_1 <= _GEN_7415;
        end
      end else begin
        valid_97_1 <= _GEN_1636;
      end
    end else begin
      valid_97_1 <= _GEN_1636;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_98_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_98_0 <= _GEN_1125;
        end else begin
          valid_98_0 <= _GEN_7416;
        end
      end else begin
        valid_98_0 <= _GEN_1125;
      end
    end else begin
      valid_98_0 <= _GEN_1125;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_98_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_98_1 <= _GEN_1637;
        end else begin
          valid_98_1 <= _GEN_7417;
        end
      end else begin
        valid_98_1 <= _GEN_1637;
      end
    end else begin
      valid_98_1 <= _GEN_1637;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_99_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_99_0 <= _GEN_1126;
        end else begin
          valid_99_0 <= _GEN_7418;
        end
      end else begin
        valid_99_0 <= _GEN_1126;
      end
    end else begin
      valid_99_0 <= _GEN_1126;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_99_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_99_1 <= _GEN_1638;
        end else begin
          valid_99_1 <= _GEN_7419;
        end
      end else begin
        valid_99_1 <= _GEN_1638;
      end
    end else begin
      valid_99_1 <= _GEN_1638;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_100_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_100_0 <= _GEN_1127;
        end else begin
          valid_100_0 <= _GEN_7420;
        end
      end else begin
        valid_100_0 <= _GEN_1127;
      end
    end else begin
      valid_100_0 <= _GEN_1127;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_100_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_100_1 <= _GEN_1639;
        end else begin
          valid_100_1 <= _GEN_7421;
        end
      end else begin
        valid_100_1 <= _GEN_1639;
      end
    end else begin
      valid_100_1 <= _GEN_1639;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_101_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_101_0 <= _GEN_1128;
        end else begin
          valid_101_0 <= _GEN_7422;
        end
      end else begin
        valid_101_0 <= _GEN_1128;
      end
    end else begin
      valid_101_0 <= _GEN_1128;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_101_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_101_1 <= _GEN_1640;
        end else begin
          valid_101_1 <= _GEN_7423;
        end
      end else begin
        valid_101_1 <= _GEN_1640;
      end
    end else begin
      valid_101_1 <= _GEN_1640;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_102_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_102_0 <= _GEN_1129;
        end else begin
          valid_102_0 <= _GEN_7424;
        end
      end else begin
        valid_102_0 <= _GEN_1129;
      end
    end else begin
      valid_102_0 <= _GEN_1129;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_102_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_102_1 <= _GEN_1641;
        end else begin
          valid_102_1 <= _GEN_7425;
        end
      end else begin
        valid_102_1 <= _GEN_1641;
      end
    end else begin
      valid_102_1 <= _GEN_1641;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_103_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_103_0 <= _GEN_1130;
        end else begin
          valid_103_0 <= _GEN_7426;
        end
      end else begin
        valid_103_0 <= _GEN_1130;
      end
    end else begin
      valid_103_0 <= _GEN_1130;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_103_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_103_1 <= _GEN_1642;
        end else begin
          valid_103_1 <= _GEN_7427;
        end
      end else begin
        valid_103_1 <= _GEN_1642;
      end
    end else begin
      valid_103_1 <= _GEN_1642;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_104_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_104_0 <= _GEN_1131;
        end else begin
          valid_104_0 <= _GEN_7428;
        end
      end else begin
        valid_104_0 <= _GEN_1131;
      end
    end else begin
      valid_104_0 <= _GEN_1131;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_104_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_104_1 <= _GEN_1643;
        end else begin
          valid_104_1 <= _GEN_7429;
        end
      end else begin
        valid_104_1 <= _GEN_1643;
      end
    end else begin
      valid_104_1 <= _GEN_1643;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_105_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_105_0 <= _GEN_1132;
        end else begin
          valid_105_0 <= _GEN_7430;
        end
      end else begin
        valid_105_0 <= _GEN_1132;
      end
    end else begin
      valid_105_0 <= _GEN_1132;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_105_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_105_1 <= _GEN_1644;
        end else begin
          valid_105_1 <= _GEN_7431;
        end
      end else begin
        valid_105_1 <= _GEN_1644;
      end
    end else begin
      valid_105_1 <= _GEN_1644;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_106_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_106_0 <= _GEN_1133;
        end else begin
          valid_106_0 <= _GEN_7432;
        end
      end else begin
        valid_106_0 <= _GEN_1133;
      end
    end else begin
      valid_106_0 <= _GEN_1133;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_106_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_106_1 <= _GEN_1645;
        end else begin
          valid_106_1 <= _GEN_7433;
        end
      end else begin
        valid_106_1 <= _GEN_1645;
      end
    end else begin
      valid_106_1 <= _GEN_1645;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_107_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_107_0 <= _GEN_1134;
        end else begin
          valid_107_0 <= _GEN_7434;
        end
      end else begin
        valid_107_0 <= _GEN_1134;
      end
    end else begin
      valid_107_0 <= _GEN_1134;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_107_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_107_1 <= _GEN_1646;
        end else begin
          valid_107_1 <= _GEN_7435;
        end
      end else begin
        valid_107_1 <= _GEN_1646;
      end
    end else begin
      valid_107_1 <= _GEN_1646;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_108_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_108_0 <= _GEN_1135;
        end else begin
          valid_108_0 <= _GEN_7436;
        end
      end else begin
        valid_108_0 <= _GEN_1135;
      end
    end else begin
      valid_108_0 <= _GEN_1135;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_108_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_108_1 <= _GEN_1647;
        end else begin
          valid_108_1 <= _GEN_7437;
        end
      end else begin
        valid_108_1 <= _GEN_1647;
      end
    end else begin
      valid_108_1 <= _GEN_1647;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_109_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_109_0 <= _GEN_1136;
        end else begin
          valid_109_0 <= _GEN_7438;
        end
      end else begin
        valid_109_0 <= _GEN_1136;
      end
    end else begin
      valid_109_0 <= _GEN_1136;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_109_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_109_1 <= _GEN_1648;
        end else begin
          valid_109_1 <= _GEN_7439;
        end
      end else begin
        valid_109_1 <= _GEN_1648;
      end
    end else begin
      valid_109_1 <= _GEN_1648;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_110_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_110_0 <= _GEN_1137;
        end else begin
          valid_110_0 <= _GEN_7440;
        end
      end else begin
        valid_110_0 <= _GEN_1137;
      end
    end else begin
      valid_110_0 <= _GEN_1137;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_110_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_110_1 <= _GEN_1649;
        end else begin
          valid_110_1 <= _GEN_7441;
        end
      end else begin
        valid_110_1 <= _GEN_1649;
      end
    end else begin
      valid_110_1 <= _GEN_1649;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_111_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_111_0 <= _GEN_1138;
        end else begin
          valid_111_0 <= _GEN_7442;
        end
      end else begin
        valid_111_0 <= _GEN_1138;
      end
    end else begin
      valid_111_0 <= _GEN_1138;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_111_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_111_1 <= _GEN_1650;
        end else begin
          valid_111_1 <= _GEN_7443;
        end
      end else begin
        valid_111_1 <= _GEN_1650;
      end
    end else begin
      valid_111_1 <= _GEN_1650;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_112_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_112_0 <= _GEN_1139;
        end else begin
          valid_112_0 <= _GEN_7444;
        end
      end else begin
        valid_112_0 <= _GEN_1139;
      end
    end else begin
      valid_112_0 <= _GEN_1139;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_112_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_112_1 <= _GEN_1651;
        end else begin
          valid_112_1 <= _GEN_7445;
        end
      end else begin
        valid_112_1 <= _GEN_1651;
      end
    end else begin
      valid_112_1 <= _GEN_1651;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_113_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_113_0 <= _GEN_1140;
        end else begin
          valid_113_0 <= _GEN_7446;
        end
      end else begin
        valid_113_0 <= _GEN_1140;
      end
    end else begin
      valid_113_0 <= _GEN_1140;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_113_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_113_1 <= _GEN_1652;
        end else begin
          valid_113_1 <= _GEN_7447;
        end
      end else begin
        valid_113_1 <= _GEN_1652;
      end
    end else begin
      valid_113_1 <= _GEN_1652;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_114_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_114_0 <= _GEN_1141;
        end else begin
          valid_114_0 <= _GEN_7448;
        end
      end else begin
        valid_114_0 <= _GEN_1141;
      end
    end else begin
      valid_114_0 <= _GEN_1141;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_114_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_114_1 <= _GEN_1653;
        end else begin
          valid_114_1 <= _GEN_7449;
        end
      end else begin
        valid_114_1 <= _GEN_1653;
      end
    end else begin
      valid_114_1 <= _GEN_1653;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_115_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_115_0 <= _GEN_1142;
        end else begin
          valid_115_0 <= _GEN_7450;
        end
      end else begin
        valid_115_0 <= _GEN_1142;
      end
    end else begin
      valid_115_0 <= _GEN_1142;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_115_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_115_1 <= _GEN_1654;
        end else begin
          valid_115_1 <= _GEN_7451;
        end
      end else begin
        valid_115_1 <= _GEN_1654;
      end
    end else begin
      valid_115_1 <= _GEN_1654;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_116_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_116_0 <= _GEN_1143;
        end else begin
          valid_116_0 <= _GEN_7452;
        end
      end else begin
        valid_116_0 <= _GEN_1143;
      end
    end else begin
      valid_116_0 <= _GEN_1143;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_116_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_116_1 <= _GEN_1655;
        end else begin
          valid_116_1 <= _GEN_7453;
        end
      end else begin
        valid_116_1 <= _GEN_1655;
      end
    end else begin
      valid_116_1 <= _GEN_1655;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_117_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_117_0 <= _GEN_1144;
        end else begin
          valid_117_0 <= _GEN_7454;
        end
      end else begin
        valid_117_0 <= _GEN_1144;
      end
    end else begin
      valid_117_0 <= _GEN_1144;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_117_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_117_1 <= _GEN_1656;
        end else begin
          valid_117_1 <= _GEN_7455;
        end
      end else begin
        valid_117_1 <= _GEN_1656;
      end
    end else begin
      valid_117_1 <= _GEN_1656;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_118_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_118_0 <= _GEN_1145;
        end else begin
          valid_118_0 <= _GEN_7456;
        end
      end else begin
        valid_118_0 <= _GEN_1145;
      end
    end else begin
      valid_118_0 <= _GEN_1145;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_118_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_118_1 <= _GEN_1657;
        end else begin
          valid_118_1 <= _GEN_7457;
        end
      end else begin
        valid_118_1 <= _GEN_1657;
      end
    end else begin
      valid_118_1 <= _GEN_1657;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_119_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_119_0 <= _GEN_1146;
        end else begin
          valid_119_0 <= _GEN_7458;
        end
      end else begin
        valid_119_0 <= _GEN_1146;
      end
    end else begin
      valid_119_0 <= _GEN_1146;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_119_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_119_1 <= _GEN_1658;
        end else begin
          valid_119_1 <= _GEN_7459;
        end
      end else begin
        valid_119_1 <= _GEN_1658;
      end
    end else begin
      valid_119_1 <= _GEN_1658;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_120_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_120_0 <= _GEN_1147;
        end else begin
          valid_120_0 <= _GEN_7460;
        end
      end else begin
        valid_120_0 <= _GEN_1147;
      end
    end else begin
      valid_120_0 <= _GEN_1147;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_120_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_120_1 <= _GEN_1659;
        end else begin
          valid_120_1 <= _GEN_7461;
        end
      end else begin
        valid_120_1 <= _GEN_1659;
      end
    end else begin
      valid_120_1 <= _GEN_1659;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_121_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_121_0 <= _GEN_1148;
        end else begin
          valid_121_0 <= _GEN_7462;
        end
      end else begin
        valid_121_0 <= _GEN_1148;
      end
    end else begin
      valid_121_0 <= _GEN_1148;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_121_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_121_1 <= _GEN_1660;
        end else begin
          valid_121_1 <= _GEN_7463;
        end
      end else begin
        valid_121_1 <= _GEN_1660;
      end
    end else begin
      valid_121_1 <= _GEN_1660;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_122_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_122_0 <= _GEN_1149;
        end else begin
          valid_122_0 <= _GEN_7464;
        end
      end else begin
        valid_122_0 <= _GEN_1149;
      end
    end else begin
      valid_122_0 <= _GEN_1149;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_122_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_122_1 <= _GEN_1661;
        end else begin
          valid_122_1 <= _GEN_7465;
        end
      end else begin
        valid_122_1 <= _GEN_1661;
      end
    end else begin
      valid_122_1 <= _GEN_1661;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_123_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_123_0 <= _GEN_1150;
        end else begin
          valid_123_0 <= _GEN_7466;
        end
      end else begin
        valid_123_0 <= _GEN_1150;
      end
    end else begin
      valid_123_0 <= _GEN_1150;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_123_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_123_1 <= _GEN_1662;
        end else begin
          valid_123_1 <= _GEN_7467;
        end
      end else begin
        valid_123_1 <= _GEN_1662;
      end
    end else begin
      valid_123_1 <= _GEN_1662;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_124_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_124_0 <= _GEN_1151;
        end else begin
          valid_124_0 <= _GEN_7468;
        end
      end else begin
        valid_124_0 <= _GEN_1151;
      end
    end else begin
      valid_124_0 <= _GEN_1151;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_124_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_124_1 <= _GEN_1663;
        end else begin
          valid_124_1 <= _GEN_7469;
        end
      end else begin
        valid_124_1 <= _GEN_1663;
      end
    end else begin
      valid_124_1 <= _GEN_1663;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_125_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_125_0 <= _GEN_1152;
        end else begin
          valid_125_0 <= _GEN_7470;
        end
      end else begin
        valid_125_0 <= _GEN_1152;
      end
    end else begin
      valid_125_0 <= _GEN_1152;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_125_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_125_1 <= _GEN_1664;
        end else begin
          valid_125_1 <= _GEN_7471;
        end
      end else begin
        valid_125_1 <= _GEN_1664;
      end
    end else begin
      valid_125_1 <= _GEN_1664;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_126_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_126_0 <= _GEN_1153;
        end else begin
          valid_126_0 <= _GEN_7472;
        end
      end else begin
        valid_126_0 <= _GEN_1153;
      end
    end else begin
      valid_126_0 <= _GEN_1153;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_126_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_126_1 <= _GEN_1665;
        end else begin
          valid_126_1 <= _GEN_7473;
        end
      end else begin
        valid_126_1 <= _GEN_1665;
      end
    end else begin
      valid_126_1 <= _GEN_1665;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_127_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_127_0 <= _GEN_1154;
        end else begin
          valid_127_0 <= _GEN_7474;
        end
      end else begin
        valid_127_0 <= _GEN_1154;
      end
    end else begin
      valid_127_0 <= _GEN_1154;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_127_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_127_1 <= _GEN_1666;
        end else begin
          valid_127_1 <= _GEN_7475;
        end
      end else begin
        valid_127_1 <= _GEN_1666;
      end
    end else begin
      valid_127_1 <= _GEN_1666;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_128_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_128_0 <= _GEN_1155;
        end else begin
          valid_128_0 <= _GEN_7476;
        end
      end else begin
        valid_128_0 <= _GEN_1155;
      end
    end else begin
      valid_128_0 <= _GEN_1155;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_128_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_128_1 <= _GEN_1667;
        end else begin
          valid_128_1 <= _GEN_7477;
        end
      end else begin
        valid_128_1 <= _GEN_1667;
      end
    end else begin
      valid_128_1 <= _GEN_1667;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_129_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_129_0 <= _GEN_1156;
        end else begin
          valid_129_0 <= _GEN_7478;
        end
      end else begin
        valid_129_0 <= _GEN_1156;
      end
    end else begin
      valid_129_0 <= _GEN_1156;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_129_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_129_1 <= _GEN_1668;
        end else begin
          valid_129_1 <= _GEN_7479;
        end
      end else begin
        valid_129_1 <= _GEN_1668;
      end
    end else begin
      valid_129_1 <= _GEN_1668;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_130_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_130_0 <= _GEN_1157;
        end else begin
          valid_130_0 <= _GEN_7480;
        end
      end else begin
        valid_130_0 <= _GEN_1157;
      end
    end else begin
      valid_130_0 <= _GEN_1157;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_130_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_130_1 <= _GEN_1669;
        end else begin
          valid_130_1 <= _GEN_7481;
        end
      end else begin
        valid_130_1 <= _GEN_1669;
      end
    end else begin
      valid_130_1 <= _GEN_1669;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_131_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_131_0 <= _GEN_1158;
        end else begin
          valid_131_0 <= _GEN_7482;
        end
      end else begin
        valid_131_0 <= _GEN_1158;
      end
    end else begin
      valid_131_0 <= _GEN_1158;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_131_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_131_1 <= _GEN_1670;
        end else begin
          valid_131_1 <= _GEN_7483;
        end
      end else begin
        valid_131_1 <= _GEN_1670;
      end
    end else begin
      valid_131_1 <= _GEN_1670;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_132_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_132_0 <= _GEN_1159;
        end else begin
          valid_132_0 <= _GEN_7484;
        end
      end else begin
        valid_132_0 <= _GEN_1159;
      end
    end else begin
      valid_132_0 <= _GEN_1159;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_132_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_132_1 <= _GEN_1671;
        end else begin
          valid_132_1 <= _GEN_7485;
        end
      end else begin
        valid_132_1 <= _GEN_1671;
      end
    end else begin
      valid_132_1 <= _GEN_1671;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_133_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_133_0 <= _GEN_1160;
        end else begin
          valid_133_0 <= _GEN_7486;
        end
      end else begin
        valid_133_0 <= _GEN_1160;
      end
    end else begin
      valid_133_0 <= _GEN_1160;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_133_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_133_1 <= _GEN_1672;
        end else begin
          valid_133_1 <= _GEN_7487;
        end
      end else begin
        valid_133_1 <= _GEN_1672;
      end
    end else begin
      valid_133_1 <= _GEN_1672;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_134_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_134_0 <= _GEN_1161;
        end else begin
          valid_134_0 <= _GEN_7488;
        end
      end else begin
        valid_134_0 <= _GEN_1161;
      end
    end else begin
      valid_134_0 <= _GEN_1161;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_134_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_134_1 <= _GEN_1673;
        end else begin
          valid_134_1 <= _GEN_7489;
        end
      end else begin
        valid_134_1 <= _GEN_1673;
      end
    end else begin
      valid_134_1 <= _GEN_1673;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_135_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_135_0 <= _GEN_1162;
        end else begin
          valid_135_0 <= _GEN_7490;
        end
      end else begin
        valid_135_0 <= _GEN_1162;
      end
    end else begin
      valid_135_0 <= _GEN_1162;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_135_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_135_1 <= _GEN_1674;
        end else begin
          valid_135_1 <= _GEN_7491;
        end
      end else begin
        valid_135_1 <= _GEN_1674;
      end
    end else begin
      valid_135_1 <= _GEN_1674;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_136_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_136_0 <= _GEN_1163;
        end else begin
          valid_136_0 <= _GEN_7492;
        end
      end else begin
        valid_136_0 <= _GEN_1163;
      end
    end else begin
      valid_136_0 <= _GEN_1163;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_136_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_136_1 <= _GEN_1675;
        end else begin
          valid_136_1 <= _GEN_7493;
        end
      end else begin
        valid_136_1 <= _GEN_1675;
      end
    end else begin
      valid_136_1 <= _GEN_1675;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_137_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_137_0 <= _GEN_1164;
        end else begin
          valid_137_0 <= _GEN_7494;
        end
      end else begin
        valid_137_0 <= _GEN_1164;
      end
    end else begin
      valid_137_0 <= _GEN_1164;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_137_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_137_1 <= _GEN_1676;
        end else begin
          valid_137_1 <= _GEN_7495;
        end
      end else begin
        valid_137_1 <= _GEN_1676;
      end
    end else begin
      valid_137_1 <= _GEN_1676;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_138_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_138_0 <= _GEN_1165;
        end else begin
          valid_138_0 <= _GEN_7496;
        end
      end else begin
        valid_138_0 <= _GEN_1165;
      end
    end else begin
      valid_138_0 <= _GEN_1165;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_138_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_138_1 <= _GEN_1677;
        end else begin
          valid_138_1 <= _GEN_7497;
        end
      end else begin
        valid_138_1 <= _GEN_1677;
      end
    end else begin
      valid_138_1 <= _GEN_1677;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_139_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_139_0 <= _GEN_1166;
        end else begin
          valid_139_0 <= _GEN_7498;
        end
      end else begin
        valid_139_0 <= _GEN_1166;
      end
    end else begin
      valid_139_0 <= _GEN_1166;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_139_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_139_1 <= _GEN_1678;
        end else begin
          valid_139_1 <= _GEN_7499;
        end
      end else begin
        valid_139_1 <= _GEN_1678;
      end
    end else begin
      valid_139_1 <= _GEN_1678;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_140_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_140_0 <= _GEN_1167;
        end else begin
          valid_140_0 <= _GEN_7500;
        end
      end else begin
        valid_140_0 <= _GEN_1167;
      end
    end else begin
      valid_140_0 <= _GEN_1167;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_140_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_140_1 <= _GEN_1679;
        end else begin
          valid_140_1 <= _GEN_7501;
        end
      end else begin
        valid_140_1 <= _GEN_1679;
      end
    end else begin
      valid_140_1 <= _GEN_1679;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_141_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_141_0 <= _GEN_1168;
        end else begin
          valid_141_0 <= _GEN_7502;
        end
      end else begin
        valid_141_0 <= _GEN_1168;
      end
    end else begin
      valid_141_0 <= _GEN_1168;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_141_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_141_1 <= _GEN_1680;
        end else begin
          valid_141_1 <= _GEN_7503;
        end
      end else begin
        valid_141_1 <= _GEN_1680;
      end
    end else begin
      valid_141_1 <= _GEN_1680;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_142_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_142_0 <= _GEN_1169;
        end else begin
          valid_142_0 <= _GEN_7504;
        end
      end else begin
        valid_142_0 <= _GEN_1169;
      end
    end else begin
      valid_142_0 <= _GEN_1169;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_142_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_142_1 <= _GEN_1681;
        end else begin
          valid_142_1 <= _GEN_7505;
        end
      end else begin
        valid_142_1 <= _GEN_1681;
      end
    end else begin
      valid_142_1 <= _GEN_1681;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_143_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_143_0 <= _GEN_1170;
        end else begin
          valid_143_0 <= _GEN_7506;
        end
      end else begin
        valid_143_0 <= _GEN_1170;
      end
    end else begin
      valid_143_0 <= _GEN_1170;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_143_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_143_1 <= _GEN_1682;
        end else begin
          valid_143_1 <= _GEN_7507;
        end
      end else begin
        valid_143_1 <= _GEN_1682;
      end
    end else begin
      valid_143_1 <= _GEN_1682;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_144_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_144_0 <= _GEN_1171;
        end else begin
          valid_144_0 <= _GEN_7508;
        end
      end else begin
        valid_144_0 <= _GEN_1171;
      end
    end else begin
      valid_144_0 <= _GEN_1171;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_144_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_144_1 <= _GEN_1683;
        end else begin
          valid_144_1 <= _GEN_7509;
        end
      end else begin
        valid_144_1 <= _GEN_1683;
      end
    end else begin
      valid_144_1 <= _GEN_1683;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_145_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_145_0 <= _GEN_1172;
        end else begin
          valid_145_0 <= _GEN_7510;
        end
      end else begin
        valid_145_0 <= _GEN_1172;
      end
    end else begin
      valid_145_0 <= _GEN_1172;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_145_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_145_1 <= _GEN_1684;
        end else begin
          valid_145_1 <= _GEN_7511;
        end
      end else begin
        valid_145_1 <= _GEN_1684;
      end
    end else begin
      valid_145_1 <= _GEN_1684;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_146_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_146_0 <= _GEN_1173;
        end else begin
          valid_146_0 <= _GEN_7512;
        end
      end else begin
        valid_146_0 <= _GEN_1173;
      end
    end else begin
      valid_146_0 <= _GEN_1173;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_146_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_146_1 <= _GEN_1685;
        end else begin
          valid_146_1 <= _GEN_7513;
        end
      end else begin
        valid_146_1 <= _GEN_1685;
      end
    end else begin
      valid_146_1 <= _GEN_1685;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_147_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_147_0 <= _GEN_1174;
        end else begin
          valid_147_0 <= _GEN_7514;
        end
      end else begin
        valid_147_0 <= _GEN_1174;
      end
    end else begin
      valid_147_0 <= _GEN_1174;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_147_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_147_1 <= _GEN_1686;
        end else begin
          valid_147_1 <= _GEN_7515;
        end
      end else begin
        valid_147_1 <= _GEN_1686;
      end
    end else begin
      valid_147_1 <= _GEN_1686;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_148_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_148_0 <= _GEN_1175;
        end else begin
          valid_148_0 <= _GEN_7516;
        end
      end else begin
        valid_148_0 <= _GEN_1175;
      end
    end else begin
      valid_148_0 <= _GEN_1175;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_148_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_148_1 <= _GEN_1687;
        end else begin
          valid_148_1 <= _GEN_7517;
        end
      end else begin
        valid_148_1 <= _GEN_1687;
      end
    end else begin
      valid_148_1 <= _GEN_1687;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_149_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_149_0 <= _GEN_1176;
        end else begin
          valid_149_0 <= _GEN_7518;
        end
      end else begin
        valid_149_0 <= _GEN_1176;
      end
    end else begin
      valid_149_0 <= _GEN_1176;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_149_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_149_1 <= _GEN_1688;
        end else begin
          valid_149_1 <= _GEN_7519;
        end
      end else begin
        valid_149_1 <= _GEN_1688;
      end
    end else begin
      valid_149_1 <= _GEN_1688;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_150_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_150_0 <= _GEN_1177;
        end else begin
          valid_150_0 <= _GEN_7520;
        end
      end else begin
        valid_150_0 <= _GEN_1177;
      end
    end else begin
      valid_150_0 <= _GEN_1177;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_150_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_150_1 <= _GEN_1689;
        end else begin
          valid_150_1 <= _GEN_7521;
        end
      end else begin
        valid_150_1 <= _GEN_1689;
      end
    end else begin
      valid_150_1 <= _GEN_1689;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_151_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_151_0 <= _GEN_1178;
        end else begin
          valid_151_0 <= _GEN_7522;
        end
      end else begin
        valid_151_0 <= _GEN_1178;
      end
    end else begin
      valid_151_0 <= _GEN_1178;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_151_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_151_1 <= _GEN_1690;
        end else begin
          valid_151_1 <= _GEN_7523;
        end
      end else begin
        valid_151_1 <= _GEN_1690;
      end
    end else begin
      valid_151_1 <= _GEN_1690;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_152_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_152_0 <= _GEN_1179;
        end else begin
          valid_152_0 <= _GEN_7524;
        end
      end else begin
        valid_152_0 <= _GEN_1179;
      end
    end else begin
      valid_152_0 <= _GEN_1179;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_152_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_152_1 <= _GEN_1691;
        end else begin
          valid_152_1 <= _GEN_7525;
        end
      end else begin
        valid_152_1 <= _GEN_1691;
      end
    end else begin
      valid_152_1 <= _GEN_1691;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_153_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_153_0 <= _GEN_1180;
        end else begin
          valid_153_0 <= _GEN_7526;
        end
      end else begin
        valid_153_0 <= _GEN_1180;
      end
    end else begin
      valid_153_0 <= _GEN_1180;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_153_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_153_1 <= _GEN_1692;
        end else begin
          valid_153_1 <= _GEN_7527;
        end
      end else begin
        valid_153_1 <= _GEN_1692;
      end
    end else begin
      valid_153_1 <= _GEN_1692;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_154_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_154_0 <= _GEN_1181;
        end else begin
          valid_154_0 <= _GEN_7528;
        end
      end else begin
        valid_154_0 <= _GEN_1181;
      end
    end else begin
      valid_154_0 <= _GEN_1181;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_154_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_154_1 <= _GEN_1693;
        end else begin
          valid_154_1 <= _GEN_7529;
        end
      end else begin
        valid_154_1 <= _GEN_1693;
      end
    end else begin
      valid_154_1 <= _GEN_1693;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_155_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_155_0 <= _GEN_1182;
        end else begin
          valid_155_0 <= _GEN_7530;
        end
      end else begin
        valid_155_0 <= _GEN_1182;
      end
    end else begin
      valid_155_0 <= _GEN_1182;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_155_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_155_1 <= _GEN_1694;
        end else begin
          valid_155_1 <= _GEN_7531;
        end
      end else begin
        valid_155_1 <= _GEN_1694;
      end
    end else begin
      valid_155_1 <= _GEN_1694;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_156_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_156_0 <= _GEN_1183;
        end else begin
          valid_156_0 <= _GEN_7532;
        end
      end else begin
        valid_156_0 <= _GEN_1183;
      end
    end else begin
      valid_156_0 <= _GEN_1183;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_156_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_156_1 <= _GEN_1695;
        end else begin
          valid_156_1 <= _GEN_7533;
        end
      end else begin
        valid_156_1 <= _GEN_1695;
      end
    end else begin
      valid_156_1 <= _GEN_1695;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_157_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_157_0 <= _GEN_1184;
        end else begin
          valid_157_0 <= _GEN_7534;
        end
      end else begin
        valid_157_0 <= _GEN_1184;
      end
    end else begin
      valid_157_0 <= _GEN_1184;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_157_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_157_1 <= _GEN_1696;
        end else begin
          valid_157_1 <= _GEN_7535;
        end
      end else begin
        valid_157_1 <= _GEN_1696;
      end
    end else begin
      valid_157_1 <= _GEN_1696;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_158_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_158_0 <= _GEN_1185;
        end else begin
          valid_158_0 <= _GEN_7536;
        end
      end else begin
        valid_158_0 <= _GEN_1185;
      end
    end else begin
      valid_158_0 <= _GEN_1185;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_158_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_158_1 <= _GEN_1697;
        end else begin
          valid_158_1 <= _GEN_7537;
        end
      end else begin
        valid_158_1 <= _GEN_1697;
      end
    end else begin
      valid_158_1 <= _GEN_1697;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_159_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_159_0 <= _GEN_1186;
        end else begin
          valid_159_0 <= _GEN_7538;
        end
      end else begin
        valid_159_0 <= _GEN_1186;
      end
    end else begin
      valid_159_0 <= _GEN_1186;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_159_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_159_1 <= _GEN_1698;
        end else begin
          valid_159_1 <= _GEN_7539;
        end
      end else begin
        valid_159_1 <= _GEN_1698;
      end
    end else begin
      valid_159_1 <= _GEN_1698;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_160_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_160_0 <= _GEN_1187;
        end else begin
          valid_160_0 <= _GEN_7540;
        end
      end else begin
        valid_160_0 <= _GEN_1187;
      end
    end else begin
      valid_160_0 <= _GEN_1187;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_160_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_160_1 <= _GEN_1699;
        end else begin
          valid_160_1 <= _GEN_7541;
        end
      end else begin
        valid_160_1 <= _GEN_1699;
      end
    end else begin
      valid_160_1 <= _GEN_1699;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_161_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_161_0 <= _GEN_1188;
        end else begin
          valid_161_0 <= _GEN_7542;
        end
      end else begin
        valid_161_0 <= _GEN_1188;
      end
    end else begin
      valid_161_0 <= _GEN_1188;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_161_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_161_1 <= _GEN_1700;
        end else begin
          valid_161_1 <= _GEN_7543;
        end
      end else begin
        valid_161_1 <= _GEN_1700;
      end
    end else begin
      valid_161_1 <= _GEN_1700;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_162_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_162_0 <= _GEN_1189;
        end else begin
          valid_162_0 <= _GEN_7544;
        end
      end else begin
        valid_162_0 <= _GEN_1189;
      end
    end else begin
      valid_162_0 <= _GEN_1189;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_162_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_162_1 <= _GEN_1701;
        end else begin
          valid_162_1 <= _GEN_7545;
        end
      end else begin
        valid_162_1 <= _GEN_1701;
      end
    end else begin
      valid_162_1 <= _GEN_1701;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_163_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_163_0 <= _GEN_1190;
        end else begin
          valid_163_0 <= _GEN_7546;
        end
      end else begin
        valid_163_0 <= _GEN_1190;
      end
    end else begin
      valid_163_0 <= _GEN_1190;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_163_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_163_1 <= _GEN_1702;
        end else begin
          valid_163_1 <= _GEN_7547;
        end
      end else begin
        valid_163_1 <= _GEN_1702;
      end
    end else begin
      valid_163_1 <= _GEN_1702;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_164_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_164_0 <= _GEN_1191;
        end else begin
          valid_164_0 <= _GEN_7548;
        end
      end else begin
        valid_164_0 <= _GEN_1191;
      end
    end else begin
      valid_164_0 <= _GEN_1191;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_164_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_164_1 <= _GEN_1703;
        end else begin
          valid_164_1 <= _GEN_7549;
        end
      end else begin
        valid_164_1 <= _GEN_1703;
      end
    end else begin
      valid_164_1 <= _GEN_1703;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_165_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_165_0 <= _GEN_1192;
        end else begin
          valid_165_0 <= _GEN_7550;
        end
      end else begin
        valid_165_0 <= _GEN_1192;
      end
    end else begin
      valid_165_0 <= _GEN_1192;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_165_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_165_1 <= _GEN_1704;
        end else begin
          valid_165_1 <= _GEN_7551;
        end
      end else begin
        valid_165_1 <= _GEN_1704;
      end
    end else begin
      valid_165_1 <= _GEN_1704;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_166_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_166_0 <= _GEN_1193;
        end else begin
          valid_166_0 <= _GEN_7552;
        end
      end else begin
        valid_166_0 <= _GEN_1193;
      end
    end else begin
      valid_166_0 <= _GEN_1193;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_166_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_166_1 <= _GEN_1705;
        end else begin
          valid_166_1 <= _GEN_7553;
        end
      end else begin
        valid_166_1 <= _GEN_1705;
      end
    end else begin
      valid_166_1 <= _GEN_1705;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_167_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_167_0 <= _GEN_1194;
        end else begin
          valid_167_0 <= _GEN_7554;
        end
      end else begin
        valid_167_0 <= _GEN_1194;
      end
    end else begin
      valid_167_0 <= _GEN_1194;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_167_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_167_1 <= _GEN_1706;
        end else begin
          valid_167_1 <= _GEN_7555;
        end
      end else begin
        valid_167_1 <= _GEN_1706;
      end
    end else begin
      valid_167_1 <= _GEN_1706;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_168_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_168_0 <= _GEN_1195;
        end else begin
          valid_168_0 <= _GEN_7556;
        end
      end else begin
        valid_168_0 <= _GEN_1195;
      end
    end else begin
      valid_168_0 <= _GEN_1195;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_168_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_168_1 <= _GEN_1707;
        end else begin
          valid_168_1 <= _GEN_7557;
        end
      end else begin
        valid_168_1 <= _GEN_1707;
      end
    end else begin
      valid_168_1 <= _GEN_1707;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_169_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_169_0 <= _GEN_1196;
        end else begin
          valid_169_0 <= _GEN_7558;
        end
      end else begin
        valid_169_0 <= _GEN_1196;
      end
    end else begin
      valid_169_0 <= _GEN_1196;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_169_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_169_1 <= _GEN_1708;
        end else begin
          valid_169_1 <= _GEN_7559;
        end
      end else begin
        valid_169_1 <= _GEN_1708;
      end
    end else begin
      valid_169_1 <= _GEN_1708;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_170_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_170_0 <= _GEN_1197;
        end else begin
          valid_170_0 <= _GEN_7560;
        end
      end else begin
        valid_170_0 <= _GEN_1197;
      end
    end else begin
      valid_170_0 <= _GEN_1197;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_170_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_170_1 <= _GEN_1709;
        end else begin
          valid_170_1 <= _GEN_7561;
        end
      end else begin
        valid_170_1 <= _GEN_1709;
      end
    end else begin
      valid_170_1 <= _GEN_1709;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_171_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_171_0 <= _GEN_1198;
        end else begin
          valid_171_0 <= _GEN_7562;
        end
      end else begin
        valid_171_0 <= _GEN_1198;
      end
    end else begin
      valid_171_0 <= _GEN_1198;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_171_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_171_1 <= _GEN_1710;
        end else begin
          valid_171_1 <= _GEN_7563;
        end
      end else begin
        valid_171_1 <= _GEN_1710;
      end
    end else begin
      valid_171_1 <= _GEN_1710;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_172_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_172_0 <= _GEN_1199;
        end else begin
          valid_172_0 <= _GEN_7564;
        end
      end else begin
        valid_172_0 <= _GEN_1199;
      end
    end else begin
      valid_172_0 <= _GEN_1199;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_172_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_172_1 <= _GEN_1711;
        end else begin
          valid_172_1 <= _GEN_7565;
        end
      end else begin
        valid_172_1 <= _GEN_1711;
      end
    end else begin
      valid_172_1 <= _GEN_1711;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_173_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_173_0 <= _GEN_1200;
        end else begin
          valid_173_0 <= _GEN_7566;
        end
      end else begin
        valid_173_0 <= _GEN_1200;
      end
    end else begin
      valid_173_0 <= _GEN_1200;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_173_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_173_1 <= _GEN_1712;
        end else begin
          valid_173_1 <= _GEN_7567;
        end
      end else begin
        valid_173_1 <= _GEN_1712;
      end
    end else begin
      valid_173_1 <= _GEN_1712;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_174_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_174_0 <= _GEN_1201;
        end else begin
          valid_174_0 <= _GEN_7568;
        end
      end else begin
        valid_174_0 <= _GEN_1201;
      end
    end else begin
      valid_174_0 <= _GEN_1201;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_174_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_174_1 <= _GEN_1713;
        end else begin
          valid_174_1 <= _GEN_7569;
        end
      end else begin
        valid_174_1 <= _GEN_1713;
      end
    end else begin
      valid_174_1 <= _GEN_1713;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_175_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_175_0 <= _GEN_1202;
        end else begin
          valid_175_0 <= _GEN_7570;
        end
      end else begin
        valid_175_0 <= _GEN_1202;
      end
    end else begin
      valid_175_0 <= _GEN_1202;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_175_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_175_1 <= _GEN_1714;
        end else begin
          valid_175_1 <= _GEN_7571;
        end
      end else begin
        valid_175_1 <= _GEN_1714;
      end
    end else begin
      valid_175_1 <= _GEN_1714;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_176_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_176_0 <= _GEN_1203;
        end else begin
          valid_176_0 <= _GEN_7572;
        end
      end else begin
        valid_176_0 <= _GEN_1203;
      end
    end else begin
      valid_176_0 <= _GEN_1203;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_176_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_176_1 <= _GEN_1715;
        end else begin
          valid_176_1 <= _GEN_7573;
        end
      end else begin
        valid_176_1 <= _GEN_1715;
      end
    end else begin
      valid_176_1 <= _GEN_1715;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_177_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_177_0 <= _GEN_1204;
        end else begin
          valid_177_0 <= _GEN_7574;
        end
      end else begin
        valid_177_0 <= _GEN_1204;
      end
    end else begin
      valid_177_0 <= _GEN_1204;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_177_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_177_1 <= _GEN_1716;
        end else begin
          valid_177_1 <= _GEN_7575;
        end
      end else begin
        valid_177_1 <= _GEN_1716;
      end
    end else begin
      valid_177_1 <= _GEN_1716;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_178_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_178_0 <= _GEN_1205;
        end else begin
          valid_178_0 <= _GEN_7576;
        end
      end else begin
        valid_178_0 <= _GEN_1205;
      end
    end else begin
      valid_178_0 <= _GEN_1205;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_178_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_178_1 <= _GEN_1717;
        end else begin
          valid_178_1 <= _GEN_7577;
        end
      end else begin
        valid_178_1 <= _GEN_1717;
      end
    end else begin
      valid_178_1 <= _GEN_1717;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_179_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_179_0 <= _GEN_1206;
        end else begin
          valid_179_0 <= _GEN_7578;
        end
      end else begin
        valid_179_0 <= _GEN_1206;
      end
    end else begin
      valid_179_0 <= _GEN_1206;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_179_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_179_1 <= _GEN_1718;
        end else begin
          valid_179_1 <= _GEN_7579;
        end
      end else begin
        valid_179_1 <= _GEN_1718;
      end
    end else begin
      valid_179_1 <= _GEN_1718;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_180_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_180_0 <= _GEN_1207;
        end else begin
          valid_180_0 <= _GEN_7580;
        end
      end else begin
        valid_180_0 <= _GEN_1207;
      end
    end else begin
      valid_180_0 <= _GEN_1207;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_180_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_180_1 <= _GEN_1719;
        end else begin
          valid_180_1 <= _GEN_7581;
        end
      end else begin
        valid_180_1 <= _GEN_1719;
      end
    end else begin
      valid_180_1 <= _GEN_1719;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_181_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_181_0 <= _GEN_1208;
        end else begin
          valid_181_0 <= _GEN_7582;
        end
      end else begin
        valid_181_0 <= _GEN_1208;
      end
    end else begin
      valid_181_0 <= _GEN_1208;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_181_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_181_1 <= _GEN_1720;
        end else begin
          valid_181_1 <= _GEN_7583;
        end
      end else begin
        valid_181_1 <= _GEN_1720;
      end
    end else begin
      valid_181_1 <= _GEN_1720;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_182_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_182_0 <= _GEN_1209;
        end else begin
          valid_182_0 <= _GEN_7584;
        end
      end else begin
        valid_182_0 <= _GEN_1209;
      end
    end else begin
      valid_182_0 <= _GEN_1209;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_182_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_182_1 <= _GEN_1721;
        end else begin
          valid_182_1 <= _GEN_7585;
        end
      end else begin
        valid_182_1 <= _GEN_1721;
      end
    end else begin
      valid_182_1 <= _GEN_1721;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_183_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_183_0 <= _GEN_1210;
        end else begin
          valid_183_0 <= _GEN_7586;
        end
      end else begin
        valid_183_0 <= _GEN_1210;
      end
    end else begin
      valid_183_0 <= _GEN_1210;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_183_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_183_1 <= _GEN_1722;
        end else begin
          valid_183_1 <= _GEN_7587;
        end
      end else begin
        valid_183_1 <= _GEN_1722;
      end
    end else begin
      valid_183_1 <= _GEN_1722;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_184_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_184_0 <= _GEN_1211;
        end else begin
          valid_184_0 <= _GEN_7588;
        end
      end else begin
        valid_184_0 <= _GEN_1211;
      end
    end else begin
      valid_184_0 <= _GEN_1211;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_184_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_184_1 <= _GEN_1723;
        end else begin
          valid_184_1 <= _GEN_7589;
        end
      end else begin
        valid_184_1 <= _GEN_1723;
      end
    end else begin
      valid_184_1 <= _GEN_1723;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_185_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_185_0 <= _GEN_1212;
        end else begin
          valid_185_0 <= _GEN_7590;
        end
      end else begin
        valid_185_0 <= _GEN_1212;
      end
    end else begin
      valid_185_0 <= _GEN_1212;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_185_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_185_1 <= _GEN_1724;
        end else begin
          valid_185_1 <= _GEN_7591;
        end
      end else begin
        valid_185_1 <= _GEN_1724;
      end
    end else begin
      valid_185_1 <= _GEN_1724;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_186_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_186_0 <= _GEN_1213;
        end else begin
          valid_186_0 <= _GEN_7592;
        end
      end else begin
        valid_186_0 <= _GEN_1213;
      end
    end else begin
      valid_186_0 <= _GEN_1213;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_186_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_186_1 <= _GEN_1725;
        end else begin
          valid_186_1 <= _GEN_7593;
        end
      end else begin
        valid_186_1 <= _GEN_1725;
      end
    end else begin
      valid_186_1 <= _GEN_1725;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_187_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_187_0 <= _GEN_1214;
        end else begin
          valid_187_0 <= _GEN_7594;
        end
      end else begin
        valid_187_0 <= _GEN_1214;
      end
    end else begin
      valid_187_0 <= _GEN_1214;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_187_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_187_1 <= _GEN_1726;
        end else begin
          valid_187_1 <= _GEN_7595;
        end
      end else begin
        valid_187_1 <= _GEN_1726;
      end
    end else begin
      valid_187_1 <= _GEN_1726;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_188_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_188_0 <= _GEN_1215;
        end else begin
          valid_188_0 <= _GEN_7596;
        end
      end else begin
        valid_188_0 <= _GEN_1215;
      end
    end else begin
      valid_188_0 <= _GEN_1215;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_188_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_188_1 <= _GEN_1727;
        end else begin
          valid_188_1 <= _GEN_7597;
        end
      end else begin
        valid_188_1 <= _GEN_1727;
      end
    end else begin
      valid_188_1 <= _GEN_1727;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_189_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_189_0 <= _GEN_1216;
        end else begin
          valid_189_0 <= _GEN_7598;
        end
      end else begin
        valid_189_0 <= _GEN_1216;
      end
    end else begin
      valid_189_0 <= _GEN_1216;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_189_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_189_1 <= _GEN_1728;
        end else begin
          valid_189_1 <= _GEN_7599;
        end
      end else begin
        valid_189_1 <= _GEN_1728;
      end
    end else begin
      valid_189_1 <= _GEN_1728;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_190_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_190_0 <= _GEN_1217;
        end else begin
          valid_190_0 <= _GEN_7600;
        end
      end else begin
        valid_190_0 <= _GEN_1217;
      end
    end else begin
      valid_190_0 <= _GEN_1217;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_190_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_190_1 <= _GEN_1729;
        end else begin
          valid_190_1 <= _GEN_7601;
        end
      end else begin
        valid_190_1 <= _GEN_1729;
      end
    end else begin
      valid_190_1 <= _GEN_1729;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_191_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_191_0 <= _GEN_1218;
        end else begin
          valid_191_0 <= _GEN_7602;
        end
      end else begin
        valid_191_0 <= _GEN_1218;
      end
    end else begin
      valid_191_0 <= _GEN_1218;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_191_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_191_1 <= _GEN_1730;
        end else begin
          valid_191_1 <= _GEN_7603;
        end
      end else begin
        valid_191_1 <= _GEN_1730;
      end
    end else begin
      valid_191_1 <= _GEN_1730;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_192_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_192_0 <= _GEN_1219;
        end else begin
          valid_192_0 <= _GEN_7604;
        end
      end else begin
        valid_192_0 <= _GEN_1219;
      end
    end else begin
      valid_192_0 <= _GEN_1219;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_192_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_192_1 <= _GEN_1731;
        end else begin
          valid_192_1 <= _GEN_7605;
        end
      end else begin
        valid_192_1 <= _GEN_1731;
      end
    end else begin
      valid_192_1 <= _GEN_1731;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_193_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_193_0 <= _GEN_1220;
        end else begin
          valid_193_0 <= _GEN_7606;
        end
      end else begin
        valid_193_0 <= _GEN_1220;
      end
    end else begin
      valid_193_0 <= _GEN_1220;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_193_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_193_1 <= _GEN_1732;
        end else begin
          valid_193_1 <= _GEN_7607;
        end
      end else begin
        valid_193_1 <= _GEN_1732;
      end
    end else begin
      valid_193_1 <= _GEN_1732;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_194_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_194_0 <= _GEN_1221;
        end else begin
          valid_194_0 <= _GEN_7608;
        end
      end else begin
        valid_194_0 <= _GEN_1221;
      end
    end else begin
      valid_194_0 <= _GEN_1221;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_194_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_194_1 <= _GEN_1733;
        end else begin
          valid_194_1 <= _GEN_7609;
        end
      end else begin
        valid_194_1 <= _GEN_1733;
      end
    end else begin
      valid_194_1 <= _GEN_1733;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_195_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_195_0 <= _GEN_1222;
        end else begin
          valid_195_0 <= _GEN_7610;
        end
      end else begin
        valid_195_0 <= _GEN_1222;
      end
    end else begin
      valid_195_0 <= _GEN_1222;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_195_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_195_1 <= _GEN_1734;
        end else begin
          valid_195_1 <= _GEN_7611;
        end
      end else begin
        valid_195_1 <= _GEN_1734;
      end
    end else begin
      valid_195_1 <= _GEN_1734;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_196_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_196_0 <= _GEN_1223;
        end else begin
          valid_196_0 <= _GEN_7612;
        end
      end else begin
        valid_196_0 <= _GEN_1223;
      end
    end else begin
      valid_196_0 <= _GEN_1223;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_196_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_196_1 <= _GEN_1735;
        end else begin
          valid_196_1 <= _GEN_7613;
        end
      end else begin
        valid_196_1 <= _GEN_1735;
      end
    end else begin
      valid_196_1 <= _GEN_1735;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_197_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_197_0 <= _GEN_1224;
        end else begin
          valid_197_0 <= _GEN_7614;
        end
      end else begin
        valid_197_0 <= _GEN_1224;
      end
    end else begin
      valid_197_0 <= _GEN_1224;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_197_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_197_1 <= _GEN_1736;
        end else begin
          valid_197_1 <= _GEN_7615;
        end
      end else begin
        valid_197_1 <= _GEN_1736;
      end
    end else begin
      valid_197_1 <= _GEN_1736;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_198_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_198_0 <= _GEN_1225;
        end else begin
          valid_198_0 <= _GEN_7616;
        end
      end else begin
        valid_198_0 <= _GEN_1225;
      end
    end else begin
      valid_198_0 <= _GEN_1225;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_198_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_198_1 <= _GEN_1737;
        end else begin
          valid_198_1 <= _GEN_7617;
        end
      end else begin
        valid_198_1 <= _GEN_1737;
      end
    end else begin
      valid_198_1 <= _GEN_1737;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_199_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_199_0 <= _GEN_1226;
        end else begin
          valid_199_0 <= _GEN_7618;
        end
      end else begin
        valid_199_0 <= _GEN_1226;
      end
    end else begin
      valid_199_0 <= _GEN_1226;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_199_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_199_1 <= _GEN_1738;
        end else begin
          valid_199_1 <= _GEN_7619;
        end
      end else begin
        valid_199_1 <= _GEN_1738;
      end
    end else begin
      valid_199_1 <= _GEN_1738;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_200_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_200_0 <= _GEN_1227;
        end else begin
          valid_200_0 <= _GEN_7620;
        end
      end else begin
        valid_200_0 <= _GEN_1227;
      end
    end else begin
      valid_200_0 <= _GEN_1227;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_200_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_200_1 <= _GEN_1739;
        end else begin
          valid_200_1 <= _GEN_7621;
        end
      end else begin
        valid_200_1 <= _GEN_1739;
      end
    end else begin
      valid_200_1 <= _GEN_1739;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_201_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_201_0 <= _GEN_1228;
        end else begin
          valid_201_0 <= _GEN_7622;
        end
      end else begin
        valid_201_0 <= _GEN_1228;
      end
    end else begin
      valid_201_0 <= _GEN_1228;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_201_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_201_1 <= _GEN_1740;
        end else begin
          valid_201_1 <= _GEN_7623;
        end
      end else begin
        valid_201_1 <= _GEN_1740;
      end
    end else begin
      valid_201_1 <= _GEN_1740;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_202_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_202_0 <= _GEN_1229;
        end else begin
          valid_202_0 <= _GEN_7624;
        end
      end else begin
        valid_202_0 <= _GEN_1229;
      end
    end else begin
      valid_202_0 <= _GEN_1229;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_202_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_202_1 <= _GEN_1741;
        end else begin
          valid_202_1 <= _GEN_7625;
        end
      end else begin
        valid_202_1 <= _GEN_1741;
      end
    end else begin
      valid_202_1 <= _GEN_1741;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_203_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_203_0 <= _GEN_1230;
        end else begin
          valid_203_0 <= _GEN_7626;
        end
      end else begin
        valid_203_0 <= _GEN_1230;
      end
    end else begin
      valid_203_0 <= _GEN_1230;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_203_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_203_1 <= _GEN_1742;
        end else begin
          valid_203_1 <= _GEN_7627;
        end
      end else begin
        valid_203_1 <= _GEN_1742;
      end
    end else begin
      valid_203_1 <= _GEN_1742;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_204_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_204_0 <= _GEN_1231;
        end else begin
          valid_204_0 <= _GEN_7628;
        end
      end else begin
        valid_204_0 <= _GEN_1231;
      end
    end else begin
      valid_204_0 <= _GEN_1231;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_204_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_204_1 <= _GEN_1743;
        end else begin
          valid_204_1 <= _GEN_7629;
        end
      end else begin
        valid_204_1 <= _GEN_1743;
      end
    end else begin
      valid_204_1 <= _GEN_1743;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_205_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_205_0 <= _GEN_1232;
        end else begin
          valid_205_0 <= _GEN_7630;
        end
      end else begin
        valid_205_0 <= _GEN_1232;
      end
    end else begin
      valid_205_0 <= _GEN_1232;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_205_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_205_1 <= _GEN_1744;
        end else begin
          valid_205_1 <= _GEN_7631;
        end
      end else begin
        valid_205_1 <= _GEN_1744;
      end
    end else begin
      valid_205_1 <= _GEN_1744;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_206_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_206_0 <= _GEN_1233;
        end else begin
          valid_206_0 <= _GEN_7632;
        end
      end else begin
        valid_206_0 <= _GEN_1233;
      end
    end else begin
      valid_206_0 <= _GEN_1233;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_206_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_206_1 <= _GEN_1745;
        end else begin
          valid_206_1 <= _GEN_7633;
        end
      end else begin
        valid_206_1 <= _GEN_1745;
      end
    end else begin
      valid_206_1 <= _GEN_1745;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_207_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_207_0 <= _GEN_1234;
        end else begin
          valid_207_0 <= _GEN_7634;
        end
      end else begin
        valid_207_0 <= _GEN_1234;
      end
    end else begin
      valid_207_0 <= _GEN_1234;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_207_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_207_1 <= _GEN_1746;
        end else begin
          valid_207_1 <= _GEN_7635;
        end
      end else begin
        valid_207_1 <= _GEN_1746;
      end
    end else begin
      valid_207_1 <= _GEN_1746;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_208_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_208_0 <= _GEN_1235;
        end else begin
          valid_208_0 <= _GEN_7636;
        end
      end else begin
        valid_208_0 <= _GEN_1235;
      end
    end else begin
      valid_208_0 <= _GEN_1235;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_208_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_208_1 <= _GEN_1747;
        end else begin
          valid_208_1 <= _GEN_7637;
        end
      end else begin
        valid_208_1 <= _GEN_1747;
      end
    end else begin
      valid_208_1 <= _GEN_1747;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_209_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_209_0 <= _GEN_1236;
        end else begin
          valid_209_0 <= _GEN_7638;
        end
      end else begin
        valid_209_0 <= _GEN_1236;
      end
    end else begin
      valid_209_0 <= _GEN_1236;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_209_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_209_1 <= _GEN_1748;
        end else begin
          valid_209_1 <= _GEN_7639;
        end
      end else begin
        valid_209_1 <= _GEN_1748;
      end
    end else begin
      valid_209_1 <= _GEN_1748;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_210_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_210_0 <= _GEN_1237;
        end else begin
          valid_210_0 <= _GEN_7640;
        end
      end else begin
        valid_210_0 <= _GEN_1237;
      end
    end else begin
      valid_210_0 <= _GEN_1237;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_210_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_210_1 <= _GEN_1749;
        end else begin
          valid_210_1 <= _GEN_7641;
        end
      end else begin
        valid_210_1 <= _GEN_1749;
      end
    end else begin
      valid_210_1 <= _GEN_1749;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_211_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_211_0 <= _GEN_1238;
        end else begin
          valid_211_0 <= _GEN_7642;
        end
      end else begin
        valid_211_0 <= _GEN_1238;
      end
    end else begin
      valid_211_0 <= _GEN_1238;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_211_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_211_1 <= _GEN_1750;
        end else begin
          valid_211_1 <= _GEN_7643;
        end
      end else begin
        valid_211_1 <= _GEN_1750;
      end
    end else begin
      valid_211_1 <= _GEN_1750;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_212_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_212_0 <= _GEN_1239;
        end else begin
          valid_212_0 <= _GEN_7644;
        end
      end else begin
        valid_212_0 <= _GEN_1239;
      end
    end else begin
      valid_212_0 <= _GEN_1239;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_212_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_212_1 <= _GEN_1751;
        end else begin
          valid_212_1 <= _GEN_7645;
        end
      end else begin
        valid_212_1 <= _GEN_1751;
      end
    end else begin
      valid_212_1 <= _GEN_1751;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_213_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_213_0 <= _GEN_1240;
        end else begin
          valid_213_0 <= _GEN_7646;
        end
      end else begin
        valid_213_0 <= _GEN_1240;
      end
    end else begin
      valid_213_0 <= _GEN_1240;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_213_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_213_1 <= _GEN_1752;
        end else begin
          valid_213_1 <= _GEN_7647;
        end
      end else begin
        valid_213_1 <= _GEN_1752;
      end
    end else begin
      valid_213_1 <= _GEN_1752;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_214_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_214_0 <= _GEN_1241;
        end else begin
          valid_214_0 <= _GEN_7648;
        end
      end else begin
        valid_214_0 <= _GEN_1241;
      end
    end else begin
      valid_214_0 <= _GEN_1241;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_214_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_214_1 <= _GEN_1753;
        end else begin
          valid_214_1 <= _GEN_7649;
        end
      end else begin
        valid_214_1 <= _GEN_1753;
      end
    end else begin
      valid_214_1 <= _GEN_1753;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_215_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_215_0 <= _GEN_1242;
        end else begin
          valid_215_0 <= _GEN_7650;
        end
      end else begin
        valid_215_0 <= _GEN_1242;
      end
    end else begin
      valid_215_0 <= _GEN_1242;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_215_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_215_1 <= _GEN_1754;
        end else begin
          valid_215_1 <= _GEN_7651;
        end
      end else begin
        valid_215_1 <= _GEN_1754;
      end
    end else begin
      valid_215_1 <= _GEN_1754;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_216_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_216_0 <= _GEN_1243;
        end else begin
          valid_216_0 <= _GEN_7652;
        end
      end else begin
        valid_216_0 <= _GEN_1243;
      end
    end else begin
      valid_216_0 <= _GEN_1243;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_216_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_216_1 <= _GEN_1755;
        end else begin
          valid_216_1 <= _GEN_7653;
        end
      end else begin
        valid_216_1 <= _GEN_1755;
      end
    end else begin
      valid_216_1 <= _GEN_1755;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_217_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_217_0 <= _GEN_1244;
        end else begin
          valid_217_0 <= _GEN_7654;
        end
      end else begin
        valid_217_0 <= _GEN_1244;
      end
    end else begin
      valid_217_0 <= _GEN_1244;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_217_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_217_1 <= _GEN_1756;
        end else begin
          valid_217_1 <= _GEN_7655;
        end
      end else begin
        valid_217_1 <= _GEN_1756;
      end
    end else begin
      valid_217_1 <= _GEN_1756;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_218_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_218_0 <= _GEN_1245;
        end else begin
          valid_218_0 <= _GEN_7656;
        end
      end else begin
        valid_218_0 <= _GEN_1245;
      end
    end else begin
      valid_218_0 <= _GEN_1245;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_218_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_218_1 <= _GEN_1757;
        end else begin
          valid_218_1 <= _GEN_7657;
        end
      end else begin
        valid_218_1 <= _GEN_1757;
      end
    end else begin
      valid_218_1 <= _GEN_1757;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_219_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_219_0 <= _GEN_1246;
        end else begin
          valid_219_0 <= _GEN_7658;
        end
      end else begin
        valid_219_0 <= _GEN_1246;
      end
    end else begin
      valid_219_0 <= _GEN_1246;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_219_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_219_1 <= _GEN_1758;
        end else begin
          valid_219_1 <= _GEN_7659;
        end
      end else begin
        valid_219_1 <= _GEN_1758;
      end
    end else begin
      valid_219_1 <= _GEN_1758;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_220_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_220_0 <= _GEN_1247;
        end else begin
          valid_220_0 <= _GEN_7660;
        end
      end else begin
        valid_220_0 <= _GEN_1247;
      end
    end else begin
      valid_220_0 <= _GEN_1247;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_220_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_220_1 <= _GEN_1759;
        end else begin
          valid_220_1 <= _GEN_7661;
        end
      end else begin
        valid_220_1 <= _GEN_1759;
      end
    end else begin
      valid_220_1 <= _GEN_1759;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_221_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_221_0 <= _GEN_1248;
        end else begin
          valid_221_0 <= _GEN_7662;
        end
      end else begin
        valid_221_0 <= _GEN_1248;
      end
    end else begin
      valid_221_0 <= _GEN_1248;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_221_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_221_1 <= _GEN_1760;
        end else begin
          valid_221_1 <= _GEN_7663;
        end
      end else begin
        valid_221_1 <= _GEN_1760;
      end
    end else begin
      valid_221_1 <= _GEN_1760;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_222_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_222_0 <= _GEN_1249;
        end else begin
          valid_222_0 <= _GEN_7664;
        end
      end else begin
        valid_222_0 <= _GEN_1249;
      end
    end else begin
      valid_222_0 <= _GEN_1249;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_222_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_222_1 <= _GEN_1761;
        end else begin
          valid_222_1 <= _GEN_7665;
        end
      end else begin
        valid_222_1 <= _GEN_1761;
      end
    end else begin
      valid_222_1 <= _GEN_1761;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_223_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_223_0 <= _GEN_1250;
        end else begin
          valid_223_0 <= _GEN_7666;
        end
      end else begin
        valid_223_0 <= _GEN_1250;
      end
    end else begin
      valid_223_0 <= _GEN_1250;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_223_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_223_1 <= _GEN_1762;
        end else begin
          valid_223_1 <= _GEN_7667;
        end
      end else begin
        valid_223_1 <= _GEN_1762;
      end
    end else begin
      valid_223_1 <= _GEN_1762;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_224_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_224_0 <= _GEN_1251;
        end else begin
          valid_224_0 <= _GEN_7668;
        end
      end else begin
        valid_224_0 <= _GEN_1251;
      end
    end else begin
      valid_224_0 <= _GEN_1251;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_224_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_224_1 <= _GEN_1763;
        end else begin
          valid_224_1 <= _GEN_7669;
        end
      end else begin
        valid_224_1 <= _GEN_1763;
      end
    end else begin
      valid_224_1 <= _GEN_1763;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_225_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_225_0 <= _GEN_1252;
        end else begin
          valid_225_0 <= _GEN_7670;
        end
      end else begin
        valid_225_0 <= _GEN_1252;
      end
    end else begin
      valid_225_0 <= _GEN_1252;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_225_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_225_1 <= _GEN_1764;
        end else begin
          valid_225_1 <= _GEN_7671;
        end
      end else begin
        valid_225_1 <= _GEN_1764;
      end
    end else begin
      valid_225_1 <= _GEN_1764;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_226_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_226_0 <= _GEN_1253;
        end else begin
          valid_226_0 <= _GEN_7672;
        end
      end else begin
        valid_226_0 <= _GEN_1253;
      end
    end else begin
      valid_226_0 <= _GEN_1253;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_226_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_226_1 <= _GEN_1765;
        end else begin
          valid_226_1 <= _GEN_7673;
        end
      end else begin
        valid_226_1 <= _GEN_1765;
      end
    end else begin
      valid_226_1 <= _GEN_1765;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_227_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_227_0 <= _GEN_1254;
        end else begin
          valid_227_0 <= _GEN_7674;
        end
      end else begin
        valid_227_0 <= _GEN_1254;
      end
    end else begin
      valid_227_0 <= _GEN_1254;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_227_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_227_1 <= _GEN_1766;
        end else begin
          valid_227_1 <= _GEN_7675;
        end
      end else begin
        valid_227_1 <= _GEN_1766;
      end
    end else begin
      valid_227_1 <= _GEN_1766;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_228_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_228_0 <= _GEN_1255;
        end else begin
          valid_228_0 <= _GEN_7676;
        end
      end else begin
        valid_228_0 <= _GEN_1255;
      end
    end else begin
      valid_228_0 <= _GEN_1255;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_228_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_228_1 <= _GEN_1767;
        end else begin
          valid_228_1 <= _GEN_7677;
        end
      end else begin
        valid_228_1 <= _GEN_1767;
      end
    end else begin
      valid_228_1 <= _GEN_1767;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_229_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_229_0 <= _GEN_1256;
        end else begin
          valid_229_0 <= _GEN_7678;
        end
      end else begin
        valid_229_0 <= _GEN_1256;
      end
    end else begin
      valid_229_0 <= _GEN_1256;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_229_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_229_1 <= _GEN_1768;
        end else begin
          valid_229_1 <= _GEN_7679;
        end
      end else begin
        valid_229_1 <= _GEN_1768;
      end
    end else begin
      valid_229_1 <= _GEN_1768;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_230_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_230_0 <= _GEN_1257;
        end else begin
          valid_230_0 <= _GEN_7680;
        end
      end else begin
        valid_230_0 <= _GEN_1257;
      end
    end else begin
      valid_230_0 <= _GEN_1257;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_230_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_230_1 <= _GEN_1769;
        end else begin
          valid_230_1 <= _GEN_7681;
        end
      end else begin
        valid_230_1 <= _GEN_1769;
      end
    end else begin
      valid_230_1 <= _GEN_1769;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_231_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_231_0 <= _GEN_1258;
        end else begin
          valid_231_0 <= _GEN_7682;
        end
      end else begin
        valid_231_0 <= _GEN_1258;
      end
    end else begin
      valid_231_0 <= _GEN_1258;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_231_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_231_1 <= _GEN_1770;
        end else begin
          valid_231_1 <= _GEN_7683;
        end
      end else begin
        valid_231_1 <= _GEN_1770;
      end
    end else begin
      valid_231_1 <= _GEN_1770;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_232_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_232_0 <= _GEN_1259;
        end else begin
          valid_232_0 <= _GEN_7684;
        end
      end else begin
        valid_232_0 <= _GEN_1259;
      end
    end else begin
      valid_232_0 <= _GEN_1259;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_232_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_232_1 <= _GEN_1771;
        end else begin
          valid_232_1 <= _GEN_7685;
        end
      end else begin
        valid_232_1 <= _GEN_1771;
      end
    end else begin
      valid_232_1 <= _GEN_1771;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_233_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_233_0 <= _GEN_1260;
        end else begin
          valid_233_0 <= _GEN_7686;
        end
      end else begin
        valid_233_0 <= _GEN_1260;
      end
    end else begin
      valid_233_0 <= _GEN_1260;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_233_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_233_1 <= _GEN_1772;
        end else begin
          valid_233_1 <= _GEN_7687;
        end
      end else begin
        valid_233_1 <= _GEN_1772;
      end
    end else begin
      valid_233_1 <= _GEN_1772;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_234_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_234_0 <= _GEN_1261;
        end else begin
          valid_234_0 <= _GEN_7688;
        end
      end else begin
        valid_234_0 <= _GEN_1261;
      end
    end else begin
      valid_234_0 <= _GEN_1261;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_234_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_234_1 <= _GEN_1773;
        end else begin
          valid_234_1 <= _GEN_7689;
        end
      end else begin
        valid_234_1 <= _GEN_1773;
      end
    end else begin
      valid_234_1 <= _GEN_1773;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_235_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_235_0 <= _GEN_1262;
        end else begin
          valid_235_0 <= _GEN_7690;
        end
      end else begin
        valid_235_0 <= _GEN_1262;
      end
    end else begin
      valid_235_0 <= _GEN_1262;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_235_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_235_1 <= _GEN_1774;
        end else begin
          valid_235_1 <= _GEN_7691;
        end
      end else begin
        valid_235_1 <= _GEN_1774;
      end
    end else begin
      valid_235_1 <= _GEN_1774;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_236_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_236_0 <= _GEN_1263;
        end else begin
          valid_236_0 <= _GEN_7692;
        end
      end else begin
        valid_236_0 <= _GEN_1263;
      end
    end else begin
      valid_236_0 <= _GEN_1263;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_236_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_236_1 <= _GEN_1775;
        end else begin
          valid_236_1 <= _GEN_7693;
        end
      end else begin
        valid_236_1 <= _GEN_1775;
      end
    end else begin
      valid_236_1 <= _GEN_1775;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_237_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_237_0 <= _GEN_1264;
        end else begin
          valid_237_0 <= _GEN_7694;
        end
      end else begin
        valid_237_0 <= _GEN_1264;
      end
    end else begin
      valid_237_0 <= _GEN_1264;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_237_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_237_1 <= _GEN_1776;
        end else begin
          valid_237_1 <= _GEN_7695;
        end
      end else begin
        valid_237_1 <= _GEN_1776;
      end
    end else begin
      valid_237_1 <= _GEN_1776;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_238_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_238_0 <= _GEN_1265;
        end else begin
          valid_238_0 <= _GEN_7696;
        end
      end else begin
        valid_238_0 <= _GEN_1265;
      end
    end else begin
      valid_238_0 <= _GEN_1265;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_238_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_238_1 <= _GEN_1777;
        end else begin
          valid_238_1 <= _GEN_7697;
        end
      end else begin
        valid_238_1 <= _GEN_1777;
      end
    end else begin
      valid_238_1 <= _GEN_1777;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_239_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_239_0 <= _GEN_1266;
        end else begin
          valid_239_0 <= _GEN_7698;
        end
      end else begin
        valid_239_0 <= _GEN_1266;
      end
    end else begin
      valid_239_0 <= _GEN_1266;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_239_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_239_1 <= _GEN_1778;
        end else begin
          valid_239_1 <= _GEN_7699;
        end
      end else begin
        valid_239_1 <= _GEN_1778;
      end
    end else begin
      valid_239_1 <= _GEN_1778;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_240_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_240_0 <= _GEN_1267;
        end else begin
          valid_240_0 <= _GEN_7700;
        end
      end else begin
        valid_240_0 <= _GEN_1267;
      end
    end else begin
      valid_240_0 <= _GEN_1267;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_240_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_240_1 <= _GEN_1779;
        end else begin
          valid_240_1 <= _GEN_7701;
        end
      end else begin
        valid_240_1 <= _GEN_1779;
      end
    end else begin
      valid_240_1 <= _GEN_1779;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_241_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_241_0 <= _GEN_1268;
        end else begin
          valid_241_0 <= _GEN_7702;
        end
      end else begin
        valid_241_0 <= _GEN_1268;
      end
    end else begin
      valid_241_0 <= _GEN_1268;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_241_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_241_1 <= _GEN_1780;
        end else begin
          valid_241_1 <= _GEN_7703;
        end
      end else begin
        valid_241_1 <= _GEN_1780;
      end
    end else begin
      valid_241_1 <= _GEN_1780;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_242_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_242_0 <= _GEN_1269;
        end else begin
          valid_242_0 <= _GEN_7704;
        end
      end else begin
        valid_242_0 <= _GEN_1269;
      end
    end else begin
      valid_242_0 <= _GEN_1269;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_242_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_242_1 <= _GEN_1781;
        end else begin
          valid_242_1 <= _GEN_7705;
        end
      end else begin
        valid_242_1 <= _GEN_1781;
      end
    end else begin
      valid_242_1 <= _GEN_1781;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_243_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_243_0 <= _GEN_1270;
        end else begin
          valid_243_0 <= _GEN_7706;
        end
      end else begin
        valid_243_0 <= _GEN_1270;
      end
    end else begin
      valid_243_0 <= _GEN_1270;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_243_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_243_1 <= _GEN_1782;
        end else begin
          valid_243_1 <= _GEN_7707;
        end
      end else begin
        valid_243_1 <= _GEN_1782;
      end
    end else begin
      valid_243_1 <= _GEN_1782;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_244_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_244_0 <= _GEN_1271;
        end else begin
          valid_244_0 <= _GEN_7708;
        end
      end else begin
        valid_244_0 <= _GEN_1271;
      end
    end else begin
      valid_244_0 <= _GEN_1271;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_244_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_244_1 <= _GEN_1783;
        end else begin
          valid_244_1 <= _GEN_7709;
        end
      end else begin
        valid_244_1 <= _GEN_1783;
      end
    end else begin
      valid_244_1 <= _GEN_1783;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_245_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_245_0 <= _GEN_1272;
        end else begin
          valid_245_0 <= _GEN_7710;
        end
      end else begin
        valid_245_0 <= _GEN_1272;
      end
    end else begin
      valid_245_0 <= _GEN_1272;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_245_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_245_1 <= _GEN_1784;
        end else begin
          valid_245_1 <= _GEN_7711;
        end
      end else begin
        valid_245_1 <= _GEN_1784;
      end
    end else begin
      valid_245_1 <= _GEN_1784;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_246_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_246_0 <= _GEN_1273;
        end else begin
          valid_246_0 <= _GEN_7712;
        end
      end else begin
        valid_246_0 <= _GEN_1273;
      end
    end else begin
      valid_246_0 <= _GEN_1273;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_246_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_246_1 <= _GEN_1785;
        end else begin
          valid_246_1 <= _GEN_7713;
        end
      end else begin
        valid_246_1 <= _GEN_1785;
      end
    end else begin
      valid_246_1 <= _GEN_1785;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_247_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_247_0 <= _GEN_1274;
        end else begin
          valid_247_0 <= _GEN_7714;
        end
      end else begin
        valid_247_0 <= _GEN_1274;
      end
    end else begin
      valid_247_0 <= _GEN_1274;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_247_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_247_1 <= _GEN_1786;
        end else begin
          valid_247_1 <= _GEN_7715;
        end
      end else begin
        valid_247_1 <= _GEN_1786;
      end
    end else begin
      valid_247_1 <= _GEN_1786;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_248_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_248_0 <= _GEN_1275;
        end else begin
          valid_248_0 <= _GEN_7716;
        end
      end else begin
        valid_248_0 <= _GEN_1275;
      end
    end else begin
      valid_248_0 <= _GEN_1275;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_248_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_248_1 <= _GEN_1787;
        end else begin
          valid_248_1 <= _GEN_7717;
        end
      end else begin
        valid_248_1 <= _GEN_1787;
      end
    end else begin
      valid_248_1 <= _GEN_1787;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_249_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_249_0 <= _GEN_1276;
        end else begin
          valid_249_0 <= _GEN_7718;
        end
      end else begin
        valid_249_0 <= _GEN_1276;
      end
    end else begin
      valid_249_0 <= _GEN_1276;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_249_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_249_1 <= _GEN_1788;
        end else begin
          valid_249_1 <= _GEN_7719;
        end
      end else begin
        valid_249_1 <= _GEN_1788;
      end
    end else begin
      valid_249_1 <= _GEN_1788;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_250_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_250_0 <= _GEN_1277;
        end else begin
          valid_250_0 <= _GEN_7720;
        end
      end else begin
        valid_250_0 <= _GEN_1277;
      end
    end else begin
      valid_250_0 <= _GEN_1277;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_250_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_250_1 <= _GEN_1789;
        end else begin
          valid_250_1 <= _GEN_7721;
        end
      end else begin
        valid_250_1 <= _GEN_1789;
      end
    end else begin
      valid_250_1 <= _GEN_1789;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_251_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_251_0 <= _GEN_1278;
        end else begin
          valid_251_0 <= _GEN_7722;
        end
      end else begin
        valid_251_0 <= _GEN_1278;
      end
    end else begin
      valid_251_0 <= _GEN_1278;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_251_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_251_1 <= _GEN_1790;
        end else begin
          valid_251_1 <= _GEN_7723;
        end
      end else begin
        valid_251_1 <= _GEN_1790;
      end
    end else begin
      valid_251_1 <= _GEN_1790;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_252_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_252_0 <= _GEN_1279;
        end else begin
          valid_252_0 <= _GEN_7724;
        end
      end else begin
        valid_252_0 <= _GEN_1279;
      end
    end else begin
      valid_252_0 <= _GEN_1279;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_252_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_252_1 <= _GEN_1791;
        end else begin
          valid_252_1 <= _GEN_7725;
        end
      end else begin
        valid_252_1 <= _GEN_1791;
      end
    end else begin
      valid_252_1 <= _GEN_1791;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_253_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_253_0 <= _GEN_1280;
        end else begin
          valid_253_0 <= _GEN_7726;
        end
      end else begin
        valid_253_0 <= _GEN_1280;
      end
    end else begin
      valid_253_0 <= _GEN_1280;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_253_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_253_1 <= _GEN_1792;
        end else begin
          valid_253_1 <= _GEN_7727;
        end
      end else begin
        valid_253_1 <= _GEN_1792;
      end
    end else begin
      valid_253_1 <= _GEN_1792;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_254_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_254_0 <= _GEN_1281;
        end else begin
          valid_254_0 <= _GEN_7728;
        end
      end else begin
        valid_254_0 <= _GEN_1281;
      end
    end else begin
      valid_254_0 <= _GEN_1281;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_254_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_254_1 <= _GEN_1793;
        end else begin
          valid_254_1 <= _GEN_7729;
        end
      end else begin
        valid_254_1 <= _GEN_1793;
      end
    end else begin
      valid_254_1 <= _GEN_1793;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_255_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_255_0 <= _GEN_1282;
        end else begin
          valid_255_0 <= _GEN_7730;
        end
      end else begin
        valid_255_0 <= _GEN_1282;
      end
    end else begin
      valid_255_0 <= _GEN_1282;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_255_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_255_1 <= _GEN_1794;
        end else begin
          valid_255_1 <= _GEN_7731;
        end
      end else begin
        valid_255_1 <= _GEN_1794;
      end
    end else begin
      valid_255_1 <= _GEN_1794;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_256_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_256_0 <= _GEN_1283;
        end else begin
          valid_256_0 <= _GEN_7732;
        end
      end else begin
        valid_256_0 <= _GEN_1283;
      end
    end else begin
      valid_256_0 <= _GEN_1283;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_256_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_256_1 <= _GEN_1795;
        end else begin
          valid_256_1 <= _GEN_7733;
        end
      end else begin
        valid_256_1 <= _GEN_1795;
      end
    end else begin
      valid_256_1 <= _GEN_1795;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_257_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_257_0 <= _GEN_1284;
        end else begin
          valid_257_0 <= _GEN_7734;
        end
      end else begin
        valid_257_0 <= _GEN_1284;
      end
    end else begin
      valid_257_0 <= _GEN_1284;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_257_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_257_1 <= _GEN_1796;
        end else begin
          valid_257_1 <= _GEN_7735;
        end
      end else begin
        valid_257_1 <= _GEN_1796;
      end
    end else begin
      valid_257_1 <= _GEN_1796;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_258_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_258_0 <= _GEN_1285;
        end else begin
          valid_258_0 <= _GEN_7736;
        end
      end else begin
        valid_258_0 <= _GEN_1285;
      end
    end else begin
      valid_258_0 <= _GEN_1285;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_258_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_258_1 <= _GEN_1797;
        end else begin
          valid_258_1 <= _GEN_7737;
        end
      end else begin
        valid_258_1 <= _GEN_1797;
      end
    end else begin
      valid_258_1 <= _GEN_1797;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_259_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_259_0 <= _GEN_1286;
        end else begin
          valid_259_0 <= _GEN_7738;
        end
      end else begin
        valid_259_0 <= _GEN_1286;
      end
    end else begin
      valid_259_0 <= _GEN_1286;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_259_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_259_1 <= _GEN_1798;
        end else begin
          valid_259_1 <= _GEN_7739;
        end
      end else begin
        valid_259_1 <= _GEN_1798;
      end
    end else begin
      valid_259_1 <= _GEN_1798;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_260_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_260_0 <= _GEN_1287;
        end else begin
          valid_260_0 <= _GEN_7740;
        end
      end else begin
        valid_260_0 <= _GEN_1287;
      end
    end else begin
      valid_260_0 <= _GEN_1287;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_260_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_260_1 <= _GEN_1799;
        end else begin
          valid_260_1 <= _GEN_7741;
        end
      end else begin
        valid_260_1 <= _GEN_1799;
      end
    end else begin
      valid_260_1 <= _GEN_1799;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_261_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_261_0 <= _GEN_1288;
        end else begin
          valid_261_0 <= _GEN_7742;
        end
      end else begin
        valid_261_0 <= _GEN_1288;
      end
    end else begin
      valid_261_0 <= _GEN_1288;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_261_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_261_1 <= _GEN_1800;
        end else begin
          valid_261_1 <= _GEN_7743;
        end
      end else begin
        valid_261_1 <= _GEN_1800;
      end
    end else begin
      valid_261_1 <= _GEN_1800;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_262_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_262_0 <= _GEN_1289;
        end else begin
          valid_262_0 <= _GEN_7744;
        end
      end else begin
        valid_262_0 <= _GEN_1289;
      end
    end else begin
      valid_262_0 <= _GEN_1289;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_262_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_262_1 <= _GEN_1801;
        end else begin
          valid_262_1 <= _GEN_7745;
        end
      end else begin
        valid_262_1 <= _GEN_1801;
      end
    end else begin
      valid_262_1 <= _GEN_1801;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_263_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_263_0 <= _GEN_1290;
        end else begin
          valid_263_0 <= _GEN_7746;
        end
      end else begin
        valid_263_0 <= _GEN_1290;
      end
    end else begin
      valid_263_0 <= _GEN_1290;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_263_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_263_1 <= _GEN_1802;
        end else begin
          valid_263_1 <= _GEN_7747;
        end
      end else begin
        valid_263_1 <= _GEN_1802;
      end
    end else begin
      valid_263_1 <= _GEN_1802;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_264_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_264_0 <= _GEN_1291;
        end else begin
          valid_264_0 <= _GEN_7748;
        end
      end else begin
        valid_264_0 <= _GEN_1291;
      end
    end else begin
      valid_264_0 <= _GEN_1291;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_264_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_264_1 <= _GEN_1803;
        end else begin
          valid_264_1 <= _GEN_7749;
        end
      end else begin
        valid_264_1 <= _GEN_1803;
      end
    end else begin
      valid_264_1 <= _GEN_1803;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_265_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_265_0 <= _GEN_1292;
        end else begin
          valid_265_0 <= _GEN_7750;
        end
      end else begin
        valid_265_0 <= _GEN_1292;
      end
    end else begin
      valid_265_0 <= _GEN_1292;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_265_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_265_1 <= _GEN_1804;
        end else begin
          valid_265_1 <= _GEN_7751;
        end
      end else begin
        valid_265_1 <= _GEN_1804;
      end
    end else begin
      valid_265_1 <= _GEN_1804;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_266_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_266_0 <= _GEN_1293;
        end else begin
          valid_266_0 <= _GEN_7752;
        end
      end else begin
        valid_266_0 <= _GEN_1293;
      end
    end else begin
      valid_266_0 <= _GEN_1293;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_266_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_266_1 <= _GEN_1805;
        end else begin
          valid_266_1 <= _GEN_7753;
        end
      end else begin
        valid_266_1 <= _GEN_1805;
      end
    end else begin
      valid_266_1 <= _GEN_1805;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_267_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_267_0 <= _GEN_1294;
        end else begin
          valid_267_0 <= _GEN_7754;
        end
      end else begin
        valid_267_0 <= _GEN_1294;
      end
    end else begin
      valid_267_0 <= _GEN_1294;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_267_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_267_1 <= _GEN_1806;
        end else begin
          valid_267_1 <= _GEN_7755;
        end
      end else begin
        valid_267_1 <= _GEN_1806;
      end
    end else begin
      valid_267_1 <= _GEN_1806;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_268_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_268_0 <= _GEN_1295;
        end else begin
          valid_268_0 <= _GEN_7756;
        end
      end else begin
        valid_268_0 <= _GEN_1295;
      end
    end else begin
      valid_268_0 <= _GEN_1295;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_268_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_268_1 <= _GEN_1807;
        end else begin
          valid_268_1 <= _GEN_7757;
        end
      end else begin
        valid_268_1 <= _GEN_1807;
      end
    end else begin
      valid_268_1 <= _GEN_1807;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_269_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_269_0 <= _GEN_1296;
        end else begin
          valid_269_0 <= _GEN_7758;
        end
      end else begin
        valid_269_0 <= _GEN_1296;
      end
    end else begin
      valid_269_0 <= _GEN_1296;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_269_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_269_1 <= _GEN_1808;
        end else begin
          valid_269_1 <= _GEN_7759;
        end
      end else begin
        valid_269_1 <= _GEN_1808;
      end
    end else begin
      valid_269_1 <= _GEN_1808;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_270_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_270_0 <= _GEN_1297;
        end else begin
          valid_270_0 <= _GEN_7760;
        end
      end else begin
        valid_270_0 <= _GEN_1297;
      end
    end else begin
      valid_270_0 <= _GEN_1297;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_270_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_270_1 <= _GEN_1809;
        end else begin
          valid_270_1 <= _GEN_7761;
        end
      end else begin
        valid_270_1 <= _GEN_1809;
      end
    end else begin
      valid_270_1 <= _GEN_1809;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_271_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_271_0 <= _GEN_1298;
        end else begin
          valid_271_0 <= _GEN_7762;
        end
      end else begin
        valid_271_0 <= _GEN_1298;
      end
    end else begin
      valid_271_0 <= _GEN_1298;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_271_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_271_1 <= _GEN_1810;
        end else begin
          valid_271_1 <= _GEN_7763;
        end
      end else begin
        valid_271_1 <= _GEN_1810;
      end
    end else begin
      valid_271_1 <= _GEN_1810;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_272_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_272_0 <= _GEN_1299;
        end else begin
          valid_272_0 <= _GEN_7764;
        end
      end else begin
        valid_272_0 <= _GEN_1299;
      end
    end else begin
      valid_272_0 <= _GEN_1299;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_272_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_272_1 <= _GEN_1811;
        end else begin
          valid_272_1 <= _GEN_7765;
        end
      end else begin
        valid_272_1 <= _GEN_1811;
      end
    end else begin
      valid_272_1 <= _GEN_1811;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_273_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_273_0 <= _GEN_1300;
        end else begin
          valid_273_0 <= _GEN_7766;
        end
      end else begin
        valid_273_0 <= _GEN_1300;
      end
    end else begin
      valid_273_0 <= _GEN_1300;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_273_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_273_1 <= _GEN_1812;
        end else begin
          valid_273_1 <= _GEN_7767;
        end
      end else begin
        valid_273_1 <= _GEN_1812;
      end
    end else begin
      valid_273_1 <= _GEN_1812;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_274_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_274_0 <= _GEN_1301;
        end else begin
          valid_274_0 <= _GEN_7768;
        end
      end else begin
        valid_274_0 <= _GEN_1301;
      end
    end else begin
      valid_274_0 <= _GEN_1301;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_274_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_274_1 <= _GEN_1813;
        end else begin
          valid_274_1 <= _GEN_7769;
        end
      end else begin
        valid_274_1 <= _GEN_1813;
      end
    end else begin
      valid_274_1 <= _GEN_1813;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_275_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_275_0 <= _GEN_1302;
        end else begin
          valid_275_0 <= _GEN_7770;
        end
      end else begin
        valid_275_0 <= _GEN_1302;
      end
    end else begin
      valid_275_0 <= _GEN_1302;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_275_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_275_1 <= _GEN_1814;
        end else begin
          valid_275_1 <= _GEN_7771;
        end
      end else begin
        valid_275_1 <= _GEN_1814;
      end
    end else begin
      valid_275_1 <= _GEN_1814;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_276_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_276_0 <= _GEN_1303;
        end else begin
          valid_276_0 <= _GEN_7772;
        end
      end else begin
        valid_276_0 <= _GEN_1303;
      end
    end else begin
      valid_276_0 <= _GEN_1303;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_276_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_276_1 <= _GEN_1815;
        end else begin
          valid_276_1 <= _GEN_7773;
        end
      end else begin
        valid_276_1 <= _GEN_1815;
      end
    end else begin
      valid_276_1 <= _GEN_1815;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_277_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_277_0 <= _GEN_1304;
        end else begin
          valid_277_0 <= _GEN_7774;
        end
      end else begin
        valid_277_0 <= _GEN_1304;
      end
    end else begin
      valid_277_0 <= _GEN_1304;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_277_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_277_1 <= _GEN_1816;
        end else begin
          valid_277_1 <= _GEN_7775;
        end
      end else begin
        valid_277_1 <= _GEN_1816;
      end
    end else begin
      valid_277_1 <= _GEN_1816;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_278_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_278_0 <= _GEN_1305;
        end else begin
          valid_278_0 <= _GEN_7776;
        end
      end else begin
        valid_278_0 <= _GEN_1305;
      end
    end else begin
      valid_278_0 <= _GEN_1305;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_278_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_278_1 <= _GEN_1817;
        end else begin
          valid_278_1 <= _GEN_7777;
        end
      end else begin
        valid_278_1 <= _GEN_1817;
      end
    end else begin
      valid_278_1 <= _GEN_1817;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_279_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_279_0 <= _GEN_1306;
        end else begin
          valid_279_0 <= _GEN_7778;
        end
      end else begin
        valid_279_0 <= _GEN_1306;
      end
    end else begin
      valid_279_0 <= _GEN_1306;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_279_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_279_1 <= _GEN_1818;
        end else begin
          valid_279_1 <= _GEN_7779;
        end
      end else begin
        valid_279_1 <= _GEN_1818;
      end
    end else begin
      valid_279_1 <= _GEN_1818;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_280_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_280_0 <= _GEN_1307;
        end else begin
          valid_280_0 <= _GEN_7780;
        end
      end else begin
        valid_280_0 <= _GEN_1307;
      end
    end else begin
      valid_280_0 <= _GEN_1307;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_280_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_280_1 <= _GEN_1819;
        end else begin
          valid_280_1 <= _GEN_7781;
        end
      end else begin
        valid_280_1 <= _GEN_1819;
      end
    end else begin
      valid_280_1 <= _GEN_1819;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_281_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_281_0 <= _GEN_1308;
        end else begin
          valid_281_0 <= _GEN_7782;
        end
      end else begin
        valid_281_0 <= _GEN_1308;
      end
    end else begin
      valid_281_0 <= _GEN_1308;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_281_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_281_1 <= _GEN_1820;
        end else begin
          valid_281_1 <= _GEN_7783;
        end
      end else begin
        valid_281_1 <= _GEN_1820;
      end
    end else begin
      valid_281_1 <= _GEN_1820;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_282_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_282_0 <= _GEN_1309;
        end else begin
          valid_282_0 <= _GEN_7784;
        end
      end else begin
        valid_282_0 <= _GEN_1309;
      end
    end else begin
      valid_282_0 <= _GEN_1309;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_282_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_282_1 <= _GEN_1821;
        end else begin
          valid_282_1 <= _GEN_7785;
        end
      end else begin
        valid_282_1 <= _GEN_1821;
      end
    end else begin
      valid_282_1 <= _GEN_1821;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_283_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_283_0 <= _GEN_1310;
        end else begin
          valid_283_0 <= _GEN_7786;
        end
      end else begin
        valid_283_0 <= _GEN_1310;
      end
    end else begin
      valid_283_0 <= _GEN_1310;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_283_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_283_1 <= _GEN_1822;
        end else begin
          valid_283_1 <= _GEN_7787;
        end
      end else begin
        valid_283_1 <= _GEN_1822;
      end
    end else begin
      valid_283_1 <= _GEN_1822;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_284_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_284_0 <= _GEN_1311;
        end else begin
          valid_284_0 <= _GEN_7788;
        end
      end else begin
        valid_284_0 <= _GEN_1311;
      end
    end else begin
      valid_284_0 <= _GEN_1311;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_284_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_284_1 <= _GEN_1823;
        end else begin
          valid_284_1 <= _GEN_7789;
        end
      end else begin
        valid_284_1 <= _GEN_1823;
      end
    end else begin
      valid_284_1 <= _GEN_1823;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_285_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_285_0 <= _GEN_1312;
        end else begin
          valid_285_0 <= _GEN_7790;
        end
      end else begin
        valid_285_0 <= _GEN_1312;
      end
    end else begin
      valid_285_0 <= _GEN_1312;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_285_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_285_1 <= _GEN_1824;
        end else begin
          valid_285_1 <= _GEN_7791;
        end
      end else begin
        valid_285_1 <= _GEN_1824;
      end
    end else begin
      valid_285_1 <= _GEN_1824;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_286_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_286_0 <= _GEN_1313;
        end else begin
          valid_286_0 <= _GEN_7792;
        end
      end else begin
        valid_286_0 <= _GEN_1313;
      end
    end else begin
      valid_286_0 <= _GEN_1313;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_286_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_286_1 <= _GEN_1825;
        end else begin
          valid_286_1 <= _GEN_7793;
        end
      end else begin
        valid_286_1 <= _GEN_1825;
      end
    end else begin
      valid_286_1 <= _GEN_1825;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_287_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_287_0 <= _GEN_1314;
        end else begin
          valid_287_0 <= _GEN_7794;
        end
      end else begin
        valid_287_0 <= _GEN_1314;
      end
    end else begin
      valid_287_0 <= _GEN_1314;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_287_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_287_1 <= _GEN_1826;
        end else begin
          valid_287_1 <= _GEN_7795;
        end
      end else begin
        valid_287_1 <= _GEN_1826;
      end
    end else begin
      valid_287_1 <= _GEN_1826;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_288_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_288_0 <= _GEN_1315;
        end else begin
          valid_288_0 <= _GEN_7796;
        end
      end else begin
        valid_288_0 <= _GEN_1315;
      end
    end else begin
      valid_288_0 <= _GEN_1315;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_288_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_288_1 <= _GEN_1827;
        end else begin
          valid_288_1 <= _GEN_7797;
        end
      end else begin
        valid_288_1 <= _GEN_1827;
      end
    end else begin
      valid_288_1 <= _GEN_1827;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_289_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_289_0 <= _GEN_1316;
        end else begin
          valid_289_0 <= _GEN_7798;
        end
      end else begin
        valid_289_0 <= _GEN_1316;
      end
    end else begin
      valid_289_0 <= _GEN_1316;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_289_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_289_1 <= _GEN_1828;
        end else begin
          valid_289_1 <= _GEN_7799;
        end
      end else begin
        valid_289_1 <= _GEN_1828;
      end
    end else begin
      valid_289_1 <= _GEN_1828;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_290_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_290_0 <= _GEN_1317;
        end else begin
          valid_290_0 <= _GEN_7800;
        end
      end else begin
        valid_290_0 <= _GEN_1317;
      end
    end else begin
      valid_290_0 <= _GEN_1317;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_290_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_290_1 <= _GEN_1829;
        end else begin
          valid_290_1 <= _GEN_7801;
        end
      end else begin
        valid_290_1 <= _GEN_1829;
      end
    end else begin
      valid_290_1 <= _GEN_1829;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_291_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_291_0 <= _GEN_1318;
        end else begin
          valid_291_0 <= _GEN_7802;
        end
      end else begin
        valid_291_0 <= _GEN_1318;
      end
    end else begin
      valid_291_0 <= _GEN_1318;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_291_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_291_1 <= _GEN_1830;
        end else begin
          valid_291_1 <= _GEN_7803;
        end
      end else begin
        valid_291_1 <= _GEN_1830;
      end
    end else begin
      valid_291_1 <= _GEN_1830;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_292_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_292_0 <= _GEN_1319;
        end else begin
          valid_292_0 <= _GEN_7804;
        end
      end else begin
        valid_292_0 <= _GEN_1319;
      end
    end else begin
      valid_292_0 <= _GEN_1319;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_292_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_292_1 <= _GEN_1831;
        end else begin
          valid_292_1 <= _GEN_7805;
        end
      end else begin
        valid_292_1 <= _GEN_1831;
      end
    end else begin
      valid_292_1 <= _GEN_1831;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_293_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_293_0 <= _GEN_1320;
        end else begin
          valid_293_0 <= _GEN_7806;
        end
      end else begin
        valid_293_0 <= _GEN_1320;
      end
    end else begin
      valid_293_0 <= _GEN_1320;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_293_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_293_1 <= _GEN_1832;
        end else begin
          valid_293_1 <= _GEN_7807;
        end
      end else begin
        valid_293_1 <= _GEN_1832;
      end
    end else begin
      valid_293_1 <= _GEN_1832;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_294_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_294_0 <= _GEN_1321;
        end else begin
          valid_294_0 <= _GEN_7808;
        end
      end else begin
        valid_294_0 <= _GEN_1321;
      end
    end else begin
      valid_294_0 <= _GEN_1321;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_294_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_294_1 <= _GEN_1833;
        end else begin
          valid_294_1 <= _GEN_7809;
        end
      end else begin
        valid_294_1 <= _GEN_1833;
      end
    end else begin
      valid_294_1 <= _GEN_1833;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_295_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_295_0 <= _GEN_1322;
        end else begin
          valid_295_0 <= _GEN_7810;
        end
      end else begin
        valid_295_0 <= _GEN_1322;
      end
    end else begin
      valid_295_0 <= _GEN_1322;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_295_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_295_1 <= _GEN_1834;
        end else begin
          valid_295_1 <= _GEN_7811;
        end
      end else begin
        valid_295_1 <= _GEN_1834;
      end
    end else begin
      valid_295_1 <= _GEN_1834;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_296_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_296_0 <= _GEN_1323;
        end else begin
          valid_296_0 <= _GEN_7812;
        end
      end else begin
        valid_296_0 <= _GEN_1323;
      end
    end else begin
      valid_296_0 <= _GEN_1323;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_296_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_296_1 <= _GEN_1835;
        end else begin
          valid_296_1 <= _GEN_7813;
        end
      end else begin
        valid_296_1 <= _GEN_1835;
      end
    end else begin
      valid_296_1 <= _GEN_1835;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_297_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_297_0 <= _GEN_1324;
        end else begin
          valid_297_0 <= _GEN_7814;
        end
      end else begin
        valid_297_0 <= _GEN_1324;
      end
    end else begin
      valid_297_0 <= _GEN_1324;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_297_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_297_1 <= _GEN_1836;
        end else begin
          valid_297_1 <= _GEN_7815;
        end
      end else begin
        valid_297_1 <= _GEN_1836;
      end
    end else begin
      valid_297_1 <= _GEN_1836;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_298_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_298_0 <= _GEN_1325;
        end else begin
          valid_298_0 <= _GEN_7816;
        end
      end else begin
        valid_298_0 <= _GEN_1325;
      end
    end else begin
      valid_298_0 <= _GEN_1325;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_298_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_298_1 <= _GEN_1837;
        end else begin
          valid_298_1 <= _GEN_7817;
        end
      end else begin
        valid_298_1 <= _GEN_1837;
      end
    end else begin
      valid_298_1 <= _GEN_1837;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_299_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_299_0 <= _GEN_1326;
        end else begin
          valid_299_0 <= _GEN_7818;
        end
      end else begin
        valid_299_0 <= _GEN_1326;
      end
    end else begin
      valid_299_0 <= _GEN_1326;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_299_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_299_1 <= _GEN_1838;
        end else begin
          valid_299_1 <= _GEN_7819;
        end
      end else begin
        valid_299_1 <= _GEN_1838;
      end
    end else begin
      valid_299_1 <= _GEN_1838;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_300_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_300_0 <= _GEN_1327;
        end else begin
          valid_300_0 <= _GEN_7820;
        end
      end else begin
        valid_300_0 <= _GEN_1327;
      end
    end else begin
      valid_300_0 <= _GEN_1327;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_300_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_300_1 <= _GEN_1839;
        end else begin
          valid_300_1 <= _GEN_7821;
        end
      end else begin
        valid_300_1 <= _GEN_1839;
      end
    end else begin
      valid_300_1 <= _GEN_1839;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_301_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_301_0 <= _GEN_1328;
        end else begin
          valid_301_0 <= _GEN_7822;
        end
      end else begin
        valid_301_0 <= _GEN_1328;
      end
    end else begin
      valid_301_0 <= _GEN_1328;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_301_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_301_1 <= _GEN_1840;
        end else begin
          valid_301_1 <= _GEN_7823;
        end
      end else begin
        valid_301_1 <= _GEN_1840;
      end
    end else begin
      valid_301_1 <= _GEN_1840;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_302_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_302_0 <= _GEN_1329;
        end else begin
          valid_302_0 <= _GEN_7824;
        end
      end else begin
        valid_302_0 <= _GEN_1329;
      end
    end else begin
      valid_302_0 <= _GEN_1329;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_302_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_302_1 <= _GEN_1841;
        end else begin
          valid_302_1 <= _GEN_7825;
        end
      end else begin
        valid_302_1 <= _GEN_1841;
      end
    end else begin
      valid_302_1 <= _GEN_1841;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_303_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_303_0 <= _GEN_1330;
        end else begin
          valid_303_0 <= _GEN_7826;
        end
      end else begin
        valid_303_0 <= _GEN_1330;
      end
    end else begin
      valid_303_0 <= _GEN_1330;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_303_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_303_1 <= _GEN_1842;
        end else begin
          valid_303_1 <= _GEN_7827;
        end
      end else begin
        valid_303_1 <= _GEN_1842;
      end
    end else begin
      valid_303_1 <= _GEN_1842;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_304_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_304_0 <= _GEN_1331;
        end else begin
          valid_304_0 <= _GEN_7828;
        end
      end else begin
        valid_304_0 <= _GEN_1331;
      end
    end else begin
      valid_304_0 <= _GEN_1331;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_304_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_304_1 <= _GEN_1843;
        end else begin
          valid_304_1 <= _GEN_7829;
        end
      end else begin
        valid_304_1 <= _GEN_1843;
      end
    end else begin
      valid_304_1 <= _GEN_1843;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_305_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_305_0 <= _GEN_1332;
        end else begin
          valid_305_0 <= _GEN_7830;
        end
      end else begin
        valid_305_0 <= _GEN_1332;
      end
    end else begin
      valid_305_0 <= _GEN_1332;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_305_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_305_1 <= _GEN_1844;
        end else begin
          valid_305_1 <= _GEN_7831;
        end
      end else begin
        valid_305_1 <= _GEN_1844;
      end
    end else begin
      valid_305_1 <= _GEN_1844;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_306_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_306_0 <= _GEN_1333;
        end else begin
          valid_306_0 <= _GEN_7832;
        end
      end else begin
        valid_306_0 <= _GEN_1333;
      end
    end else begin
      valid_306_0 <= _GEN_1333;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_306_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_306_1 <= _GEN_1845;
        end else begin
          valid_306_1 <= _GEN_7833;
        end
      end else begin
        valid_306_1 <= _GEN_1845;
      end
    end else begin
      valid_306_1 <= _GEN_1845;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_307_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_307_0 <= _GEN_1334;
        end else begin
          valid_307_0 <= _GEN_7834;
        end
      end else begin
        valid_307_0 <= _GEN_1334;
      end
    end else begin
      valid_307_0 <= _GEN_1334;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_307_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_307_1 <= _GEN_1846;
        end else begin
          valid_307_1 <= _GEN_7835;
        end
      end else begin
        valid_307_1 <= _GEN_1846;
      end
    end else begin
      valid_307_1 <= _GEN_1846;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_308_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_308_0 <= _GEN_1335;
        end else begin
          valid_308_0 <= _GEN_7836;
        end
      end else begin
        valid_308_0 <= _GEN_1335;
      end
    end else begin
      valid_308_0 <= _GEN_1335;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_308_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_308_1 <= _GEN_1847;
        end else begin
          valid_308_1 <= _GEN_7837;
        end
      end else begin
        valid_308_1 <= _GEN_1847;
      end
    end else begin
      valid_308_1 <= _GEN_1847;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_309_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_309_0 <= _GEN_1336;
        end else begin
          valid_309_0 <= _GEN_7838;
        end
      end else begin
        valid_309_0 <= _GEN_1336;
      end
    end else begin
      valid_309_0 <= _GEN_1336;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_309_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_309_1 <= _GEN_1848;
        end else begin
          valid_309_1 <= _GEN_7839;
        end
      end else begin
        valid_309_1 <= _GEN_1848;
      end
    end else begin
      valid_309_1 <= _GEN_1848;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_310_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_310_0 <= _GEN_1337;
        end else begin
          valid_310_0 <= _GEN_7840;
        end
      end else begin
        valid_310_0 <= _GEN_1337;
      end
    end else begin
      valid_310_0 <= _GEN_1337;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_310_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_310_1 <= _GEN_1849;
        end else begin
          valid_310_1 <= _GEN_7841;
        end
      end else begin
        valid_310_1 <= _GEN_1849;
      end
    end else begin
      valid_310_1 <= _GEN_1849;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_311_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_311_0 <= _GEN_1338;
        end else begin
          valid_311_0 <= _GEN_7842;
        end
      end else begin
        valid_311_0 <= _GEN_1338;
      end
    end else begin
      valid_311_0 <= _GEN_1338;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_311_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_311_1 <= _GEN_1850;
        end else begin
          valid_311_1 <= _GEN_7843;
        end
      end else begin
        valid_311_1 <= _GEN_1850;
      end
    end else begin
      valid_311_1 <= _GEN_1850;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_312_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_312_0 <= _GEN_1339;
        end else begin
          valid_312_0 <= _GEN_7844;
        end
      end else begin
        valid_312_0 <= _GEN_1339;
      end
    end else begin
      valid_312_0 <= _GEN_1339;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_312_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_312_1 <= _GEN_1851;
        end else begin
          valid_312_1 <= _GEN_7845;
        end
      end else begin
        valid_312_1 <= _GEN_1851;
      end
    end else begin
      valid_312_1 <= _GEN_1851;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_313_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_313_0 <= _GEN_1340;
        end else begin
          valid_313_0 <= _GEN_7846;
        end
      end else begin
        valid_313_0 <= _GEN_1340;
      end
    end else begin
      valid_313_0 <= _GEN_1340;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_313_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_313_1 <= _GEN_1852;
        end else begin
          valid_313_1 <= _GEN_7847;
        end
      end else begin
        valid_313_1 <= _GEN_1852;
      end
    end else begin
      valid_313_1 <= _GEN_1852;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_314_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_314_0 <= _GEN_1341;
        end else begin
          valid_314_0 <= _GEN_7848;
        end
      end else begin
        valid_314_0 <= _GEN_1341;
      end
    end else begin
      valid_314_0 <= _GEN_1341;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_314_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_314_1 <= _GEN_1853;
        end else begin
          valid_314_1 <= _GEN_7849;
        end
      end else begin
        valid_314_1 <= _GEN_1853;
      end
    end else begin
      valid_314_1 <= _GEN_1853;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_315_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_315_0 <= _GEN_1342;
        end else begin
          valid_315_0 <= _GEN_7850;
        end
      end else begin
        valid_315_0 <= _GEN_1342;
      end
    end else begin
      valid_315_0 <= _GEN_1342;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_315_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_315_1 <= _GEN_1854;
        end else begin
          valid_315_1 <= _GEN_7851;
        end
      end else begin
        valid_315_1 <= _GEN_1854;
      end
    end else begin
      valid_315_1 <= _GEN_1854;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_316_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_316_0 <= _GEN_1343;
        end else begin
          valid_316_0 <= _GEN_7852;
        end
      end else begin
        valid_316_0 <= _GEN_1343;
      end
    end else begin
      valid_316_0 <= _GEN_1343;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_316_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_316_1 <= _GEN_1855;
        end else begin
          valid_316_1 <= _GEN_7853;
        end
      end else begin
        valid_316_1 <= _GEN_1855;
      end
    end else begin
      valid_316_1 <= _GEN_1855;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_317_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_317_0 <= _GEN_1344;
        end else begin
          valid_317_0 <= _GEN_7854;
        end
      end else begin
        valid_317_0 <= _GEN_1344;
      end
    end else begin
      valid_317_0 <= _GEN_1344;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_317_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_317_1 <= _GEN_1856;
        end else begin
          valid_317_1 <= _GEN_7855;
        end
      end else begin
        valid_317_1 <= _GEN_1856;
      end
    end else begin
      valid_317_1 <= _GEN_1856;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_318_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_318_0 <= _GEN_1345;
        end else begin
          valid_318_0 <= _GEN_7856;
        end
      end else begin
        valid_318_0 <= _GEN_1345;
      end
    end else begin
      valid_318_0 <= _GEN_1345;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_318_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_318_1 <= _GEN_1857;
        end else begin
          valid_318_1 <= _GEN_7857;
        end
      end else begin
        valid_318_1 <= _GEN_1857;
      end
    end else begin
      valid_318_1 <= _GEN_1857;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_319_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_319_0 <= _GEN_1346;
        end else begin
          valid_319_0 <= _GEN_7858;
        end
      end else begin
        valid_319_0 <= _GEN_1346;
      end
    end else begin
      valid_319_0 <= _GEN_1346;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_319_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_319_1 <= _GEN_1858;
        end else begin
          valid_319_1 <= _GEN_7859;
        end
      end else begin
        valid_319_1 <= _GEN_1858;
      end
    end else begin
      valid_319_1 <= _GEN_1858;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_320_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_320_0 <= _GEN_1347;
        end else begin
          valid_320_0 <= _GEN_7860;
        end
      end else begin
        valid_320_0 <= _GEN_1347;
      end
    end else begin
      valid_320_0 <= _GEN_1347;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_320_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_320_1 <= _GEN_1859;
        end else begin
          valid_320_1 <= _GEN_7861;
        end
      end else begin
        valid_320_1 <= _GEN_1859;
      end
    end else begin
      valid_320_1 <= _GEN_1859;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_321_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_321_0 <= _GEN_1348;
        end else begin
          valid_321_0 <= _GEN_7862;
        end
      end else begin
        valid_321_0 <= _GEN_1348;
      end
    end else begin
      valid_321_0 <= _GEN_1348;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_321_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_321_1 <= _GEN_1860;
        end else begin
          valid_321_1 <= _GEN_7863;
        end
      end else begin
        valid_321_1 <= _GEN_1860;
      end
    end else begin
      valid_321_1 <= _GEN_1860;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_322_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_322_0 <= _GEN_1349;
        end else begin
          valid_322_0 <= _GEN_7864;
        end
      end else begin
        valid_322_0 <= _GEN_1349;
      end
    end else begin
      valid_322_0 <= _GEN_1349;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_322_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_322_1 <= _GEN_1861;
        end else begin
          valid_322_1 <= _GEN_7865;
        end
      end else begin
        valid_322_1 <= _GEN_1861;
      end
    end else begin
      valid_322_1 <= _GEN_1861;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_323_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_323_0 <= _GEN_1350;
        end else begin
          valid_323_0 <= _GEN_7866;
        end
      end else begin
        valid_323_0 <= _GEN_1350;
      end
    end else begin
      valid_323_0 <= _GEN_1350;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_323_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_323_1 <= _GEN_1862;
        end else begin
          valid_323_1 <= _GEN_7867;
        end
      end else begin
        valid_323_1 <= _GEN_1862;
      end
    end else begin
      valid_323_1 <= _GEN_1862;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_324_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_324_0 <= _GEN_1351;
        end else begin
          valid_324_0 <= _GEN_7868;
        end
      end else begin
        valid_324_0 <= _GEN_1351;
      end
    end else begin
      valid_324_0 <= _GEN_1351;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_324_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_324_1 <= _GEN_1863;
        end else begin
          valid_324_1 <= _GEN_7869;
        end
      end else begin
        valid_324_1 <= _GEN_1863;
      end
    end else begin
      valid_324_1 <= _GEN_1863;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_325_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_325_0 <= _GEN_1352;
        end else begin
          valid_325_0 <= _GEN_7870;
        end
      end else begin
        valid_325_0 <= _GEN_1352;
      end
    end else begin
      valid_325_0 <= _GEN_1352;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_325_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_325_1 <= _GEN_1864;
        end else begin
          valid_325_1 <= _GEN_7871;
        end
      end else begin
        valid_325_1 <= _GEN_1864;
      end
    end else begin
      valid_325_1 <= _GEN_1864;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_326_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_326_0 <= _GEN_1353;
        end else begin
          valid_326_0 <= _GEN_7872;
        end
      end else begin
        valid_326_0 <= _GEN_1353;
      end
    end else begin
      valid_326_0 <= _GEN_1353;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_326_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_326_1 <= _GEN_1865;
        end else begin
          valid_326_1 <= _GEN_7873;
        end
      end else begin
        valid_326_1 <= _GEN_1865;
      end
    end else begin
      valid_326_1 <= _GEN_1865;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_327_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_327_0 <= _GEN_1354;
        end else begin
          valid_327_0 <= _GEN_7874;
        end
      end else begin
        valid_327_0 <= _GEN_1354;
      end
    end else begin
      valid_327_0 <= _GEN_1354;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_327_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_327_1 <= _GEN_1866;
        end else begin
          valid_327_1 <= _GEN_7875;
        end
      end else begin
        valid_327_1 <= _GEN_1866;
      end
    end else begin
      valid_327_1 <= _GEN_1866;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_328_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_328_0 <= _GEN_1355;
        end else begin
          valid_328_0 <= _GEN_7876;
        end
      end else begin
        valid_328_0 <= _GEN_1355;
      end
    end else begin
      valid_328_0 <= _GEN_1355;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_328_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_328_1 <= _GEN_1867;
        end else begin
          valid_328_1 <= _GEN_7877;
        end
      end else begin
        valid_328_1 <= _GEN_1867;
      end
    end else begin
      valid_328_1 <= _GEN_1867;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_329_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_329_0 <= _GEN_1356;
        end else begin
          valid_329_0 <= _GEN_7878;
        end
      end else begin
        valid_329_0 <= _GEN_1356;
      end
    end else begin
      valid_329_0 <= _GEN_1356;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_329_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_329_1 <= _GEN_1868;
        end else begin
          valid_329_1 <= _GEN_7879;
        end
      end else begin
        valid_329_1 <= _GEN_1868;
      end
    end else begin
      valid_329_1 <= _GEN_1868;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_330_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_330_0 <= _GEN_1357;
        end else begin
          valid_330_0 <= _GEN_7880;
        end
      end else begin
        valid_330_0 <= _GEN_1357;
      end
    end else begin
      valid_330_0 <= _GEN_1357;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_330_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_330_1 <= _GEN_1869;
        end else begin
          valid_330_1 <= _GEN_7881;
        end
      end else begin
        valid_330_1 <= _GEN_1869;
      end
    end else begin
      valid_330_1 <= _GEN_1869;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_331_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_331_0 <= _GEN_1358;
        end else begin
          valid_331_0 <= _GEN_7882;
        end
      end else begin
        valid_331_0 <= _GEN_1358;
      end
    end else begin
      valid_331_0 <= _GEN_1358;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_331_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_331_1 <= _GEN_1870;
        end else begin
          valid_331_1 <= _GEN_7883;
        end
      end else begin
        valid_331_1 <= _GEN_1870;
      end
    end else begin
      valid_331_1 <= _GEN_1870;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_332_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_332_0 <= _GEN_1359;
        end else begin
          valid_332_0 <= _GEN_7884;
        end
      end else begin
        valid_332_0 <= _GEN_1359;
      end
    end else begin
      valid_332_0 <= _GEN_1359;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_332_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_332_1 <= _GEN_1871;
        end else begin
          valid_332_1 <= _GEN_7885;
        end
      end else begin
        valid_332_1 <= _GEN_1871;
      end
    end else begin
      valid_332_1 <= _GEN_1871;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_333_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_333_0 <= _GEN_1360;
        end else begin
          valid_333_0 <= _GEN_7886;
        end
      end else begin
        valid_333_0 <= _GEN_1360;
      end
    end else begin
      valid_333_0 <= _GEN_1360;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_333_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_333_1 <= _GEN_1872;
        end else begin
          valid_333_1 <= _GEN_7887;
        end
      end else begin
        valid_333_1 <= _GEN_1872;
      end
    end else begin
      valid_333_1 <= _GEN_1872;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_334_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_334_0 <= _GEN_1361;
        end else begin
          valid_334_0 <= _GEN_7888;
        end
      end else begin
        valid_334_0 <= _GEN_1361;
      end
    end else begin
      valid_334_0 <= _GEN_1361;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_334_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_334_1 <= _GEN_1873;
        end else begin
          valid_334_1 <= _GEN_7889;
        end
      end else begin
        valid_334_1 <= _GEN_1873;
      end
    end else begin
      valid_334_1 <= _GEN_1873;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_335_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_335_0 <= _GEN_1362;
        end else begin
          valid_335_0 <= _GEN_7890;
        end
      end else begin
        valid_335_0 <= _GEN_1362;
      end
    end else begin
      valid_335_0 <= _GEN_1362;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_335_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_335_1 <= _GEN_1874;
        end else begin
          valid_335_1 <= _GEN_7891;
        end
      end else begin
        valid_335_1 <= _GEN_1874;
      end
    end else begin
      valid_335_1 <= _GEN_1874;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_336_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_336_0 <= _GEN_1363;
        end else begin
          valid_336_0 <= _GEN_7892;
        end
      end else begin
        valid_336_0 <= _GEN_1363;
      end
    end else begin
      valid_336_0 <= _GEN_1363;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_336_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_336_1 <= _GEN_1875;
        end else begin
          valid_336_1 <= _GEN_7893;
        end
      end else begin
        valid_336_1 <= _GEN_1875;
      end
    end else begin
      valid_336_1 <= _GEN_1875;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_337_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_337_0 <= _GEN_1364;
        end else begin
          valid_337_0 <= _GEN_7894;
        end
      end else begin
        valid_337_0 <= _GEN_1364;
      end
    end else begin
      valid_337_0 <= _GEN_1364;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_337_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_337_1 <= _GEN_1876;
        end else begin
          valid_337_1 <= _GEN_7895;
        end
      end else begin
        valid_337_1 <= _GEN_1876;
      end
    end else begin
      valid_337_1 <= _GEN_1876;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_338_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_338_0 <= _GEN_1365;
        end else begin
          valid_338_0 <= _GEN_7896;
        end
      end else begin
        valid_338_0 <= _GEN_1365;
      end
    end else begin
      valid_338_0 <= _GEN_1365;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_338_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_338_1 <= _GEN_1877;
        end else begin
          valid_338_1 <= _GEN_7897;
        end
      end else begin
        valid_338_1 <= _GEN_1877;
      end
    end else begin
      valid_338_1 <= _GEN_1877;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_339_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_339_0 <= _GEN_1366;
        end else begin
          valid_339_0 <= _GEN_7898;
        end
      end else begin
        valid_339_0 <= _GEN_1366;
      end
    end else begin
      valid_339_0 <= _GEN_1366;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_339_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_339_1 <= _GEN_1878;
        end else begin
          valid_339_1 <= _GEN_7899;
        end
      end else begin
        valid_339_1 <= _GEN_1878;
      end
    end else begin
      valid_339_1 <= _GEN_1878;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_340_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_340_0 <= _GEN_1367;
        end else begin
          valid_340_0 <= _GEN_7900;
        end
      end else begin
        valid_340_0 <= _GEN_1367;
      end
    end else begin
      valid_340_0 <= _GEN_1367;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_340_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_340_1 <= _GEN_1879;
        end else begin
          valid_340_1 <= _GEN_7901;
        end
      end else begin
        valid_340_1 <= _GEN_1879;
      end
    end else begin
      valid_340_1 <= _GEN_1879;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_341_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_341_0 <= _GEN_1368;
        end else begin
          valid_341_0 <= _GEN_7902;
        end
      end else begin
        valid_341_0 <= _GEN_1368;
      end
    end else begin
      valid_341_0 <= _GEN_1368;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_341_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_341_1 <= _GEN_1880;
        end else begin
          valid_341_1 <= _GEN_7903;
        end
      end else begin
        valid_341_1 <= _GEN_1880;
      end
    end else begin
      valid_341_1 <= _GEN_1880;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_342_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_342_0 <= _GEN_1369;
        end else begin
          valid_342_0 <= _GEN_7904;
        end
      end else begin
        valid_342_0 <= _GEN_1369;
      end
    end else begin
      valid_342_0 <= _GEN_1369;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_342_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_342_1 <= _GEN_1881;
        end else begin
          valid_342_1 <= _GEN_7905;
        end
      end else begin
        valid_342_1 <= _GEN_1881;
      end
    end else begin
      valid_342_1 <= _GEN_1881;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_343_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_343_0 <= _GEN_1370;
        end else begin
          valid_343_0 <= _GEN_7906;
        end
      end else begin
        valid_343_0 <= _GEN_1370;
      end
    end else begin
      valid_343_0 <= _GEN_1370;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_343_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_343_1 <= _GEN_1882;
        end else begin
          valid_343_1 <= _GEN_7907;
        end
      end else begin
        valid_343_1 <= _GEN_1882;
      end
    end else begin
      valid_343_1 <= _GEN_1882;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_344_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_344_0 <= _GEN_1371;
        end else begin
          valid_344_0 <= _GEN_7908;
        end
      end else begin
        valid_344_0 <= _GEN_1371;
      end
    end else begin
      valid_344_0 <= _GEN_1371;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_344_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_344_1 <= _GEN_1883;
        end else begin
          valid_344_1 <= _GEN_7909;
        end
      end else begin
        valid_344_1 <= _GEN_1883;
      end
    end else begin
      valid_344_1 <= _GEN_1883;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_345_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_345_0 <= _GEN_1372;
        end else begin
          valid_345_0 <= _GEN_7910;
        end
      end else begin
        valid_345_0 <= _GEN_1372;
      end
    end else begin
      valid_345_0 <= _GEN_1372;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_345_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_345_1 <= _GEN_1884;
        end else begin
          valid_345_1 <= _GEN_7911;
        end
      end else begin
        valid_345_1 <= _GEN_1884;
      end
    end else begin
      valid_345_1 <= _GEN_1884;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_346_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_346_0 <= _GEN_1373;
        end else begin
          valid_346_0 <= _GEN_7912;
        end
      end else begin
        valid_346_0 <= _GEN_1373;
      end
    end else begin
      valid_346_0 <= _GEN_1373;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_346_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_346_1 <= _GEN_1885;
        end else begin
          valid_346_1 <= _GEN_7913;
        end
      end else begin
        valid_346_1 <= _GEN_1885;
      end
    end else begin
      valid_346_1 <= _GEN_1885;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_347_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_347_0 <= _GEN_1374;
        end else begin
          valid_347_0 <= _GEN_7914;
        end
      end else begin
        valid_347_0 <= _GEN_1374;
      end
    end else begin
      valid_347_0 <= _GEN_1374;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_347_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_347_1 <= _GEN_1886;
        end else begin
          valid_347_1 <= _GEN_7915;
        end
      end else begin
        valid_347_1 <= _GEN_1886;
      end
    end else begin
      valid_347_1 <= _GEN_1886;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_348_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_348_0 <= _GEN_1375;
        end else begin
          valid_348_0 <= _GEN_7916;
        end
      end else begin
        valid_348_0 <= _GEN_1375;
      end
    end else begin
      valid_348_0 <= _GEN_1375;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_348_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_348_1 <= _GEN_1887;
        end else begin
          valid_348_1 <= _GEN_7917;
        end
      end else begin
        valid_348_1 <= _GEN_1887;
      end
    end else begin
      valid_348_1 <= _GEN_1887;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_349_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_349_0 <= _GEN_1376;
        end else begin
          valid_349_0 <= _GEN_7918;
        end
      end else begin
        valid_349_0 <= _GEN_1376;
      end
    end else begin
      valid_349_0 <= _GEN_1376;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_349_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_349_1 <= _GEN_1888;
        end else begin
          valid_349_1 <= _GEN_7919;
        end
      end else begin
        valid_349_1 <= _GEN_1888;
      end
    end else begin
      valid_349_1 <= _GEN_1888;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_350_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_350_0 <= _GEN_1377;
        end else begin
          valid_350_0 <= _GEN_7920;
        end
      end else begin
        valid_350_0 <= _GEN_1377;
      end
    end else begin
      valid_350_0 <= _GEN_1377;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_350_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_350_1 <= _GEN_1889;
        end else begin
          valid_350_1 <= _GEN_7921;
        end
      end else begin
        valid_350_1 <= _GEN_1889;
      end
    end else begin
      valid_350_1 <= _GEN_1889;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_351_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_351_0 <= _GEN_1378;
        end else begin
          valid_351_0 <= _GEN_7922;
        end
      end else begin
        valid_351_0 <= _GEN_1378;
      end
    end else begin
      valid_351_0 <= _GEN_1378;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_351_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_351_1 <= _GEN_1890;
        end else begin
          valid_351_1 <= _GEN_7923;
        end
      end else begin
        valid_351_1 <= _GEN_1890;
      end
    end else begin
      valid_351_1 <= _GEN_1890;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_352_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_352_0 <= _GEN_1379;
        end else begin
          valid_352_0 <= _GEN_7924;
        end
      end else begin
        valid_352_0 <= _GEN_1379;
      end
    end else begin
      valid_352_0 <= _GEN_1379;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_352_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_352_1 <= _GEN_1891;
        end else begin
          valid_352_1 <= _GEN_7925;
        end
      end else begin
        valid_352_1 <= _GEN_1891;
      end
    end else begin
      valid_352_1 <= _GEN_1891;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_353_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_353_0 <= _GEN_1380;
        end else begin
          valid_353_0 <= _GEN_7926;
        end
      end else begin
        valid_353_0 <= _GEN_1380;
      end
    end else begin
      valid_353_0 <= _GEN_1380;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_353_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_353_1 <= _GEN_1892;
        end else begin
          valid_353_1 <= _GEN_7927;
        end
      end else begin
        valid_353_1 <= _GEN_1892;
      end
    end else begin
      valid_353_1 <= _GEN_1892;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_354_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_354_0 <= _GEN_1381;
        end else begin
          valid_354_0 <= _GEN_7928;
        end
      end else begin
        valid_354_0 <= _GEN_1381;
      end
    end else begin
      valid_354_0 <= _GEN_1381;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_354_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_354_1 <= _GEN_1893;
        end else begin
          valid_354_1 <= _GEN_7929;
        end
      end else begin
        valid_354_1 <= _GEN_1893;
      end
    end else begin
      valid_354_1 <= _GEN_1893;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_355_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_355_0 <= _GEN_1382;
        end else begin
          valid_355_0 <= _GEN_7930;
        end
      end else begin
        valid_355_0 <= _GEN_1382;
      end
    end else begin
      valid_355_0 <= _GEN_1382;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_355_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_355_1 <= _GEN_1894;
        end else begin
          valid_355_1 <= _GEN_7931;
        end
      end else begin
        valid_355_1 <= _GEN_1894;
      end
    end else begin
      valid_355_1 <= _GEN_1894;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_356_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_356_0 <= _GEN_1383;
        end else begin
          valid_356_0 <= _GEN_7932;
        end
      end else begin
        valid_356_0 <= _GEN_1383;
      end
    end else begin
      valid_356_0 <= _GEN_1383;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_356_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_356_1 <= _GEN_1895;
        end else begin
          valid_356_1 <= _GEN_7933;
        end
      end else begin
        valid_356_1 <= _GEN_1895;
      end
    end else begin
      valid_356_1 <= _GEN_1895;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_357_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_357_0 <= _GEN_1384;
        end else begin
          valid_357_0 <= _GEN_7934;
        end
      end else begin
        valid_357_0 <= _GEN_1384;
      end
    end else begin
      valid_357_0 <= _GEN_1384;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_357_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_357_1 <= _GEN_1896;
        end else begin
          valid_357_1 <= _GEN_7935;
        end
      end else begin
        valid_357_1 <= _GEN_1896;
      end
    end else begin
      valid_357_1 <= _GEN_1896;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_358_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_358_0 <= _GEN_1385;
        end else begin
          valid_358_0 <= _GEN_7936;
        end
      end else begin
        valid_358_0 <= _GEN_1385;
      end
    end else begin
      valid_358_0 <= _GEN_1385;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_358_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_358_1 <= _GEN_1897;
        end else begin
          valid_358_1 <= _GEN_7937;
        end
      end else begin
        valid_358_1 <= _GEN_1897;
      end
    end else begin
      valid_358_1 <= _GEN_1897;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_359_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_359_0 <= _GEN_1386;
        end else begin
          valid_359_0 <= _GEN_7938;
        end
      end else begin
        valid_359_0 <= _GEN_1386;
      end
    end else begin
      valid_359_0 <= _GEN_1386;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_359_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_359_1 <= _GEN_1898;
        end else begin
          valid_359_1 <= _GEN_7939;
        end
      end else begin
        valid_359_1 <= _GEN_1898;
      end
    end else begin
      valid_359_1 <= _GEN_1898;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_360_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_360_0 <= _GEN_1387;
        end else begin
          valid_360_0 <= _GEN_7940;
        end
      end else begin
        valid_360_0 <= _GEN_1387;
      end
    end else begin
      valid_360_0 <= _GEN_1387;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_360_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_360_1 <= _GEN_1899;
        end else begin
          valid_360_1 <= _GEN_7941;
        end
      end else begin
        valid_360_1 <= _GEN_1899;
      end
    end else begin
      valid_360_1 <= _GEN_1899;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_361_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_361_0 <= _GEN_1388;
        end else begin
          valid_361_0 <= _GEN_7942;
        end
      end else begin
        valid_361_0 <= _GEN_1388;
      end
    end else begin
      valid_361_0 <= _GEN_1388;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_361_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_361_1 <= _GEN_1900;
        end else begin
          valid_361_1 <= _GEN_7943;
        end
      end else begin
        valid_361_1 <= _GEN_1900;
      end
    end else begin
      valid_361_1 <= _GEN_1900;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_362_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_362_0 <= _GEN_1389;
        end else begin
          valid_362_0 <= _GEN_7944;
        end
      end else begin
        valid_362_0 <= _GEN_1389;
      end
    end else begin
      valid_362_0 <= _GEN_1389;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_362_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_362_1 <= _GEN_1901;
        end else begin
          valid_362_1 <= _GEN_7945;
        end
      end else begin
        valid_362_1 <= _GEN_1901;
      end
    end else begin
      valid_362_1 <= _GEN_1901;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_363_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_363_0 <= _GEN_1390;
        end else begin
          valid_363_0 <= _GEN_7946;
        end
      end else begin
        valid_363_0 <= _GEN_1390;
      end
    end else begin
      valid_363_0 <= _GEN_1390;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_363_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_363_1 <= _GEN_1902;
        end else begin
          valid_363_1 <= _GEN_7947;
        end
      end else begin
        valid_363_1 <= _GEN_1902;
      end
    end else begin
      valid_363_1 <= _GEN_1902;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_364_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_364_0 <= _GEN_1391;
        end else begin
          valid_364_0 <= _GEN_7948;
        end
      end else begin
        valid_364_0 <= _GEN_1391;
      end
    end else begin
      valid_364_0 <= _GEN_1391;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_364_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_364_1 <= _GEN_1903;
        end else begin
          valid_364_1 <= _GEN_7949;
        end
      end else begin
        valid_364_1 <= _GEN_1903;
      end
    end else begin
      valid_364_1 <= _GEN_1903;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_365_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_365_0 <= _GEN_1392;
        end else begin
          valid_365_0 <= _GEN_7950;
        end
      end else begin
        valid_365_0 <= _GEN_1392;
      end
    end else begin
      valid_365_0 <= _GEN_1392;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_365_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_365_1 <= _GEN_1904;
        end else begin
          valid_365_1 <= _GEN_7951;
        end
      end else begin
        valid_365_1 <= _GEN_1904;
      end
    end else begin
      valid_365_1 <= _GEN_1904;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_366_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_366_0 <= _GEN_1393;
        end else begin
          valid_366_0 <= _GEN_7952;
        end
      end else begin
        valid_366_0 <= _GEN_1393;
      end
    end else begin
      valid_366_0 <= _GEN_1393;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_366_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_366_1 <= _GEN_1905;
        end else begin
          valid_366_1 <= _GEN_7953;
        end
      end else begin
        valid_366_1 <= _GEN_1905;
      end
    end else begin
      valid_366_1 <= _GEN_1905;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_367_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_367_0 <= _GEN_1394;
        end else begin
          valid_367_0 <= _GEN_7954;
        end
      end else begin
        valid_367_0 <= _GEN_1394;
      end
    end else begin
      valid_367_0 <= _GEN_1394;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_367_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_367_1 <= _GEN_1906;
        end else begin
          valid_367_1 <= _GEN_7955;
        end
      end else begin
        valid_367_1 <= _GEN_1906;
      end
    end else begin
      valid_367_1 <= _GEN_1906;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_368_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_368_0 <= _GEN_1395;
        end else begin
          valid_368_0 <= _GEN_7956;
        end
      end else begin
        valid_368_0 <= _GEN_1395;
      end
    end else begin
      valid_368_0 <= _GEN_1395;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_368_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_368_1 <= _GEN_1907;
        end else begin
          valid_368_1 <= _GEN_7957;
        end
      end else begin
        valid_368_1 <= _GEN_1907;
      end
    end else begin
      valid_368_1 <= _GEN_1907;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_369_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_369_0 <= _GEN_1396;
        end else begin
          valid_369_0 <= _GEN_7958;
        end
      end else begin
        valid_369_0 <= _GEN_1396;
      end
    end else begin
      valid_369_0 <= _GEN_1396;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_369_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_369_1 <= _GEN_1908;
        end else begin
          valid_369_1 <= _GEN_7959;
        end
      end else begin
        valid_369_1 <= _GEN_1908;
      end
    end else begin
      valid_369_1 <= _GEN_1908;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_370_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_370_0 <= _GEN_1397;
        end else begin
          valid_370_0 <= _GEN_7960;
        end
      end else begin
        valid_370_0 <= _GEN_1397;
      end
    end else begin
      valid_370_0 <= _GEN_1397;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_370_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_370_1 <= _GEN_1909;
        end else begin
          valid_370_1 <= _GEN_7961;
        end
      end else begin
        valid_370_1 <= _GEN_1909;
      end
    end else begin
      valid_370_1 <= _GEN_1909;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_371_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_371_0 <= _GEN_1398;
        end else begin
          valid_371_0 <= _GEN_7962;
        end
      end else begin
        valid_371_0 <= _GEN_1398;
      end
    end else begin
      valid_371_0 <= _GEN_1398;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_371_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_371_1 <= _GEN_1910;
        end else begin
          valid_371_1 <= _GEN_7963;
        end
      end else begin
        valid_371_1 <= _GEN_1910;
      end
    end else begin
      valid_371_1 <= _GEN_1910;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_372_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_372_0 <= _GEN_1399;
        end else begin
          valid_372_0 <= _GEN_7964;
        end
      end else begin
        valid_372_0 <= _GEN_1399;
      end
    end else begin
      valid_372_0 <= _GEN_1399;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_372_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_372_1 <= _GEN_1911;
        end else begin
          valid_372_1 <= _GEN_7965;
        end
      end else begin
        valid_372_1 <= _GEN_1911;
      end
    end else begin
      valid_372_1 <= _GEN_1911;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_373_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_373_0 <= _GEN_1400;
        end else begin
          valid_373_0 <= _GEN_7966;
        end
      end else begin
        valid_373_0 <= _GEN_1400;
      end
    end else begin
      valid_373_0 <= _GEN_1400;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_373_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_373_1 <= _GEN_1912;
        end else begin
          valid_373_1 <= _GEN_7967;
        end
      end else begin
        valid_373_1 <= _GEN_1912;
      end
    end else begin
      valid_373_1 <= _GEN_1912;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_374_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_374_0 <= _GEN_1401;
        end else begin
          valid_374_0 <= _GEN_7968;
        end
      end else begin
        valid_374_0 <= _GEN_1401;
      end
    end else begin
      valid_374_0 <= _GEN_1401;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_374_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_374_1 <= _GEN_1913;
        end else begin
          valid_374_1 <= _GEN_7969;
        end
      end else begin
        valid_374_1 <= _GEN_1913;
      end
    end else begin
      valid_374_1 <= _GEN_1913;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_375_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_375_0 <= _GEN_1402;
        end else begin
          valid_375_0 <= _GEN_7970;
        end
      end else begin
        valid_375_0 <= _GEN_1402;
      end
    end else begin
      valid_375_0 <= _GEN_1402;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_375_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_375_1 <= _GEN_1914;
        end else begin
          valid_375_1 <= _GEN_7971;
        end
      end else begin
        valid_375_1 <= _GEN_1914;
      end
    end else begin
      valid_375_1 <= _GEN_1914;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_376_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_376_0 <= _GEN_1403;
        end else begin
          valid_376_0 <= _GEN_7972;
        end
      end else begin
        valid_376_0 <= _GEN_1403;
      end
    end else begin
      valid_376_0 <= _GEN_1403;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_376_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_376_1 <= _GEN_1915;
        end else begin
          valid_376_1 <= _GEN_7973;
        end
      end else begin
        valid_376_1 <= _GEN_1915;
      end
    end else begin
      valid_376_1 <= _GEN_1915;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_377_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_377_0 <= _GEN_1404;
        end else begin
          valid_377_0 <= _GEN_7974;
        end
      end else begin
        valid_377_0 <= _GEN_1404;
      end
    end else begin
      valid_377_0 <= _GEN_1404;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_377_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_377_1 <= _GEN_1916;
        end else begin
          valid_377_1 <= _GEN_7975;
        end
      end else begin
        valid_377_1 <= _GEN_1916;
      end
    end else begin
      valid_377_1 <= _GEN_1916;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_378_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_378_0 <= _GEN_1405;
        end else begin
          valid_378_0 <= _GEN_7976;
        end
      end else begin
        valid_378_0 <= _GEN_1405;
      end
    end else begin
      valid_378_0 <= _GEN_1405;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_378_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_378_1 <= _GEN_1917;
        end else begin
          valid_378_1 <= _GEN_7977;
        end
      end else begin
        valid_378_1 <= _GEN_1917;
      end
    end else begin
      valid_378_1 <= _GEN_1917;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_379_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_379_0 <= _GEN_1406;
        end else begin
          valid_379_0 <= _GEN_7978;
        end
      end else begin
        valid_379_0 <= _GEN_1406;
      end
    end else begin
      valid_379_0 <= _GEN_1406;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_379_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_379_1 <= _GEN_1918;
        end else begin
          valid_379_1 <= _GEN_7979;
        end
      end else begin
        valid_379_1 <= _GEN_1918;
      end
    end else begin
      valid_379_1 <= _GEN_1918;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_380_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_380_0 <= _GEN_1407;
        end else begin
          valid_380_0 <= _GEN_7980;
        end
      end else begin
        valid_380_0 <= _GEN_1407;
      end
    end else begin
      valid_380_0 <= _GEN_1407;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_380_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_380_1 <= _GEN_1919;
        end else begin
          valid_380_1 <= _GEN_7981;
        end
      end else begin
        valid_380_1 <= _GEN_1919;
      end
    end else begin
      valid_380_1 <= _GEN_1919;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_381_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_381_0 <= _GEN_1408;
        end else begin
          valid_381_0 <= _GEN_7982;
        end
      end else begin
        valid_381_0 <= _GEN_1408;
      end
    end else begin
      valid_381_0 <= _GEN_1408;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_381_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_381_1 <= _GEN_1920;
        end else begin
          valid_381_1 <= _GEN_7983;
        end
      end else begin
        valid_381_1 <= _GEN_1920;
      end
    end else begin
      valid_381_1 <= _GEN_1920;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_382_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_382_0 <= _GEN_1409;
        end else begin
          valid_382_0 <= _GEN_7984;
        end
      end else begin
        valid_382_0 <= _GEN_1409;
      end
    end else begin
      valid_382_0 <= _GEN_1409;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_382_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_382_1 <= _GEN_1921;
        end else begin
          valid_382_1 <= _GEN_7985;
        end
      end else begin
        valid_382_1 <= _GEN_1921;
      end
    end else begin
      valid_382_1 <= _GEN_1921;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_383_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_383_0 <= _GEN_1410;
        end else begin
          valid_383_0 <= _GEN_7986;
        end
      end else begin
        valid_383_0 <= _GEN_1410;
      end
    end else begin
      valid_383_0 <= _GEN_1410;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_383_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_383_1 <= _GEN_1922;
        end else begin
          valid_383_1 <= _GEN_7987;
        end
      end else begin
        valid_383_1 <= _GEN_1922;
      end
    end else begin
      valid_383_1 <= _GEN_1922;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_384_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_384_0 <= _GEN_1411;
        end else begin
          valid_384_0 <= _GEN_7988;
        end
      end else begin
        valid_384_0 <= _GEN_1411;
      end
    end else begin
      valid_384_0 <= _GEN_1411;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_384_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_384_1 <= _GEN_1923;
        end else begin
          valid_384_1 <= _GEN_7989;
        end
      end else begin
        valid_384_1 <= _GEN_1923;
      end
    end else begin
      valid_384_1 <= _GEN_1923;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_385_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_385_0 <= _GEN_1412;
        end else begin
          valid_385_0 <= _GEN_7990;
        end
      end else begin
        valid_385_0 <= _GEN_1412;
      end
    end else begin
      valid_385_0 <= _GEN_1412;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_385_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_385_1 <= _GEN_1924;
        end else begin
          valid_385_1 <= _GEN_7991;
        end
      end else begin
        valid_385_1 <= _GEN_1924;
      end
    end else begin
      valid_385_1 <= _GEN_1924;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_386_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_386_0 <= _GEN_1413;
        end else begin
          valid_386_0 <= _GEN_7992;
        end
      end else begin
        valid_386_0 <= _GEN_1413;
      end
    end else begin
      valid_386_0 <= _GEN_1413;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_386_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_386_1 <= _GEN_1925;
        end else begin
          valid_386_1 <= _GEN_7993;
        end
      end else begin
        valid_386_1 <= _GEN_1925;
      end
    end else begin
      valid_386_1 <= _GEN_1925;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_387_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_387_0 <= _GEN_1414;
        end else begin
          valid_387_0 <= _GEN_7994;
        end
      end else begin
        valid_387_0 <= _GEN_1414;
      end
    end else begin
      valid_387_0 <= _GEN_1414;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_387_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_387_1 <= _GEN_1926;
        end else begin
          valid_387_1 <= _GEN_7995;
        end
      end else begin
        valid_387_1 <= _GEN_1926;
      end
    end else begin
      valid_387_1 <= _GEN_1926;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_388_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_388_0 <= _GEN_1415;
        end else begin
          valid_388_0 <= _GEN_7996;
        end
      end else begin
        valid_388_0 <= _GEN_1415;
      end
    end else begin
      valid_388_0 <= _GEN_1415;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_388_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_388_1 <= _GEN_1927;
        end else begin
          valid_388_1 <= _GEN_7997;
        end
      end else begin
        valid_388_1 <= _GEN_1927;
      end
    end else begin
      valid_388_1 <= _GEN_1927;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_389_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_389_0 <= _GEN_1416;
        end else begin
          valid_389_0 <= _GEN_7998;
        end
      end else begin
        valid_389_0 <= _GEN_1416;
      end
    end else begin
      valid_389_0 <= _GEN_1416;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_389_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_389_1 <= _GEN_1928;
        end else begin
          valid_389_1 <= _GEN_7999;
        end
      end else begin
        valid_389_1 <= _GEN_1928;
      end
    end else begin
      valid_389_1 <= _GEN_1928;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_390_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_390_0 <= _GEN_1417;
        end else begin
          valid_390_0 <= _GEN_8000;
        end
      end else begin
        valid_390_0 <= _GEN_1417;
      end
    end else begin
      valid_390_0 <= _GEN_1417;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_390_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_390_1 <= _GEN_1929;
        end else begin
          valid_390_1 <= _GEN_8001;
        end
      end else begin
        valid_390_1 <= _GEN_1929;
      end
    end else begin
      valid_390_1 <= _GEN_1929;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_391_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_391_0 <= _GEN_1418;
        end else begin
          valid_391_0 <= _GEN_8002;
        end
      end else begin
        valid_391_0 <= _GEN_1418;
      end
    end else begin
      valid_391_0 <= _GEN_1418;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_391_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_391_1 <= _GEN_1930;
        end else begin
          valid_391_1 <= _GEN_8003;
        end
      end else begin
        valid_391_1 <= _GEN_1930;
      end
    end else begin
      valid_391_1 <= _GEN_1930;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_392_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_392_0 <= _GEN_1419;
        end else begin
          valid_392_0 <= _GEN_8004;
        end
      end else begin
        valid_392_0 <= _GEN_1419;
      end
    end else begin
      valid_392_0 <= _GEN_1419;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_392_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_392_1 <= _GEN_1931;
        end else begin
          valid_392_1 <= _GEN_8005;
        end
      end else begin
        valid_392_1 <= _GEN_1931;
      end
    end else begin
      valid_392_1 <= _GEN_1931;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_393_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_393_0 <= _GEN_1420;
        end else begin
          valid_393_0 <= _GEN_8006;
        end
      end else begin
        valid_393_0 <= _GEN_1420;
      end
    end else begin
      valid_393_0 <= _GEN_1420;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_393_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_393_1 <= _GEN_1932;
        end else begin
          valid_393_1 <= _GEN_8007;
        end
      end else begin
        valid_393_1 <= _GEN_1932;
      end
    end else begin
      valid_393_1 <= _GEN_1932;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_394_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_394_0 <= _GEN_1421;
        end else begin
          valid_394_0 <= _GEN_8008;
        end
      end else begin
        valid_394_0 <= _GEN_1421;
      end
    end else begin
      valid_394_0 <= _GEN_1421;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_394_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_394_1 <= _GEN_1933;
        end else begin
          valid_394_1 <= _GEN_8009;
        end
      end else begin
        valid_394_1 <= _GEN_1933;
      end
    end else begin
      valid_394_1 <= _GEN_1933;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_395_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_395_0 <= _GEN_1422;
        end else begin
          valid_395_0 <= _GEN_8010;
        end
      end else begin
        valid_395_0 <= _GEN_1422;
      end
    end else begin
      valid_395_0 <= _GEN_1422;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_395_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_395_1 <= _GEN_1934;
        end else begin
          valid_395_1 <= _GEN_8011;
        end
      end else begin
        valid_395_1 <= _GEN_1934;
      end
    end else begin
      valid_395_1 <= _GEN_1934;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_396_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_396_0 <= _GEN_1423;
        end else begin
          valid_396_0 <= _GEN_8012;
        end
      end else begin
        valid_396_0 <= _GEN_1423;
      end
    end else begin
      valid_396_0 <= _GEN_1423;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_396_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_396_1 <= _GEN_1935;
        end else begin
          valid_396_1 <= _GEN_8013;
        end
      end else begin
        valid_396_1 <= _GEN_1935;
      end
    end else begin
      valid_396_1 <= _GEN_1935;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_397_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_397_0 <= _GEN_1424;
        end else begin
          valid_397_0 <= _GEN_8014;
        end
      end else begin
        valid_397_0 <= _GEN_1424;
      end
    end else begin
      valid_397_0 <= _GEN_1424;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_397_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_397_1 <= _GEN_1936;
        end else begin
          valid_397_1 <= _GEN_8015;
        end
      end else begin
        valid_397_1 <= _GEN_1936;
      end
    end else begin
      valid_397_1 <= _GEN_1936;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_398_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_398_0 <= _GEN_1425;
        end else begin
          valid_398_0 <= _GEN_8016;
        end
      end else begin
        valid_398_0 <= _GEN_1425;
      end
    end else begin
      valid_398_0 <= _GEN_1425;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_398_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_398_1 <= _GEN_1937;
        end else begin
          valid_398_1 <= _GEN_8017;
        end
      end else begin
        valid_398_1 <= _GEN_1937;
      end
    end else begin
      valid_398_1 <= _GEN_1937;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_399_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_399_0 <= _GEN_1426;
        end else begin
          valid_399_0 <= _GEN_8018;
        end
      end else begin
        valid_399_0 <= _GEN_1426;
      end
    end else begin
      valid_399_0 <= _GEN_1426;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_399_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_399_1 <= _GEN_1938;
        end else begin
          valid_399_1 <= _GEN_8019;
        end
      end else begin
        valid_399_1 <= _GEN_1938;
      end
    end else begin
      valid_399_1 <= _GEN_1938;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_400_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_400_0 <= _GEN_1427;
        end else begin
          valid_400_0 <= _GEN_8020;
        end
      end else begin
        valid_400_0 <= _GEN_1427;
      end
    end else begin
      valid_400_0 <= _GEN_1427;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_400_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_400_1 <= _GEN_1939;
        end else begin
          valid_400_1 <= _GEN_8021;
        end
      end else begin
        valid_400_1 <= _GEN_1939;
      end
    end else begin
      valid_400_1 <= _GEN_1939;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_401_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_401_0 <= _GEN_1428;
        end else begin
          valid_401_0 <= _GEN_8022;
        end
      end else begin
        valid_401_0 <= _GEN_1428;
      end
    end else begin
      valid_401_0 <= _GEN_1428;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_401_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_401_1 <= _GEN_1940;
        end else begin
          valid_401_1 <= _GEN_8023;
        end
      end else begin
        valid_401_1 <= _GEN_1940;
      end
    end else begin
      valid_401_1 <= _GEN_1940;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_402_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_402_0 <= _GEN_1429;
        end else begin
          valid_402_0 <= _GEN_8024;
        end
      end else begin
        valid_402_0 <= _GEN_1429;
      end
    end else begin
      valid_402_0 <= _GEN_1429;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_402_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_402_1 <= _GEN_1941;
        end else begin
          valid_402_1 <= _GEN_8025;
        end
      end else begin
        valid_402_1 <= _GEN_1941;
      end
    end else begin
      valid_402_1 <= _GEN_1941;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_403_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_403_0 <= _GEN_1430;
        end else begin
          valid_403_0 <= _GEN_8026;
        end
      end else begin
        valid_403_0 <= _GEN_1430;
      end
    end else begin
      valid_403_0 <= _GEN_1430;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_403_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_403_1 <= _GEN_1942;
        end else begin
          valid_403_1 <= _GEN_8027;
        end
      end else begin
        valid_403_1 <= _GEN_1942;
      end
    end else begin
      valid_403_1 <= _GEN_1942;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_404_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_404_0 <= _GEN_1431;
        end else begin
          valid_404_0 <= _GEN_8028;
        end
      end else begin
        valid_404_0 <= _GEN_1431;
      end
    end else begin
      valid_404_0 <= _GEN_1431;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_404_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_404_1 <= _GEN_1943;
        end else begin
          valid_404_1 <= _GEN_8029;
        end
      end else begin
        valid_404_1 <= _GEN_1943;
      end
    end else begin
      valid_404_1 <= _GEN_1943;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_405_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_405_0 <= _GEN_1432;
        end else begin
          valid_405_0 <= _GEN_8030;
        end
      end else begin
        valid_405_0 <= _GEN_1432;
      end
    end else begin
      valid_405_0 <= _GEN_1432;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_405_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_405_1 <= _GEN_1944;
        end else begin
          valid_405_1 <= _GEN_8031;
        end
      end else begin
        valid_405_1 <= _GEN_1944;
      end
    end else begin
      valid_405_1 <= _GEN_1944;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_406_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_406_0 <= _GEN_1433;
        end else begin
          valid_406_0 <= _GEN_8032;
        end
      end else begin
        valid_406_0 <= _GEN_1433;
      end
    end else begin
      valid_406_0 <= _GEN_1433;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_406_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_406_1 <= _GEN_1945;
        end else begin
          valid_406_1 <= _GEN_8033;
        end
      end else begin
        valid_406_1 <= _GEN_1945;
      end
    end else begin
      valid_406_1 <= _GEN_1945;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_407_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_407_0 <= _GEN_1434;
        end else begin
          valid_407_0 <= _GEN_8034;
        end
      end else begin
        valid_407_0 <= _GEN_1434;
      end
    end else begin
      valid_407_0 <= _GEN_1434;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_407_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_407_1 <= _GEN_1946;
        end else begin
          valid_407_1 <= _GEN_8035;
        end
      end else begin
        valid_407_1 <= _GEN_1946;
      end
    end else begin
      valid_407_1 <= _GEN_1946;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_408_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_408_0 <= _GEN_1435;
        end else begin
          valid_408_0 <= _GEN_8036;
        end
      end else begin
        valid_408_0 <= _GEN_1435;
      end
    end else begin
      valid_408_0 <= _GEN_1435;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_408_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_408_1 <= _GEN_1947;
        end else begin
          valid_408_1 <= _GEN_8037;
        end
      end else begin
        valid_408_1 <= _GEN_1947;
      end
    end else begin
      valid_408_1 <= _GEN_1947;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_409_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_409_0 <= _GEN_1436;
        end else begin
          valid_409_0 <= _GEN_8038;
        end
      end else begin
        valid_409_0 <= _GEN_1436;
      end
    end else begin
      valid_409_0 <= _GEN_1436;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_409_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_409_1 <= _GEN_1948;
        end else begin
          valid_409_1 <= _GEN_8039;
        end
      end else begin
        valid_409_1 <= _GEN_1948;
      end
    end else begin
      valid_409_1 <= _GEN_1948;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_410_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_410_0 <= _GEN_1437;
        end else begin
          valid_410_0 <= _GEN_8040;
        end
      end else begin
        valid_410_0 <= _GEN_1437;
      end
    end else begin
      valid_410_0 <= _GEN_1437;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_410_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_410_1 <= _GEN_1949;
        end else begin
          valid_410_1 <= _GEN_8041;
        end
      end else begin
        valid_410_1 <= _GEN_1949;
      end
    end else begin
      valid_410_1 <= _GEN_1949;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_411_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_411_0 <= _GEN_1438;
        end else begin
          valid_411_0 <= _GEN_8042;
        end
      end else begin
        valid_411_0 <= _GEN_1438;
      end
    end else begin
      valid_411_0 <= _GEN_1438;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_411_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_411_1 <= _GEN_1950;
        end else begin
          valid_411_1 <= _GEN_8043;
        end
      end else begin
        valid_411_1 <= _GEN_1950;
      end
    end else begin
      valid_411_1 <= _GEN_1950;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_412_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_412_0 <= _GEN_1439;
        end else begin
          valid_412_0 <= _GEN_8044;
        end
      end else begin
        valid_412_0 <= _GEN_1439;
      end
    end else begin
      valid_412_0 <= _GEN_1439;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_412_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_412_1 <= _GEN_1951;
        end else begin
          valid_412_1 <= _GEN_8045;
        end
      end else begin
        valid_412_1 <= _GEN_1951;
      end
    end else begin
      valid_412_1 <= _GEN_1951;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_413_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_413_0 <= _GEN_1440;
        end else begin
          valid_413_0 <= _GEN_8046;
        end
      end else begin
        valid_413_0 <= _GEN_1440;
      end
    end else begin
      valid_413_0 <= _GEN_1440;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_413_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_413_1 <= _GEN_1952;
        end else begin
          valid_413_1 <= _GEN_8047;
        end
      end else begin
        valid_413_1 <= _GEN_1952;
      end
    end else begin
      valid_413_1 <= _GEN_1952;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_414_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_414_0 <= _GEN_1441;
        end else begin
          valid_414_0 <= _GEN_8048;
        end
      end else begin
        valid_414_0 <= _GEN_1441;
      end
    end else begin
      valid_414_0 <= _GEN_1441;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_414_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_414_1 <= _GEN_1953;
        end else begin
          valid_414_1 <= _GEN_8049;
        end
      end else begin
        valid_414_1 <= _GEN_1953;
      end
    end else begin
      valid_414_1 <= _GEN_1953;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_415_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_415_0 <= _GEN_1442;
        end else begin
          valid_415_0 <= _GEN_8050;
        end
      end else begin
        valid_415_0 <= _GEN_1442;
      end
    end else begin
      valid_415_0 <= _GEN_1442;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_415_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_415_1 <= _GEN_1954;
        end else begin
          valid_415_1 <= _GEN_8051;
        end
      end else begin
        valid_415_1 <= _GEN_1954;
      end
    end else begin
      valid_415_1 <= _GEN_1954;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_416_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_416_0 <= _GEN_1443;
        end else begin
          valid_416_0 <= _GEN_8052;
        end
      end else begin
        valid_416_0 <= _GEN_1443;
      end
    end else begin
      valid_416_0 <= _GEN_1443;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_416_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_416_1 <= _GEN_1955;
        end else begin
          valid_416_1 <= _GEN_8053;
        end
      end else begin
        valid_416_1 <= _GEN_1955;
      end
    end else begin
      valid_416_1 <= _GEN_1955;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_417_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_417_0 <= _GEN_1444;
        end else begin
          valid_417_0 <= _GEN_8054;
        end
      end else begin
        valid_417_0 <= _GEN_1444;
      end
    end else begin
      valid_417_0 <= _GEN_1444;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_417_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_417_1 <= _GEN_1956;
        end else begin
          valid_417_1 <= _GEN_8055;
        end
      end else begin
        valid_417_1 <= _GEN_1956;
      end
    end else begin
      valid_417_1 <= _GEN_1956;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_418_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_418_0 <= _GEN_1445;
        end else begin
          valid_418_0 <= _GEN_8056;
        end
      end else begin
        valid_418_0 <= _GEN_1445;
      end
    end else begin
      valid_418_0 <= _GEN_1445;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_418_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_418_1 <= _GEN_1957;
        end else begin
          valid_418_1 <= _GEN_8057;
        end
      end else begin
        valid_418_1 <= _GEN_1957;
      end
    end else begin
      valid_418_1 <= _GEN_1957;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_419_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_419_0 <= _GEN_1446;
        end else begin
          valid_419_0 <= _GEN_8058;
        end
      end else begin
        valid_419_0 <= _GEN_1446;
      end
    end else begin
      valid_419_0 <= _GEN_1446;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_419_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_419_1 <= _GEN_1958;
        end else begin
          valid_419_1 <= _GEN_8059;
        end
      end else begin
        valid_419_1 <= _GEN_1958;
      end
    end else begin
      valid_419_1 <= _GEN_1958;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_420_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_420_0 <= _GEN_1447;
        end else begin
          valid_420_0 <= _GEN_8060;
        end
      end else begin
        valid_420_0 <= _GEN_1447;
      end
    end else begin
      valid_420_0 <= _GEN_1447;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_420_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_420_1 <= _GEN_1959;
        end else begin
          valid_420_1 <= _GEN_8061;
        end
      end else begin
        valid_420_1 <= _GEN_1959;
      end
    end else begin
      valid_420_1 <= _GEN_1959;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_421_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_421_0 <= _GEN_1448;
        end else begin
          valid_421_0 <= _GEN_8062;
        end
      end else begin
        valid_421_0 <= _GEN_1448;
      end
    end else begin
      valid_421_0 <= _GEN_1448;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_421_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_421_1 <= _GEN_1960;
        end else begin
          valid_421_1 <= _GEN_8063;
        end
      end else begin
        valid_421_1 <= _GEN_1960;
      end
    end else begin
      valid_421_1 <= _GEN_1960;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_422_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_422_0 <= _GEN_1449;
        end else begin
          valid_422_0 <= _GEN_8064;
        end
      end else begin
        valid_422_0 <= _GEN_1449;
      end
    end else begin
      valid_422_0 <= _GEN_1449;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_422_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_422_1 <= _GEN_1961;
        end else begin
          valid_422_1 <= _GEN_8065;
        end
      end else begin
        valid_422_1 <= _GEN_1961;
      end
    end else begin
      valid_422_1 <= _GEN_1961;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_423_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_423_0 <= _GEN_1450;
        end else begin
          valid_423_0 <= _GEN_8066;
        end
      end else begin
        valid_423_0 <= _GEN_1450;
      end
    end else begin
      valid_423_0 <= _GEN_1450;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_423_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_423_1 <= _GEN_1962;
        end else begin
          valid_423_1 <= _GEN_8067;
        end
      end else begin
        valid_423_1 <= _GEN_1962;
      end
    end else begin
      valid_423_1 <= _GEN_1962;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_424_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_424_0 <= _GEN_1451;
        end else begin
          valid_424_0 <= _GEN_8068;
        end
      end else begin
        valid_424_0 <= _GEN_1451;
      end
    end else begin
      valid_424_0 <= _GEN_1451;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_424_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_424_1 <= _GEN_1963;
        end else begin
          valid_424_1 <= _GEN_8069;
        end
      end else begin
        valid_424_1 <= _GEN_1963;
      end
    end else begin
      valid_424_1 <= _GEN_1963;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_425_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_425_0 <= _GEN_1452;
        end else begin
          valid_425_0 <= _GEN_8070;
        end
      end else begin
        valid_425_0 <= _GEN_1452;
      end
    end else begin
      valid_425_0 <= _GEN_1452;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_425_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_425_1 <= _GEN_1964;
        end else begin
          valid_425_1 <= _GEN_8071;
        end
      end else begin
        valid_425_1 <= _GEN_1964;
      end
    end else begin
      valid_425_1 <= _GEN_1964;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_426_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_426_0 <= _GEN_1453;
        end else begin
          valid_426_0 <= _GEN_8072;
        end
      end else begin
        valid_426_0 <= _GEN_1453;
      end
    end else begin
      valid_426_0 <= _GEN_1453;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_426_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_426_1 <= _GEN_1965;
        end else begin
          valid_426_1 <= _GEN_8073;
        end
      end else begin
        valid_426_1 <= _GEN_1965;
      end
    end else begin
      valid_426_1 <= _GEN_1965;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_427_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_427_0 <= _GEN_1454;
        end else begin
          valid_427_0 <= _GEN_8074;
        end
      end else begin
        valid_427_0 <= _GEN_1454;
      end
    end else begin
      valid_427_0 <= _GEN_1454;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_427_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_427_1 <= _GEN_1966;
        end else begin
          valid_427_1 <= _GEN_8075;
        end
      end else begin
        valid_427_1 <= _GEN_1966;
      end
    end else begin
      valid_427_1 <= _GEN_1966;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_428_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_428_0 <= _GEN_1455;
        end else begin
          valid_428_0 <= _GEN_8076;
        end
      end else begin
        valid_428_0 <= _GEN_1455;
      end
    end else begin
      valid_428_0 <= _GEN_1455;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_428_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_428_1 <= _GEN_1967;
        end else begin
          valid_428_1 <= _GEN_8077;
        end
      end else begin
        valid_428_1 <= _GEN_1967;
      end
    end else begin
      valid_428_1 <= _GEN_1967;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_429_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_429_0 <= _GEN_1456;
        end else begin
          valid_429_0 <= _GEN_8078;
        end
      end else begin
        valid_429_0 <= _GEN_1456;
      end
    end else begin
      valid_429_0 <= _GEN_1456;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_429_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_429_1 <= _GEN_1968;
        end else begin
          valid_429_1 <= _GEN_8079;
        end
      end else begin
        valid_429_1 <= _GEN_1968;
      end
    end else begin
      valid_429_1 <= _GEN_1968;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_430_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_430_0 <= _GEN_1457;
        end else begin
          valid_430_0 <= _GEN_8080;
        end
      end else begin
        valid_430_0 <= _GEN_1457;
      end
    end else begin
      valid_430_0 <= _GEN_1457;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_430_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_430_1 <= _GEN_1969;
        end else begin
          valid_430_1 <= _GEN_8081;
        end
      end else begin
        valid_430_1 <= _GEN_1969;
      end
    end else begin
      valid_430_1 <= _GEN_1969;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_431_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_431_0 <= _GEN_1458;
        end else begin
          valid_431_0 <= _GEN_8082;
        end
      end else begin
        valid_431_0 <= _GEN_1458;
      end
    end else begin
      valid_431_0 <= _GEN_1458;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_431_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_431_1 <= _GEN_1970;
        end else begin
          valid_431_1 <= _GEN_8083;
        end
      end else begin
        valid_431_1 <= _GEN_1970;
      end
    end else begin
      valid_431_1 <= _GEN_1970;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_432_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_432_0 <= _GEN_1459;
        end else begin
          valid_432_0 <= _GEN_8084;
        end
      end else begin
        valid_432_0 <= _GEN_1459;
      end
    end else begin
      valid_432_0 <= _GEN_1459;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_432_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_432_1 <= _GEN_1971;
        end else begin
          valid_432_1 <= _GEN_8085;
        end
      end else begin
        valid_432_1 <= _GEN_1971;
      end
    end else begin
      valid_432_1 <= _GEN_1971;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_433_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_433_0 <= _GEN_1460;
        end else begin
          valid_433_0 <= _GEN_8086;
        end
      end else begin
        valid_433_0 <= _GEN_1460;
      end
    end else begin
      valid_433_0 <= _GEN_1460;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_433_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_433_1 <= _GEN_1972;
        end else begin
          valid_433_1 <= _GEN_8087;
        end
      end else begin
        valid_433_1 <= _GEN_1972;
      end
    end else begin
      valid_433_1 <= _GEN_1972;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_434_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_434_0 <= _GEN_1461;
        end else begin
          valid_434_0 <= _GEN_8088;
        end
      end else begin
        valid_434_0 <= _GEN_1461;
      end
    end else begin
      valid_434_0 <= _GEN_1461;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_434_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_434_1 <= _GEN_1973;
        end else begin
          valid_434_1 <= _GEN_8089;
        end
      end else begin
        valid_434_1 <= _GEN_1973;
      end
    end else begin
      valid_434_1 <= _GEN_1973;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_435_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_435_0 <= _GEN_1462;
        end else begin
          valid_435_0 <= _GEN_8090;
        end
      end else begin
        valid_435_0 <= _GEN_1462;
      end
    end else begin
      valid_435_0 <= _GEN_1462;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_435_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_435_1 <= _GEN_1974;
        end else begin
          valid_435_1 <= _GEN_8091;
        end
      end else begin
        valid_435_1 <= _GEN_1974;
      end
    end else begin
      valid_435_1 <= _GEN_1974;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_436_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_436_0 <= _GEN_1463;
        end else begin
          valid_436_0 <= _GEN_8092;
        end
      end else begin
        valid_436_0 <= _GEN_1463;
      end
    end else begin
      valid_436_0 <= _GEN_1463;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_436_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_436_1 <= _GEN_1975;
        end else begin
          valid_436_1 <= _GEN_8093;
        end
      end else begin
        valid_436_1 <= _GEN_1975;
      end
    end else begin
      valid_436_1 <= _GEN_1975;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_437_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_437_0 <= _GEN_1464;
        end else begin
          valid_437_0 <= _GEN_8094;
        end
      end else begin
        valid_437_0 <= _GEN_1464;
      end
    end else begin
      valid_437_0 <= _GEN_1464;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_437_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_437_1 <= _GEN_1976;
        end else begin
          valid_437_1 <= _GEN_8095;
        end
      end else begin
        valid_437_1 <= _GEN_1976;
      end
    end else begin
      valid_437_1 <= _GEN_1976;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_438_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_438_0 <= _GEN_1465;
        end else begin
          valid_438_0 <= _GEN_8096;
        end
      end else begin
        valid_438_0 <= _GEN_1465;
      end
    end else begin
      valid_438_0 <= _GEN_1465;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_438_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_438_1 <= _GEN_1977;
        end else begin
          valid_438_1 <= _GEN_8097;
        end
      end else begin
        valid_438_1 <= _GEN_1977;
      end
    end else begin
      valid_438_1 <= _GEN_1977;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_439_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_439_0 <= _GEN_1466;
        end else begin
          valid_439_0 <= _GEN_8098;
        end
      end else begin
        valid_439_0 <= _GEN_1466;
      end
    end else begin
      valid_439_0 <= _GEN_1466;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_439_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_439_1 <= _GEN_1978;
        end else begin
          valid_439_1 <= _GEN_8099;
        end
      end else begin
        valid_439_1 <= _GEN_1978;
      end
    end else begin
      valid_439_1 <= _GEN_1978;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_440_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_440_0 <= _GEN_1467;
        end else begin
          valid_440_0 <= _GEN_8100;
        end
      end else begin
        valid_440_0 <= _GEN_1467;
      end
    end else begin
      valid_440_0 <= _GEN_1467;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_440_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_440_1 <= _GEN_1979;
        end else begin
          valid_440_1 <= _GEN_8101;
        end
      end else begin
        valid_440_1 <= _GEN_1979;
      end
    end else begin
      valid_440_1 <= _GEN_1979;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_441_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_441_0 <= _GEN_1468;
        end else begin
          valid_441_0 <= _GEN_8102;
        end
      end else begin
        valid_441_0 <= _GEN_1468;
      end
    end else begin
      valid_441_0 <= _GEN_1468;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_441_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_441_1 <= _GEN_1980;
        end else begin
          valid_441_1 <= _GEN_8103;
        end
      end else begin
        valid_441_1 <= _GEN_1980;
      end
    end else begin
      valid_441_1 <= _GEN_1980;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_442_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_442_0 <= _GEN_1469;
        end else begin
          valid_442_0 <= _GEN_8104;
        end
      end else begin
        valid_442_0 <= _GEN_1469;
      end
    end else begin
      valid_442_0 <= _GEN_1469;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_442_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_442_1 <= _GEN_1981;
        end else begin
          valid_442_1 <= _GEN_8105;
        end
      end else begin
        valid_442_1 <= _GEN_1981;
      end
    end else begin
      valid_442_1 <= _GEN_1981;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_443_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_443_0 <= _GEN_1470;
        end else begin
          valid_443_0 <= _GEN_8106;
        end
      end else begin
        valid_443_0 <= _GEN_1470;
      end
    end else begin
      valid_443_0 <= _GEN_1470;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_443_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_443_1 <= _GEN_1982;
        end else begin
          valid_443_1 <= _GEN_8107;
        end
      end else begin
        valid_443_1 <= _GEN_1982;
      end
    end else begin
      valid_443_1 <= _GEN_1982;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_444_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_444_0 <= _GEN_1471;
        end else begin
          valid_444_0 <= _GEN_8108;
        end
      end else begin
        valid_444_0 <= _GEN_1471;
      end
    end else begin
      valid_444_0 <= _GEN_1471;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_444_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_444_1 <= _GEN_1983;
        end else begin
          valid_444_1 <= _GEN_8109;
        end
      end else begin
        valid_444_1 <= _GEN_1983;
      end
    end else begin
      valid_444_1 <= _GEN_1983;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_445_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_445_0 <= _GEN_1472;
        end else begin
          valid_445_0 <= _GEN_8110;
        end
      end else begin
        valid_445_0 <= _GEN_1472;
      end
    end else begin
      valid_445_0 <= _GEN_1472;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_445_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_445_1 <= _GEN_1984;
        end else begin
          valid_445_1 <= _GEN_8111;
        end
      end else begin
        valid_445_1 <= _GEN_1984;
      end
    end else begin
      valid_445_1 <= _GEN_1984;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_446_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_446_0 <= _GEN_1473;
        end else begin
          valid_446_0 <= _GEN_8112;
        end
      end else begin
        valid_446_0 <= _GEN_1473;
      end
    end else begin
      valid_446_0 <= _GEN_1473;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_446_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_446_1 <= _GEN_1985;
        end else begin
          valid_446_1 <= _GEN_8113;
        end
      end else begin
        valid_446_1 <= _GEN_1985;
      end
    end else begin
      valid_446_1 <= _GEN_1985;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_447_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_447_0 <= _GEN_1474;
        end else begin
          valid_447_0 <= _GEN_8114;
        end
      end else begin
        valid_447_0 <= _GEN_1474;
      end
    end else begin
      valid_447_0 <= _GEN_1474;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_447_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_447_1 <= _GEN_1986;
        end else begin
          valid_447_1 <= _GEN_8115;
        end
      end else begin
        valid_447_1 <= _GEN_1986;
      end
    end else begin
      valid_447_1 <= _GEN_1986;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_448_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_448_0 <= _GEN_1475;
        end else begin
          valid_448_0 <= _GEN_8116;
        end
      end else begin
        valid_448_0 <= _GEN_1475;
      end
    end else begin
      valid_448_0 <= _GEN_1475;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_448_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_448_1 <= _GEN_1987;
        end else begin
          valid_448_1 <= _GEN_8117;
        end
      end else begin
        valid_448_1 <= _GEN_1987;
      end
    end else begin
      valid_448_1 <= _GEN_1987;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_449_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_449_0 <= _GEN_1476;
        end else begin
          valid_449_0 <= _GEN_8118;
        end
      end else begin
        valid_449_0 <= _GEN_1476;
      end
    end else begin
      valid_449_0 <= _GEN_1476;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_449_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_449_1 <= _GEN_1988;
        end else begin
          valid_449_1 <= _GEN_8119;
        end
      end else begin
        valid_449_1 <= _GEN_1988;
      end
    end else begin
      valid_449_1 <= _GEN_1988;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_450_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_450_0 <= _GEN_1477;
        end else begin
          valid_450_0 <= _GEN_8120;
        end
      end else begin
        valid_450_0 <= _GEN_1477;
      end
    end else begin
      valid_450_0 <= _GEN_1477;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_450_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_450_1 <= _GEN_1989;
        end else begin
          valid_450_1 <= _GEN_8121;
        end
      end else begin
        valid_450_1 <= _GEN_1989;
      end
    end else begin
      valid_450_1 <= _GEN_1989;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_451_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_451_0 <= _GEN_1478;
        end else begin
          valid_451_0 <= _GEN_8122;
        end
      end else begin
        valid_451_0 <= _GEN_1478;
      end
    end else begin
      valid_451_0 <= _GEN_1478;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_451_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_451_1 <= _GEN_1990;
        end else begin
          valid_451_1 <= _GEN_8123;
        end
      end else begin
        valid_451_1 <= _GEN_1990;
      end
    end else begin
      valid_451_1 <= _GEN_1990;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_452_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_452_0 <= _GEN_1479;
        end else begin
          valid_452_0 <= _GEN_8124;
        end
      end else begin
        valid_452_0 <= _GEN_1479;
      end
    end else begin
      valid_452_0 <= _GEN_1479;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_452_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_452_1 <= _GEN_1991;
        end else begin
          valid_452_1 <= _GEN_8125;
        end
      end else begin
        valid_452_1 <= _GEN_1991;
      end
    end else begin
      valid_452_1 <= _GEN_1991;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_453_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_453_0 <= _GEN_1480;
        end else begin
          valid_453_0 <= _GEN_8126;
        end
      end else begin
        valid_453_0 <= _GEN_1480;
      end
    end else begin
      valid_453_0 <= _GEN_1480;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_453_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_453_1 <= _GEN_1992;
        end else begin
          valid_453_1 <= _GEN_8127;
        end
      end else begin
        valid_453_1 <= _GEN_1992;
      end
    end else begin
      valid_453_1 <= _GEN_1992;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_454_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_454_0 <= _GEN_1481;
        end else begin
          valid_454_0 <= _GEN_8128;
        end
      end else begin
        valid_454_0 <= _GEN_1481;
      end
    end else begin
      valid_454_0 <= _GEN_1481;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_454_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_454_1 <= _GEN_1993;
        end else begin
          valid_454_1 <= _GEN_8129;
        end
      end else begin
        valid_454_1 <= _GEN_1993;
      end
    end else begin
      valid_454_1 <= _GEN_1993;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_455_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_455_0 <= _GEN_1482;
        end else begin
          valid_455_0 <= _GEN_8130;
        end
      end else begin
        valid_455_0 <= _GEN_1482;
      end
    end else begin
      valid_455_0 <= _GEN_1482;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_455_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_455_1 <= _GEN_1994;
        end else begin
          valid_455_1 <= _GEN_8131;
        end
      end else begin
        valid_455_1 <= _GEN_1994;
      end
    end else begin
      valid_455_1 <= _GEN_1994;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_456_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_456_0 <= _GEN_1483;
        end else begin
          valid_456_0 <= _GEN_8132;
        end
      end else begin
        valid_456_0 <= _GEN_1483;
      end
    end else begin
      valid_456_0 <= _GEN_1483;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_456_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_456_1 <= _GEN_1995;
        end else begin
          valid_456_1 <= _GEN_8133;
        end
      end else begin
        valid_456_1 <= _GEN_1995;
      end
    end else begin
      valid_456_1 <= _GEN_1995;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_457_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_457_0 <= _GEN_1484;
        end else begin
          valid_457_0 <= _GEN_8134;
        end
      end else begin
        valid_457_0 <= _GEN_1484;
      end
    end else begin
      valid_457_0 <= _GEN_1484;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_457_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_457_1 <= _GEN_1996;
        end else begin
          valid_457_1 <= _GEN_8135;
        end
      end else begin
        valid_457_1 <= _GEN_1996;
      end
    end else begin
      valid_457_1 <= _GEN_1996;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_458_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_458_0 <= _GEN_1485;
        end else begin
          valid_458_0 <= _GEN_8136;
        end
      end else begin
        valid_458_0 <= _GEN_1485;
      end
    end else begin
      valid_458_0 <= _GEN_1485;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_458_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_458_1 <= _GEN_1997;
        end else begin
          valid_458_1 <= _GEN_8137;
        end
      end else begin
        valid_458_1 <= _GEN_1997;
      end
    end else begin
      valid_458_1 <= _GEN_1997;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_459_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_459_0 <= _GEN_1486;
        end else begin
          valid_459_0 <= _GEN_8138;
        end
      end else begin
        valid_459_0 <= _GEN_1486;
      end
    end else begin
      valid_459_0 <= _GEN_1486;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_459_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_459_1 <= _GEN_1998;
        end else begin
          valid_459_1 <= _GEN_8139;
        end
      end else begin
        valid_459_1 <= _GEN_1998;
      end
    end else begin
      valid_459_1 <= _GEN_1998;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_460_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_460_0 <= _GEN_1487;
        end else begin
          valid_460_0 <= _GEN_8140;
        end
      end else begin
        valid_460_0 <= _GEN_1487;
      end
    end else begin
      valid_460_0 <= _GEN_1487;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_460_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_460_1 <= _GEN_1999;
        end else begin
          valid_460_1 <= _GEN_8141;
        end
      end else begin
        valid_460_1 <= _GEN_1999;
      end
    end else begin
      valid_460_1 <= _GEN_1999;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_461_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_461_0 <= _GEN_1488;
        end else begin
          valid_461_0 <= _GEN_8142;
        end
      end else begin
        valid_461_0 <= _GEN_1488;
      end
    end else begin
      valid_461_0 <= _GEN_1488;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_461_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_461_1 <= _GEN_2000;
        end else begin
          valid_461_1 <= _GEN_8143;
        end
      end else begin
        valid_461_1 <= _GEN_2000;
      end
    end else begin
      valid_461_1 <= _GEN_2000;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_462_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_462_0 <= _GEN_1489;
        end else begin
          valid_462_0 <= _GEN_8144;
        end
      end else begin
        valid_462_0 <= _GEN_1489;
      end
    end else begin
      valid_462_0 <= _GEN_1489;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_462_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_462_1 <= _GEN_2001;
        end else begin
          valid_462_1 <= _GEN_8145;
        end
      end else begin
        valid_462_1 <= _GEN_2001;
      end
    end else begin
      valid_462_1 <= _GEN_2001;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_463_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_463_0 <= _GEN_1490;
        end else begin
          valid_463_0 <= _GEN_8146;
        end
      end else begin
        valid_463_0 <= _GEN_1490;
      end
    end else begin
      valid_463_0 <= _GEN_1490;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_463_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_463_1 <= _GEN_2002;
        end else begin
          valid_463_1 <= _GEN_8147;
        end
      end else begin
        valid_463_1 <= _GEN_2002;
      end
    end else begin
      valid_463_1 <= _GEN_2002;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_464_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_464_0 <= _GEN_1491;
        end else begin
          valid_464_0 <= _GEN_8148;
        end
      end else begin
        valid_464_0 <= _GEN_1491;
      end
    end else begin
      valid_464_0 <= _GEN_1491;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_464_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_464_1 <= _GEN_2003;
        end else begin
          valid_464_1 <= _GEN_8149;
        end
      end else begin
        valid_464_1 <= _GEN_2003;
      end
    end else begin
      valid_464_1 <= _GEN_2003;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_465_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_465_0 <= _GEN_1492;
        end else begin
          valid_465_0 <= _GEN_8150;
        end
      end else begin
        valid_465_0 <= _GEN_1492;
      end
    end else begin
      valid_465_0 <= _GEN_1492;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_465_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_465_1 <= _GEN_2004;
        end else begin
          valid_465_1 <= _GEN_8151;
        end
      end else begin
        valid_465_1 <= _GEN_2004;
      end
    end else begin
      valid_465_1 <= _GEN_2004;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_466_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_466_0 <= _GEN_1493;
        end else begin
          valid_466_0 <= _GEN_8152;
        end
      end else begin
        valid_466_0 <= _GEN_1493;
      end
    end else begin
      valid_466_0 <= _GEN_1493;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_466_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_466_1 <= _GEN_2005;
        end else begin
          valid_466_1 <= _GEN_8153;
        end
      end else begin
        valid_466_1 <= _GEN_2005;
      end
    end else begin
      valid_466_1 <= _GEN_2005;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_467_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_467_0 <= _GEN_1494;
        end else begin
          valid_467_0 <= _GEN_8154;
        end
      end else begin
        valid_467_0 <= _GEN_1494;
      end
    end else begin
      valid_467_0 <= _GEN_1494;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_467_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_467_1 <= _GEN_2006;
        end else begin
          valid_467_1 <= _GEN_8155;
        end
      end else begin
        valid_467_1 <= _GEN_2006;
      end
    end else begin
      valid_467_1 <= _GEN_2006;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_468_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_468_0 <= _GEN_1495;
        end else begin
          valid_468_0 <= _GEN_8156;
        end
      end else begin
        valid_468_0 <= _GEN_1495;
      end
    end else begin
      valid_468_0 <= _GEN_1495;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_468_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_468_1 <= _GEN_2007;
        end else begin
          valid_468_1 <= _GEN_8157;
        end
      end else begin
        valid_468_1 <= _GEN_2007;
      end
    end else begin
      valid_468_1 <= _GEN_2007;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_469_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_469_0 <= _GEN_1496;
        end else begin
          valid_469_0 <= _GEN_8158;
        end
      end else begin
        valid_469_0 <= _GEN_1496;
      end
    end else begin
      valid_469_0 <= _GEN_1496;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_469_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_469_1 <= _GEN_2008;
        end else begin
          valid_469_1 <= _GEN_8159;
        end
      end else begin
        valid_469_1 <= _GEN_2008;
      end
    end else begin
      valid_469_1 <= _GEN_2008;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_470_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_470_0 <= _GEN_1497;
        end else begin
          valid_470_0 <= _GEN_8160;
        end
      end else begin
        valid_470_0 <= _GEN_1497;
      end
    end else begin
      valid_470_0 <= _GEN_1497;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_470_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_470_1 <= _GEN_2009;
        end else begin
          valid_470_1 <= _GEN_8161;
        end
      end else begin
        valid_470_1 <= _GEN_2009;
      end
    end else begin
      valid_470_1 <= _GEN_2009;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_471_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_471_0 <= _GEN_1498;
        end else begin
          valid_471_0 <= _GEN_8162;
        end
      end else begin
        valid_471_0 <= _GEN_1498;
      end
    end else begin
      valid_471_0 <= _GEN_1498;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_471_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_471_1 <= _GEN_2010;
        end else begin
          valid_471_1 <= _GEN_8163;
        end
      end else begin
        valid_471_1 <= _GEN_2010;
      end
    end else begin
      valid_471_1 <= _GEN_2010;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_472_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_472_0 <= _GEN_1499;
        end else begin
          valid_472_0 <= _GEN_8164;
        end
      end else begin
        valid_472_0 <= _GEN_1499;
      end
    end else begin
      valid_472_0 <= _GEN_1499;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_472_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_472_1 <= _GEN_2011;
        end else begin
          valid_472_1 <= _GEN_8165;
        end
      end else begin
        valid_472_1 <= _GEN_2011;
      end
    end else begin
      valid_472_1 <= _GEN_2011;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_473_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_473_0 <= _GEN_1500;
        end else begin
          valid_473_0 <= _GEN_8166;
        end
      end else begin
        valid_473_0 <= _GEN_1500;
      end
    end else begin
      valid_473_0 <= _GEN_1500;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_473_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_473_1 <= _GEN_2012;
        end else begin
          valid_473_1 <= _GEN_8167;
        end
      end else begin
        valid_473_1 <= _GEN_2012;
      end
    end else begin
      valid_473_1 <= _GEN_2012;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_474_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_474_0 <= _GEN_1501;
        end else begin
          valid_474_0 <= _GEN_8168;
        end
      end else begin
        valid_474_0 <= _GEN_1501;
      end
    end else begin
      valid_474_0 <= _GEN_1501;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_474_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_474_1 <= _GEN_2013;
        end else begin
          valid_474_1 <= _GEN_8169;
        end
      end else begin
        valid_474_1 <= _GEN_2013;
      end
    end else begin
      valid_474_1 <= _GEN_2013;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_475_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_475_0 <= _GEN_1502;
        end else begin
          valid_475_0 <= _GEN_8170;
        end
      end else begin
        valid_475_0 <= _GEN_1502;
      end
    end else begin
      valid_475_0 <= _GEN_1502;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_475_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_475_1 <= _GEN_2014;
        end else begin
          valid_475_1 <= _GEN_8171;
        end
      end else begin
        valid_475_1 <= _GEN_2014;
      end
    end else begin
      valid_475_1 <= _GEN_2014;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_476_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_476_0 <= _GEN_1503;
        end else begin
          valid_476_0 <= _GEN_8172;
        end
      end else begin
        valid_476_0 <= _GEN_1503;
      end
    end else begin
      valid_476_0 <= _GEN_1503;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_476_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_476_1 <= _GEN_2015;
        end else begin
          valid_476_1 <= _GEN_8173;
        end
      end else begin
        valid_476_1 <= _GEN_2015;
      end
    end else begin
      valid_476_1 <= _GEN_2015;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_477_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_477_0 <= _GEN_1504;
        end else begin
          valid_477_0 <= _GEN_8174;
        end
      end else begin
        valid_477_0 <= _GEN_1504;
      end
    end else begin
      valid_477_0 <= _GEN_1504;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_477_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_477_1 <= _GEN_2016;
        end else begin
          valid_477_1 <= _GEN_8175;
        end
      end else begin
        valid_477_1 <= _GEN_2016;
      end
    end else begin
      valid_477_1 <= _GEN_2016;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_478_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_478_0 <= _GEN_1505;
        end else begin
          valid_478_0 <= _GEN_8176;
        end
      end else begin
        valid_478_0 <= _GEN_1505;
      end
    end else begin
      valid_478_0 <= _GEN_1505;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_478_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_478_1 <= _GEN_2017;
        end else begin
          valid_478_1 <= _GEN_8177;
        end
      end else begin
        valid_478_1 <= _GEN_2017;
      end
    end else begin
      valid_478_1 <= _GEN_2017;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_479_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_479_0 <= _GEN_1506;
        end else begin
          valid_479_0 <= _GEN_8178;
        end
      end else begin
        valid_479_0 <= _GEN_1506;
      end
    end else begin
      valid_479_0 <= _GEN_1506;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_479_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_479_1 <= _GEN_2018;
        end else begin
          valid_479_1 <= _GEN_8179;
        end
      end else begin
        valid_479_1 <= _GEN_2018;
      end
    end else begin
      valid_479_1 <= _GEN_2018;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_480_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_480_0 <= _GEN_1507;
        end else begin
          valid_480_0 <= _GEN_8180;
        end
      end else begin
        valid_480_0 <= _GEN_1507;
      end
    end else begin
      valid_480_0 <= _GEN_1507;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_480_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_480_1 <= _GEN_2019;
        end else begin
          valid_480_1 <= _GEN_8181;
        end
      end else begin
        valid_480_1 <= _GEN_2019;
      end
    end else begin
      valid_480_1 <= _GEN_2019;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_481_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_481_0 <= _GEN_1508;
        end else begin
          valid_481_0 <= _GEN_8182;
        end
      end else begin
        valid_481_0 <= _GEN_1508;
      end
    end else begin
      valid_481_0 <= _GEN_1508;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_481_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_481_1 <= _GEN_2020;
        end else begin
          valid_481_1 <= _GEN_8183;
        end
      end else begin
        valid_481_1 <= _GEN_2020;
      end
    end else begin
      valid_481_1 <= _GEN_2020;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_482_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_482_0 <= _GEN_1509;
        end else begin
          valid_482_0 <= _GEN_8184;
        end
      end else begin
        valid_482_0 <= _GEN_1509;
      end
    end else begin
      valid_482_0 <= _GEN_1509;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_482_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_482_1 <= _GEN_2021;
        end else begin
          valid_482_1 <= _GEN_8185;
        end
      end else begin
        valid_482_1 <= _GEN_2021;
      end
    end else begin
      valid_482_1 <= _GEN_2021;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_483_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_483_0 <= _GEN_1510;
        end else begin
          valid_483_0 <= _GEN_8186;
        end
      end else begin
        valid_483_0 <= _GEN_1510;
      end
    end else begin
      valid_483_0 <= _GEN_1510;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_483_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_483_1 <= _GEN_2022;
        end else begin
          valid_483_1 <= _GEN_8187;
        end
      end else begin
        valid_483_1 <= _GEN_2022;
      end
    end else begin
      valid_483_1 <= _GEN_2022;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_484_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_484_0 <= _GEN_1511;
        end else begin
          valid_484_0 <= _GEN_8188;
        end
      end else begin
        valid_484_0 <= _GEN_1511;
      end
    end else begin
      valid_484_0 <= _GEN_1511;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_484_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_484_1 <= _GEN_2023;
        end else begin
          valid_484_1 <= _GEN_8189;
        end
      end else begin
        valid_484_1 <= _GEN_2023;
      end
    end else begin
      valid_484_1 <= _GEN_2023;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_485_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_485_0 <= _GEN_1512;
        end else begin
          valid_485_0 <= _GEN_8190;
        end
      end else begin
        valid_485_0 <= _GEN_1512;
      end
    end else begin
      valid_485_0 <= _GEN_1512;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_485_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_485_1 <= _GEN_2024;
        end else begin
          valid_485_1 <= _GEN_8191;
        end
      end else begin
        valid_485_1 <= _GEN_2024;
      end
    end else begin
      valid_485_1 <= _GEN_2024;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_486_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_486_0 <= _GEN_1513;
        end else begin
          valid_486_0 <= _GEN_8192;
        end
      end else begin
        valid_486_0 <= _GEN_1513;
      end
    end else begin
      valid_486_0 <= _GEN_1513;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_486_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_486_1 <= _GEN_2025;
        end else begin
          valid_486_1 <= _GEN_8193;
        end
      end else begin
        valid_486_1 <= _GEN_2025;
      end
    end else begin
      valid_486_1 <= _GEN_2025;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_487_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_487_0 <= _GEN_1514;
        end else begin
          valid_487_0 <= _GEN_8194;
        end
      end else begin
        valid_487_0 <= _GEN_1514;
      end
    end else begin
      valid_487_0 <= _GEN_1514;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_487_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_487_1 <= _GEN_2026;
        end else begin
          valid_487_1 <= _GEN_8195;
        end
      end else begin
        valid_487_1 <= _GEN_2026;
      end
    end else begin
      valid_487_1 <= _GEN_2026;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_488_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_488_0 <= _GEN_1515;
        end else begin
          valid_488_0 <= _GEN_8196;
        end
      end else begin
        valid_488_0 <= _GEN_1515;
      end
    end else begin
      valid_488_0 <= _GEN_1515;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_488_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_488_1 <= _GEN_2027;
        end else begin
          valid_488_1 <= _GEN_8197;
        end
      end else begin
        valid_488_1 <= _GEN_2027;
      end
    end else begin
      valid_488_1 <= _GEN_2027;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_489_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_489_0 <= _GEN_1516;
        end else begin
          valid_489_0 <= _GEN_8198;
        end
      end else begin
        valid_489_0 <= _GEN_1516;
      end
    end else begin
      valid_489_0 <= _GEN_1516;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_489_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_489_1 <= _GEN_2028;
        end else begin
          valid_489_1 <= _GEN_8199;
        end
      end else begin
        valid_489_1 <= _GEN_2028;
      end
    end else begin
      valid_489_1 <= _GEN_2028;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_490_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_490_0 <= _GEN_1517;
        end else begin
          valid_490_0 <= _GEN_8200;
        end
      end else begin
        valid_490_0 <= _GEN_1517;
      end
    end else begin
      valid_490_0 <= _GEN_1517;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_490_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_490_1 <= _GEN_2029;
        end else begin
          valid_490_1 <= _GEN_8201;
        end
      end else begin
        valid_490_1 <= _GEN_2029;
      end
    end else begin
      valid_490_1 <= _GEN_2029;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_491_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_491_0 <= _GEN_1518;
        end else begin
          valid_491_0 <= _GEN_8202;
        end
      end else begin
        valid_491_0 <= _GEN_1518;
      end
    end else begin
      valid_491_0 <= _GEN_1518;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_491_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_491_1 <= _GEN_2030;
        end else begin
          valid_491_1 <= _GEN_8203;
        end
      end else begin
        valid_491_1 <= _GEN_2030;
      end
    end else begin
      valid_491_1 <= _GEN_2030;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_492_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_492_0 <= _GEN_1519;
        end else begin
          valid_492_0 <= _GEN_8204;
        end
      end else begin
        valid_492_0 <= _GEN_1519;
      end
    end else begin
      valid_492_0 <= _GEN_1519;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_492_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_492_1 <= _GEN_2031;
        end else begin
          valid_492_1 <= _GEN_8205;
        end
      end else begin
        valid_492_1 <= _GEN_2031;
      end
    end else begin
      valid_492_1 <= _GEN_2031;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_493_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_493_0 <= _GEN_1520;
        end else begin
          valid_493_0 <= _GEN_8206;
        end
      end else begin
        valid_493_0 <= _GEN_1520;
      end
    end else begin
      valid_493_0 <= _GEN_1520;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_493_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_493_1 <= _GEN_2032;
        end else begin
          valid_493_1 <= _GEN_8207;
        end
      end else begin
        valid_493_1 <= _GEN_2032;
      end
    end else begin
      valid_493_1 <= _GEN_2032;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_494_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_494_0 <= _GEN_1521;
        end else begin
          valid_494_0 <= _GEN_8208;
        end
      end else begin
        valid_494_0 <= _GEN_1521;
      end
    end else begin
      valid_494_0 <= _GEN_1521;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_494_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_494_1 <= _GEN_2033;
        end else begin
          valid_494_1 <= _GEN_8209;
        end
      end else begin
        valid_494_1 <= _GEN_2033;
      end
    end else begin
      valid_494_1 <= _GEN_2033;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_495_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_495_0 <= _GEN_1522;
        end else begin
          valid_495_0 <= _GEN_8210;
        end
      end else begin
        valid_495_0 <= _GEN_1522;
      end
    end else begin
      valid_495_0 <= _GEN_1522;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_495_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_495_1 <= _GEN_2034;
        end else begin
          valid_495_1 <= _GEN_8211;
        end
      end else begin
        valid_495_1 <= _GEN_2034;
      end
    end else begin
      valid_495_1 <= _GEN_2034;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_496_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_496_0 <= _GEN_1523;
        end else begin
          valid_496_0 <= _GEN_8212;
        end
      end else begin
        valid_496_0 <= _GEN_1523;
      end
    end else begin
      valid_496_0 <= _GEN_1523;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_496_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_496_1 <= _GEN_2035;
        end else begin
          valid_496_1 <= _GEN_8213;
        end
      end else begin
        valid_496_1 <= _GEN_2035;
      end
    end else begin
      valid_496_1 <= _GEN_2035;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_497_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_497_0 <= _GEN_1524;
        end else begin
          valid_497_0 <= _GEN_8214;
        end
      end else begin
        valid_497_0 <= _GEN_1524;
      end
    end else begin
      valid_497_0 <= _GEN_1524;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_497_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_497_1 <= _GEN_2036;
        end else begin
          valid_497_1 <= _GEN_8215;
        end
      end else begin
        valid_497_1 <= _GEN_2036;
      end
    end else begin
      valid_497_1 <= _GEN_2036;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_498_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_498_0 <= _GEN_1525;
        end else begin
          valid_498_0 <= _GEN_8216;
        end
      end else begin
        valid_498_0 <= _GEN_1525;
      end
    end else begin
      valid_498_0 <= _GEN_1525;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_498_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_498_1 <= _GEN_2037;
        end else begin
          valid_498_1 <= _GEN_8217;
        end
      end else begin
        valid_498_1 <= _GEN_2037;
      end
    end else begin
      valid_498_1 <= _GEN_2037;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_499_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_499_0 <= _GEN_1526;
        end else begin
          valid_499_0 <= _GEN_8218;
        end
      end else begin
        valid_499_0 <= _GEN_1526;
      end
    end else begin
      valid_499_0 <= _GEN_1526;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_499_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_499_1 <= _GEN_2038;
        end else begin
          valid_499_1 <= _GEN_8219;
        end
      end else begin
        valid_499_1 <= _GEN_2038;
      end
    end else begin
      valid_499_1 <= _GEN_2038;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_500_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_500_0 <= _GEN_1527;
        end else begin
          valid_500_0 <= _GEN_8220;
        end
      end else begin
        valid_500_0 <= _GEN_1527;
      end
    end else begin
      valid_500_0 <= _GEN_1527;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_500_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_500_1 <= _GEN_2039;
        end else begin
          valid_500_1 <= _GEN_8221;
        end
      end else begin
        valid_500_1 <= _GEN_2039;
      end
    end else begin
      valid_500_1 <= _GEN_2039;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_501_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_501_0 <= _GEN_1528;
        end else begin
          valid_501_0 <= _GEN_8222;
        end
      end else begin
        valid_501_0 <= _GEN_1528;
      end
    end else begin
      valid_501_0 <= _GEN_1528;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_501_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_501_1 <= _GEN_2040;
        end else begin
          valid_501_1 <= _GEN_8223;
        end
      end else begin
        valid_501_1 <= _GEN_2040;
      end
    end else begin
      valid_501_1 <= _GEN_2040;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_502_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_502_0 <= _GEN_1529;
        end else begin
          valid_502_0 <= _GEN_8224;
        end
      end else begin
        valid_502_0 <= _GEN_1529;
      end
    end else begin
      valid_502_0 <= _GEN_1529;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_502_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_502_1 <= _GEN_2041;
        end else begin
          valid_502_1 <= _GEN_8225;
        end
      end else begin
        valid_502_1 <= _GEN_2041;
      end
    end else begin
      valid_502_1 <= _GEN_2041;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_503_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_503_0 <= _GEN_1530;
        end else begin
          valid_503_0 <= _GEN_8226;
        end
      end else begin
        valid_503_0 <= _GEN_1530;
      end
    end else begin
      valid_503_0 <= _GEN_1530;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_503_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_503_1 <= _GEN_2042;
        end else begin
          valid_503_1 <= _GEN_8227;
        end
      end else begin
        valid_503_1 <= _GEN_2042;
      end
    end else begin
      valid_503_1 <= _GEN_2042;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_504_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_504_0 <= _GEN_1531;
        end else begin
          valid_504_0 <= _GEN_8228;
        end
      end else begin
        valid_504_0 <= _GEN_1531;
      end
    end else begin
      valid_504_0 <= _GEN_1531;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_504_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_504_1 <= _GEN_2043;
        end else begin
          valid_504_1 <= _GEN_8229;
        end
      end else begin
        valid_504_1 <= _GEN_2043;
      end
    end else begin
      valid_504_1 <= _GEN_2043;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_505_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_505_0 <= _GEN_1532;
        end else begin
          valid_505_0 <= _GEN_8230;
        end
      end else begin
        valid_505_0 <= _GEN_1532;
      end
    end else begin
      valid_505_0 <= _GEN_1532;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_505_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_505_1 <= _GEN_2044;
        end else begin
          valid_505_1 <= _GEN_8231;
        end
      end else begin
        valid_505_1 <= _GEN_2044;
      end
    end else begin
      valid_505_1 <= _GEN_2044;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_506_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_506_0 <= _GEN_1533;
        end else begin
          valid_506_0 <= _GEN_8232;
        end
      end else begin
        valid_506_0 <= _GEN_1533;
      end
    end else begin
      valid_506_0 <= _GEN_1533;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_506_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_506_1 <= _GEN_2045;
        end else begin
          valid_506_1 <= _GEN_8233;
        end
      end else begin
        valid_506_1 <= _GEN_2045;
      end
    end else begin
      valid_506_1 <= _GEN_2045;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_507_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_507_0 <= _GEN_1534;
        end else begin
          valid_507_0 <= _GEN_8234;
        end
      end else begin
        valid_507_0 <= _GEN_1534;
      end
    end else begin
      valid_507_0 <= _GEN_1534;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_507_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_507_1 <= _GEN_2046;
        end else begin
          valid_507_1 <= _GEN_8235;
        end
      end else begin
        valid_507_1 <= _GEN_2046;
      end
    end else begin
      valid_507_1 <= _GEN_2046;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_508_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_508_0 <= _GEN_1535;
        end else begin
          valid_508_0 <= _GEN_8236;
        end
      end else begin
        valid_508_0 <= _GEN_1535;
      end
    end else begin
      valid_508_0 <= _GEN_1535;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_508_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_508_1 <= _GEN_2047;
        end else begin
          valid_508_1 <= _GEN_8237;
        end
      end else begin
        valid_508_1 <= _GEN_2047;
      end
    end else begin
      valid_508_1 <= _GEN_2047;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_509_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_509_0 <= _GEN_1536;
        end else begin
          valid_509_0 <= _GEN_8238;
        end
      end else begin
        valid_509_0 <= _GEN_1536;
      end
    end else begin
      valid_509_0 <= _GEN_1536;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_509_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_509_1 <= _GEN_2048;
        end else begin
          valid_509_1 <= _GEN_8239;
        end
      end else begin
        valid_509_1 <= _GEN_2048;
      end
    end else begin
      valid_509_1 <= _GEN_2048;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_510_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_510_0 <= _GEN_1537;
        end else begin
          valid_510_0 <= _GEN_8240;
        end
      end else begin
        valid_510_0 <= _GEN_1537;
      end
    end else begin
      valid_510_0 <= _GEN_1537;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_510_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_510_1 <= _GEN_2049;
        end else begin
          valid_510_1 <= _GEN_8241;
        end
      end else begin
        valid_510_1 <= _GEN_2049;
      end
    end else begin
      valid_510_1 <= _GEN_2049;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_511_0 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_511_0 <= _GEN_1538;
        end else begin
          valid_511_0 <= _GEN_8242;
        end
      end else begin
        valid_511_0 <= _GEN_1538;
      end
    end else begin
      valid_511_0 <= _GEN_1538;
    end
    if (reset) begin // @[ICache.scala 52:22]
      valid_511_1 <= 1'h0; // @[ICache.scala 52:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (_io_cpu_tlb2_vpn_T_2) begin // @[ICache.scala 167:31]
          valid_511_1 <= _GEN_2050;
        end else begin
          valid_511_1 <= _GEN_8243;
        end
      end else begin
        valid_511_1 <= _GEN_2050;
      end
    end else begin
      valid_511_1 <= _GEN_2050;
    end
    if (reset) begin // @[ICache.scala 61:27]
      data_wstrb_0_0 <= 4'h0; // @[ICache.scala 61:27]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          data_wstrb_0_0 <= _GEN_7213;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        data_wstrb_0_0 <= _GEN_11941;
      end
    end
    if (reset) begin // @[ICache.scala 61:27]
      data_wstrb_0_1 <= 4'h0; // @[ICache.scala 61:27]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          data_wstrb_0_1 <= _GEN_7215;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        data_wstrb_0_1 <= _GEN_11943;
      end
    end
    if (reset) begin // @[ICache.scala 61:27]
      data_wstrb_1_0 <= 4'h0; // @[ICache.scala 61:27]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          data_wstrb_1_0 <= _GEN_7214;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        data_wstrb_1_0 <= _GEN_11942;
      end
    end
    if (reset) begin // @[ICache.scala 61:27]
      data_wstrb_1_1 <= 4'h0; // @[ICache.scala 61:27]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          data_wstrb_1_1 <= _GEN_7216;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        data_wstrb_1_1 <= _GEN_11944;
      end
    end
    if (reset) begin // @[ICache.scala 64:26]
      tag_wstrb_0 <= 1'h0; // @[ICache.scala 64:26]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          tag_wstrb_0 <= _GEN_7217;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        tag_wstrb_0 <= _GEN_11945;
      end
    end
    if (reset) begin // @[ICache.scala 64:26]
      tag_wstrb_1 <= 1'h0; // @[ICache.scala 64:26]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          tag_wstrb_1 <= _GEN_7218;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        tag_wstrb_1 <= _GEN_11946;
      end
    end
    if (reset) begin // @[ICache.scala 65:26]
      tag_wdata <= 20'h0; // @[ICache.scala 65:26]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          tag_wdata <= _GEN_7219;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_0 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_0 <= _GEN_8245;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_1 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_1 <= _GEN_8246;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_2 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_2 <= _GEN_8247;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_3 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_3 <= _GEN_8248;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_4 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_4 <= _GEN_8249;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_5 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_5 <= _GEN_8250;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_6 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_6 <= _GEN_8251;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_7 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_7 <= _GEN_8252;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_8 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_8 <= _GEN_8253;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_9 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_9 <= _GEN_8254;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_10 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_10 <= _GEN_8255;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_11 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_11 <= _GEN_8256;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_12 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_12 <= _GEN_8257;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_13 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_13 <= _GEN_8258;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_14 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_14 <= _GEN_8259;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_15 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_15 <= _GEN_8260;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_16 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_16 <= _GEN_8261;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_17 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_17 <= _GEN_8262;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_18 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_18 <= _GEN_8263;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_19 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_19 <= _GEN_8264;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_20 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_20 <= _GEN_8265;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_21 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_21 <= _GEN_8266;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_22 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_22 <= _GEN_8267;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_23 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_23 <= _GEN_8268;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_24 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_24 <= _GEN_8269;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_25 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_25 <= _GEN_8270;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_26 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_26 <= _GEN_8271;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_27 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_27 <= _GEN_8272;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_28 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_28 <= _GEN_8273;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_29 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_29 <= _GEN_8274;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_30 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_30 <= _GEN_8275;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_31 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_31 <= _GEN_8276;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_32 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_32 <= _GEN_8277;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_33 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_33 <= _GEN_8278;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_34 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_34 <= _GEN_8279;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_35 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_35 <= _GEN_8280;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_36 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_36 <= _GEN_8281;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_37 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_37 <= _GEN_8282;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_38 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_38 <= _GEN_8283;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_39 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_39 <= _GEN_8284;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_40 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_40 <= _GEN_8285;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_41 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_41 <= _GEN_8286;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_42 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_42 <= _GEN_8287;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_43 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_43 <= _GEN_8288;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_44 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_44 <= _GEN_8289;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_45 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_45 <= _GEN_8290;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_46 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_46 <= _GEN_8291;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_47 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_47 <= _GEN_8292;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_48 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_48 <= _GEN_8293;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_49 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_49 <= _GEN_8294;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_50 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_50 <= _GEN_8295;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_51 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_51 <= _GEN_8296;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_52 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_52 <= _GEN_8297;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_53 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_53 <= _GEN_8298;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_54 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_54 <= _GEN_8299;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_55 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_55 <= _GEN_8300;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_56 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_56 <= _GEN_8301;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_57 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_57 <= _GEN_8302;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_58 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_58 <= _GEN_8303;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_59 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_59 <= _GEN_8304;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_60 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_60 <= _GEN_8305;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_61 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_61 <= _GEN_8306;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_62 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_62 <= _GEN_8307;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_63 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_63 <= _GEN_8308;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_64 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_64 <= _GEN_8309;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_65 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_65 <= _GEN_8310;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_66 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_66 <= _GEN_8311;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_67 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_67 <= _GEN_8312;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_68 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_68 <= _GEN_8313;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_69 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_69 <= _GEN_8314;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_70 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_70 <= _GEN_8315;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_71 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_71 <= _GEN_8316;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_72 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_72 <= _GEN_8317;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_73 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_73 <= _GEN_8318;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_74 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_74 <= _GEN_8319;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_75 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_75 <= _GEN_8320;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_76 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_76 <= _GEN_8321;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_77 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_77 <= _GEN_8322;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_78 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_78 <= _GEN_8323;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_79 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_79 <= _GEN_8324;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_80 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_80 <= _GEN_8325;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_81 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_81 <= _GEN_8326;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_82 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_82 <= _GEN_8327;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_83 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_83 <= _GEN_8328;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_84 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_84 <= _GEN_8329;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_85 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_85 <= _GEN_8330;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_86 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_86 <= _GEN_8331;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_87 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_87 <= _GEN_8332;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_88 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_88 <= _GEN_8333;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_89 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_89 <= _GEN_8334;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_90 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_90 <= _GEN_8335;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_91 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_91 <= _GEN_8336;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_92 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_92 <= _GEN_8337;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_93 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_93 <= _GEN_8338;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_94 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_94 <= _GEN_8339;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_95 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_95 <= _GEN_8340;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_96 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_96 <= _GEN_8341;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_97 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_97 <= _GEN_8342;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_98 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_98 <= _GEN_8343;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_99 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_99 <= _GEN_8344;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_100 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_100 <= _GEN_8345;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_101 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_101 <= _GEN_8346;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_102 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_102 <= _GEN_8347;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_103 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_103 <= _GEN_8348;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_104 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_104 <= _GEN_8349;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_105 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_105 <= _GEN_8350;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_106 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_106 <= _GEN_8351;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_107 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_107 <= _GEN_8352;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_108 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_108 <= _GEN_8353;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_109 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_109 <= _GEN_8354;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_110 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_110 <= _GEN_8355;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_111 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_111 <= _GEN_8356;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_112 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_112 <= _GEN_8357;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_113 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_113 <= _GEN_8358;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_114 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_114 <= _GEN_8359;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_115 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_115 <= _GEN_8360;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_116 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_116 <= _GEN_8361;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_117 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_117 <= _GEN_8362;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_118 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_118 <= _GEN_8363;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_119 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_119 <= _GEN_8364;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_120 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_120 <= _GEN_8365;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_121 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_121 <= _GEN_8366;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_122 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_122 <= _GEN_8367;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_123 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_123 <= _GEN_8368;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_124 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_124 <= _GEN_8369;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_125 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_125 <= _GEN_8370;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_126 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_126 <= _GEN_8371;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_127 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_127 <= _GEN_8372;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_128 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_128 <= _GEN_8373;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_129 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_129 <= _GEN_8374;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_130 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_130 <= _GEN_8375;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_131 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_131 <= _GEN_8376;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_132 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_132 <= _GEN_8377;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_133 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_133 <= _GEN_8378;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_134 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_134 <= _GEN_8379;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_135 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_135 <= _GEN_8380;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_136 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_136 <= _GEN_8381;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_137 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_137 <= _GEN_8382;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_138 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_138 <= _GEN_8383;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_139 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_139 <= _GEN_8384;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_140 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_140 <= _GEN_8385;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_141 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_141 <= _GEN_8386;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_142 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_142 <= _GEN_8387;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_143 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_143 <= _GEN_8388;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_144 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_144 <= _GEN_8389;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_145 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_145 <= _GEN_8390;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_146 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_146 <= _GEN_8391;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_147 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_147 <= _GEN_8392;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_148 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_148 <= _GEN_8393;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_149 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_149 <= _GEN_8394;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_150 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_150 <= _GEN_8395;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_151 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_151 <= _GEN_8396;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_152 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_152 <= _GEN_8397;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_153 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_153 <= _GEN_8398;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_154 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_154 <= _GEN_8399;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_155 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_155 <= _GEN_8400;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_156 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_156 <= _GEN_8401;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_157 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_157 <= _GEN_8402;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_158 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_158 <= _GEN_8403;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_159 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_159 <= _GEN_8404;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_160 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_160 <= _GEN_8405;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_161 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_161 <= _GEN_8406;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_162 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_162 <= _GEN_8407;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_163 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_163 <= _GEN_8408;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_164 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_164 <= _GEN_8409;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_165 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_165 <= _GEN_8410;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_166 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_166 <= _GEN_8411;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_167 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_167 <= _GEN_8412;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_168 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_168 <= _GEN_8413;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_169 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_169 <= _GEN_8414;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_170 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_170 <= _GEN_8415;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_171 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_171 <= _GEN_8416;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_172 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_172 <= _GEN_8417;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_173 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_173 <= _GEN_8418;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_174 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_174 <= _GEN_8419;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_175 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_175 <= _GEN_8420;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_176 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_176 <= _GEN_8421;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_177 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_177 <= _GEN_8422;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_178 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_178 <= _GEN_8423;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_179 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_179 <= _GEN_8424;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_180 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_180 <= _GEN_8425;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_181 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_181 <= _GEN_8426;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_182 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_182 <= _GEN_8427;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_183 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_183 <= _GEN_8428;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_184 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_184 <= _GEN_8429;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_185 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_185 <= _GEN_8430;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_186 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_186 <= _GEN_8431;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_187 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_187 <= _GEN_8432;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_188 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_188 <= _GEN_8433;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_189 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_189 <= _GEN_8434;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_190 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_190 <= _GEN_8435;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_191 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_191 <= _GEN_8436;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_192 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_192 <= _GEN_8437;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_193 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_193 <= _GEN_8438;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_194 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_194 <= _GEN_8439;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_195 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_195 <= _GEN_8440;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_196 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_196 <= _GEN_8441;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_197 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_197 <= _GEN_8442;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_198 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_198 <= _GEN_8443;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_199 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_199 <= _GEN_8444;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_200 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_200 <= _GEN_8445;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_201 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_201 <= _GEN_8446;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_202 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_202 <= _GEN_8447;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_203 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_203 <= _GEN_8448;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_204 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_204 <= _GEN_8449;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_205 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_205 <= _GEN_8450;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_206 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_206 <= _GEN_8451;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_207 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_207 <= _GEN_8452;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_208 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_208 <= _GEN_8453;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_209 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_209 <= _GEN_8454;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_210 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_210 <= _GEN_8455;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_211 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_211 <= _GEN_8456;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_212 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_212 <= _GEN_8457;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_213 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_213 <= _GEN_8458;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_214 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_214 <= _GEN_8459;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_215 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_215 <= _GEN_8460;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_216 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_216 <= _GEN_8461;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_217 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_217 <= _GEN_8462;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_218 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_218 <= _GEN_8463;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_219 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_219 <= _GEN_8464;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_220 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_220 <= _GEN_8465;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_221 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_221 <= _GEN_8466;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_222 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_222 <= _GEN_8467;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_223 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_223 <= _GEN_8468;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_224 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_224 <= _GEN_8469;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_225 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_225 <= _GEN_8470;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_226 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_226 <= _GEN_8471;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_227 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_227 <= _GEN_8472;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_228 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_228 <= _GEN_8473;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_229 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_229 <= _GEN_8474;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_230 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_230 <= _GEN_8475;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_231 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_231 <= _GEN_8476;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_232 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_232 <= _GEN_8477;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_233 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_233 <= _GEN_8478;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_234 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_234 <= _GEN_8479;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_235 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_235 <= _GEN_8480;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_236 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_236 <= _GEN_8481;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_237 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_237 <= _GEN_8482;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_238 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_238 <= _GEN_8483;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_239 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_239 <= _GEN_8484;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_240 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_240 <= _GEN_8485;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_241 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_241 <= _GEN_8486;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_242 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_242 <= _GEN_8487;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_243 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_243 <= _GEN_8488;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_244 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_244 <= _GEN_8489;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_245 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_245 <= _GEN_8490;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_246 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_246 <= _GEN_8491;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_247 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_247 <= _GEN_8492;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_248 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_248 <= _GEN_8493;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_249 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_249 <= _GEN_8494;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_250 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_250 <= _GEN_8495;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_251 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_251 <= _GEN_8496;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_252 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_252 <= _GEN_8497;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_253 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_253 <= _GEN_8498;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_254 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_254 <= _GEN_8499;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_255 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_255 <= _GEN_8500;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_256 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_256 <= _GEN_8501;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_257 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_257 <= _GEN_8502;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_258 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_258 <= _GEN_8503;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_259 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_259 <= _GEN_8504;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_260 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_260 <= _GEN_8505;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_261 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_261 <= _GEN_8506;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_262 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_262 <= _GEN_8507;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_263 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_263 <= _GEN_8508;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_264 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_264 <= _GEN_8509;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_265 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_265 <= _GEN_8510;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_266 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_266 <= _GEN_8511;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_267 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_267 <= _GEN_8512;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_268 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_268 <= _GEN_8513;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_269 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_269 <= _GEN_8514;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_270 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_270 <= _GEN_8515;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_271 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_271 <= _GEN_8516;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_272 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_272 <= _GEN_8517;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_273 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_273 <= _GEN_8518;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_274 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_274 <= _GEN_8519;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_275 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_275 <= _GEN_8520;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_276 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_276 <= _GEN_8521;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_277 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_277 <= _GEN_8522;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_278 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_278 <= _GEN_8523;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_279 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_279 <= _GEN_8524;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_280 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_280 <= _GEN_8525;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_281 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_281 <= _GEN_8526;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_282 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_282 <= _GEN_8527;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_283 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_283 <= _GEN_8528;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_284 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_284 <= _GEN_8529;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_285 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_285 <= _GEN_8530;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_286 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_286 <= _GEN_8531;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_287 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_287 <= _GEN_8532;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_288 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_288 <= _GEN_8533;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_289 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_289 <= _GEN_8534;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_290 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_290 <= _GEN_8535;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_291 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_291 <= _GEN_8536;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_292 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_292 <= _GEN_8537;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_293 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_293 <= _GEN_8538;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_294 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_294 <= _GEN_8539;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_295 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_295 <= _GEN_8540;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_296 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_296 <= _GEN_8541;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_297 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_297 <= _GEN_8542;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_298 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_298 <= _GEN_8543;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_299 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_299 <= _GEN_8544;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_300 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_300 <= _GEN_8545;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_301 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_301 <= _GEN_8546;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_302 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_302 <= _GEN_8547;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_303 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_303 <= _GEN_8548;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_304 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_304 <= _GEN_8549;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_305 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_305 <= _GEN_8550;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_306 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_306 <= _GEN_8551;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_307 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_307 <= _GEN_8552;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_308 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_308 <= _GEN_8553;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_309 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_309 <= _GEN_8554;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_310 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_310 <= _GEN_8555;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_311 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_311 <= _GEN_8556;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_312 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_312 <= _GEN_8557;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_313 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_313 <= _GEN_8558;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_314 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_314 <= _GEN_8559;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_315 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_315 <= _GEN_8560;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_316 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_316 <= _GEN_8561;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_317 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_317 <= _GEN_8562;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_318 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_318 <= _GEN_8563;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_319 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_319 <= _GEN_8564;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_320 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_320 <= _GEN_8565;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_321 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_321 <= _GEN_8566;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_322 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_322 <= _GEN_8567;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_323 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_323 <= _GEN_8568;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_324 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_324 <= _GEN_8569;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_325 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_325 <= _GEN_8570;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_326 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_326 <= _GEN_8571;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_327 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_327 <= _GEN_8572;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_328 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_328 <= _GEN_8573;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_329 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_329 <= _GEN_8574;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_330 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_330 <= _GEN_8575;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_331 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_331 <= _GEN_8576;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_332 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_332 <= _GEN_8577;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_333 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_333 <= _GEN_8578;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_334 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_334 <= _GEN_8579;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_335 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_335 <= _GEN_8580;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_336 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_336 <= _GEN_8581;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_337 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_337 <= _GEN_8582;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_338 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_338 <= _GEN_8583;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_339 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_339 <= _GEN_8584;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_340 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_340 <= _GEN_8585;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_341 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_341 <= _GEN_8586;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_342 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_342 <= _GEN_8587;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_343 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_343 <= _GEN_8588;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_344 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_344 <= _GEN_8589;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_345 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_345 <= _GEN_8590;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_346 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_346 <= _GEN_8591;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_347 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_347 <= _GEN_8592;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_348 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_348 <= _GEN_8593;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_349 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_349 <= _GEN_8594;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_350 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_350 <= _GEN_8595;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_351 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_351 <= _GEN_8596;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_352 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_352 <= _GEN_8597;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_353 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_353 <= _GEN_8598;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_354 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_354 <= _GEN_8599;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_355 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_355 <= _GEN_8600;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_356 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_356 <= _GEN_8601;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_357 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_357 <= _GEN_8602;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_358 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_358 <= _GEN_8603;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_359 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_359 <= _GEN_8604;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_360 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_360 <= _GEN_8605;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_361 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_361 <= _GEN_8606;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_362 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_362 <= _GEN_8607;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_363 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_363 <= _GEN_8608;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_364 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_364 <= _GEN_8609;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_365 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_365 <= _GEN_8610;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_366 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_366 <= _GEN_8611;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_367 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_367 <= _GEN_8612;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_368 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_368 <= _GEN_8613;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_369 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_369 <= _GEN_8614;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_370 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_370 <= _GEN_8615;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_371 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_371 <= _GEN_8616;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_372 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_372 <= _GEN_8617;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_373 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_373 <= _GEN_8618;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_374 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_374 <= _GEN_8619;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_375 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_375 <= _GEN_8620;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_376 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_376 <= _GEN_8621;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_377 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_377 <= _GEN_8622;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_378 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_378 <= _GEN_8623;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_379 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_379 <= _GEN_8624;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_380 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_380 <= _GEN_8625;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_381 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_381 <= _GEN_8626;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_382 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_382 <= _GEN_8627;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_383 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_383 <= _GEN_8628;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_384 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_384 <= _GEN_8629;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_385 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_385 <= _GEN_8630;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_386 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_386 <= _GEN_8631;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_387 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_387 <= _GEN_8632;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_388 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_388 <= _GEN_8633;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_389 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_389 <= _GEN_8634;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_390 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_390 <= _GEN_8635;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_391 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_391 <= _GEN_8636;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_392 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_392 <= _GEN_8637;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_393 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_393 <= _GEN_8638;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_394 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_394 <= _GEN_8639;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_395 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_395 <= _GEN_8640;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_396 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_396 <= _GEN_8641;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_397 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_397 <= _GEN_8642;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_398 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_398 <= _GEN_8643;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_399 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_399 <= _GEN_8644;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_400 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_400 <= _GEN_8645;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_401 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_401 <= _GEN_8646;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_402 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_402 <= _GEN_8647;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_403 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_403 <= _GEN_8648;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_404 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_404 <= _GEN_8649;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_405 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_405 <= _GEN_8650;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_406 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_406 <= _GEN_8651;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_407 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_407 <= _GEN_8652;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_408 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_408 <= _GEN_8653;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_409 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_409 <= _GEN_8654;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_410 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_410 <= _GEN_8655;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_411 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_411 <= _GEN_8656;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_412 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_412 <= _GEN_8657;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_413 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_413 <= _GEN_8658;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_414 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_414 <= _GEN_8659;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_415 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_415 <= _GEN_8660;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_416 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_416 <= _GEN_8661;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_417 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_417 <= _GEN_8662;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_418 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_418 <= _GEN_8663;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_419 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_419 <= _GEN_8664;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_420 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_420 <= _GEN_8665;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_421 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_421 <= _GEN_8666;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_422 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_422 <= _GEN_8667;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_423 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_423 <= _GEN_8668;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_424 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_424 <= _GEN_8669;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_425 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_425 <= _GEN_8670;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_426 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_426 <= _GEN_8671;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_427 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_427 <= _GEN_8672;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_428 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_428 <= _GEN_8673;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_429 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_429 <= _GEN_8674;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_430 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_430 <= _GEN_8675;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_431 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_431 <= _GEN_8676;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_432 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_432 <= _GEN_8677;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_433 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_433 <= _GEN_8678;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_434 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_434 <= _GEN_8679;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_435 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_435 <= _GEN_8680;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_436 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_436 <= _GEN_8681;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_437 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_437 <= _GEN_8682;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_438 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_438 <= _GEN_8683;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_439 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_439 <= _GEN_8684;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_440 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_440 <= _GEN_8685;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_441 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_441 <= _GEN_8686;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_442 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_442 <= _GEN_8687;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_443 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_443 <= _GEN_8688;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_444 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_444 <= _GEN_8689;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_445 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_445 <= _GEN_8690;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_446 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_446 <= _GEN_8691;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_447 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_447 <= _GEN_8692;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_448 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_448 <= _GEN_8693;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_449 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_449 <= _GEN_8694;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_450 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_450 <= _GEN_8695;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_451 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_451 <= _GEN_8696;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_452 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_452 <= _GEN_8697;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_453 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_453 <= _GEN_8698;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_454 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_454 <= _GEN_8699;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_455 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_455 <= _GEN_8700;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_456 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_456 <= _GEN_8701;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_457 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_457 <= _GEN_8702;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_458 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_458 <= _GEN_8703;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_459 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_459 <= _GEN_8704;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_460 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_460 <= _GEN_8705;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_461 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_461 <= _GEN_8706;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_462 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_462 <= _GEN_8707;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_463 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_463 <= _GEN_8708;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_464 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_464 <= _GEN_8709;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_465 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_465 <= _GEN_8710;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_466 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_466 <= _GEN_8711;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_467 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_467 <= _GEN_8712;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_468 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_468 <= _GEN_8713;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_469 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_469 <= _GEN_8714;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_470 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_470 <= _GEN_8715;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_471 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_471 <= _GEN_8716;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_472 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_472 <= _GEN_8717;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_473 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_473 <= _GEN_8718;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_474 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_474 <= _GEN_8719;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_475 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_475 <= _GEN_8720;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_476 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_476 <= _GEN_8721;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_477 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_477 <= _GEN_8722;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_478 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_478 <= _GEN_8723;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_479 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_479 <= _GEN_8724;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_480 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_480 <= _GEN_8725;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_481 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_481 <= _GEN_8726;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_482 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_482 <= _GEN_8727;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_483 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_483 <= _GEN_8728;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_484 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_484 <= _GEN_8729;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_485 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_485 <= _GEN_8730;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_486 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_486 <= _GEN_8731;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_487 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_487 <= _GEN_8732;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_488 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_488 <= _GEN_8733;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_489 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_489 <= _GEN_8734;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_490 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_490 <= _GEN_8735;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_491 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_491 <= _GEN_8736;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_492 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_492 <= _GEN_8737;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_493 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_493 <= _GEN_8738;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_494 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_494 <= _GEN_8739;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_495 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_495 <= _GEN_8740;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_496 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_496 <= _GEN_8741;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_497 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_497 <= _GEN_8742;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_498 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_498 <= _GEN_8743;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_499 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_499 <= _GEN_8744;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_500 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_500 <= _GEN_8745;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_501 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_501 <= _GEN_8746;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_502 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_502 <= _GEN_8747;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_503 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_503 <= _GEN_8748;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_504 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_504 <= _GEN_8749;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_505 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_505 <= _GEN_8750;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_506 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_506 <= _GEN_8751;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_507 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_507 <= _GEN_8752;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_508 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_508 <= _GEN_8753;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_509 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_509 <= _GEN_8754;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_510 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_510 <= _GEN_8755;
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:20]
      lru_511 <= 1'h0; // @[ICache.scala 68:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          lru_511 <= _GEN_8756;
        end
      end
    end
    if (reset) begin // @[ICache.scala 71:20]
      tlb_vpn <= 20'h0; // @[ICache.scala 71:20]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 164:17]
      if (3'h1 == state) begin // @[ICache.scala 164:17]
        if (io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_v_1 | ~inst_vpn[12] & io_cpu_tlb2_entry_v_0)) begin // @[ICache.scala 201:118]
          tlb_vpn <= {{1'd0}, io_cpu_tlb2_vpn}; // @[ICache.scala 203:22]
        end
      end
    end
    if (reset) begin // @[ICache.scala 71:20]
      tlb_ppn <= 20'h0; // @[ICache.scala 71:20]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 164:17]
      if (3'h1 == state) begin // @[ICache.scala 164:17]
        if (io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_v_1 | ~inst_vpn[12] & io_cpu_tlb2_entry_v_0)) begin // @[ICache.scala 201:118]
          tlb_ppn <= _GEN_11867; // @[ICache.scala 204:22]
        end
      end
    end
    if (reset) begin // @[ICache.scala 71:20]
      tlb_uncached <= 1'h0; // @[ICache.scala 71:20]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 164:17]
      if (3'h1 == state) begin // @[ICache.scala 164:17]
        if (io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_v_1 | ~inst_vpn[12] & io_cpu_tlb2_entry_v_0)) begin // @[ICache.scala 201:118]
          tlb_uncached <= _GEN_11869; // @[ICache.scala 205:22]
        end
      end
    end
    if (reset) begin // @[ICache.scala 71:20]
      tlb_valid <= 1'h0; // @[ICache.scala 71:20]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      tlb_valid <= _GEN_2;
    end else if (3'h1 == state) begin // @[ICache.scala 164:17]
      tlb_valid <= _GEN_11874;
    end else begin
      tlb_valid <= _GEN_2;
    end
    if (reset) begin // @[ICache.scala 95:21]
      rset <= 6'h0; // @[ICache.scala 95:21]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          rset <= _GEN_7212;
        end
      end
    end
    if (reset) begin // @[ICache.scala 113:22]
      saved_0_inst <= 32'h0; // @[ICache.scala 113:22]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 164:17]
      if (3'h1 == state) begin // @[ICache.scala 164:17]
        if (!(io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_v_1 | ~inst_vpn[12] & io_cpu_tlb2_entry_v_0))) begin // @[ICache.scala 201:118]
          saved_0_inst <= 32'h0; // @[ICache.scala 210:24]
        end
      end else if (3'h2 == state) begin // @[ICache.scala 164:17]
        saved_0_inst <= _GEN_11887;
      end
    end
    if (reset) begin // @[ICache.scala 113:22]
      saved_0_valid <= 1'h0; // @[ICache.scala 113:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          saved_0_valid <= _GEN_8758;
        end
      end
    end else if (3'h1 == state) begin // @[ICache.scala 164:17]
      if (!(io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_v_1 | ~inst_vpn[12] & io_cpu_tlb2_entry_v_0))) begin // @[ICache.scala 201:118]
        saved_0_valid <= 1'h1; // @[ICache.scala 211:24]
      end
    end else if (3'h2 == state) begin // @[ICache.scala 164:17]
      saved_0_valid <= _GEN_11888;
    end else begin
      saved_0_valid <= _GEN_11949;
    end
    if (reset) begin // @[ICache.scala 113:22]
      saved_1_inst <= 32'h0; // @[ICache.scala 113:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          saved_1_inst <= _GEN_8757;
        end
      end
    end
    if (reset) begin // @[ICache.scala 113:22]
      saved_1_valid <= 1'h0; // @[ICache.scala 113:22]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          saved_1_valid <= _GEN_8759;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        saved_1_valid <= _GEN_11950;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      axi_cnt_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          axi_cnt_value <= _GEN_8244;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        axi_cnt_value <= _GEN_11940;
      end
    end
    if (reset) begin // @[ICache.scala 149:24]
      ar_addr <= 32'h0; // @[ICache.scala 149:24]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          ar_addr <= _GEN_7208;
        end
      end
    end
    if (reset) begin // @[ICache.scala 149:24]
      ar_len <= 8'h0; // @[ICache.scala 149:24]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          ar_len <= _GEN_7209;
        end
      end
    end
    if (reset) begin // @[ICache.scala 149:24]
      ar_size <= 3'h0; // @[ICache.scala 149:24]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          ar_size <= _GEN_7210;
        end
      end
    end
    if (reset) begin // @[ICache.scala 150:24]
      arvalid <= 1'h0; // @[ICache.scala 150:24]
    end else if (3'h0 == state) begin // @[ICache.scala 164:17]
      if (io_cpu_req) begin // @[ICache.scala 166:24]
        if (!(_io_cpu_tlb2_vpn_T_2)) begin // @[ICache.scala 167:31]
          arvalid <= _GEN_7211;
        end
      end
    end else if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
      if (3'h2 == state) begin // @[ICache.scala 164:17]
        arvalid <= _GEN_11884;
      end else begin
        arvalid <= _GEN_11938;
      end
    end
    if (reset) begin // @[ICache.scala 155:23]
      rready <= 1'h0; // @[ICache.scala 155:23]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 164:17]
      if (!(3'h1 == state)) begin // @[ICache.scala 164:17]
        if (3'h2 == state) begin // @[ICache.scala 164:17]
          rready <= _GEN_11885;
        end else begin
          rready <= _GEN_11939;
        end
      end
    end
    if (reset) begin // @[ICache.scala 159:29]
      tlb1_invalid <= 1'h0; // @[ICache.scala 159:29]
    end else if (!(3'h0 == state)) begin // @[ICache.scala 164:17]
      if (3'h1 == state) begin // @[ICache.scala 164:17]
        if (!(io_cpu_tlb2_found & (inst_vpn[12] & io_cpu_tlb2_entry_v_1 | ~inst_vpn[12] & io_cpu_tlb2_entry_v_0))) begin // @[ICache.scala 201:118]
          tlb1_invalid <= 1'h1; // @[ICache.scala 209:24]
        end
      end else if (!(3'h2 == state)) begin // @[ICache.scala 164:17]
        tlb1_invalid <= _GEN_11948;
      end
    end
    if (_io_cpu_tlb2_vpn_T_3) begin // @[Reg.scala 20:18]
      io_cpu_tlb2_vpn_r <= inst_vpn; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  valid_0_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  valid_0_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_1_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_1_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_2_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_2_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_3_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_3_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_4_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_4_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_5_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_5_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_6_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_6_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_7_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_7_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_8_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_8_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_9_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_9_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_10_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_10_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_11_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_11_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_12_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_12_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_13_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_13_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_14_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_14_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_15_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_15_1 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_16_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_16_1 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_17_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_17_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_18_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_18_1 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_19_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_19_1 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_20_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_20_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_21_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_21_1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_22_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_22_1 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_23_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_23_1 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_24_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_24_1 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_25_0 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_25_1 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_26_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_26_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_27_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_27_1 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_28_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_28_1 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_29_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_29_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_30_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_30_1 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_31_0 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_31_1 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_32_0 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_32_1 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_33_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_33_1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_34_0 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_34_1 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_35_0 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_35_1 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_36_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_36_1 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_37_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_37_1 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_38_0 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_38_1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_39_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_39_1 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_40_0 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_40_1 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_41_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_41_1 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_42_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_42_1 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_43_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_43_1 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_44_0 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_44_1 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_45_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_45_1 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_46_0 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_46_1 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_47_0 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_47_1 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_48_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_48_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_49_0 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_49_1 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_50_0 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_50_1 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_51_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_51_1 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_52_0 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_52_1 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_53_0 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_53_1 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_54_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_54_1 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_55_0 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_55_1 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_56_0 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_56_1 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_57_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_57_1 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_58_0 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_58_1 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_59_0 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_59_1 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_60_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_60_1 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_61_0 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_61_1 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_62_0 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_62_1 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_63_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_63_1 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_64_0 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_64_1 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_65_0 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_65_1 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_66_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_66_1 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_67_0 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_67_1 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_68_0 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_68_1 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_69_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_69_1 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_70_0 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_70_1 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_71_0 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_71_1 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_72_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_72_1 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_73_0 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_73_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_74_0 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_74_1 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_75_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_75_1 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_76_0 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_76_1 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_77_0 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_77_1 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_78_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_78_1 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_79_0 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_79_1 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_80_0 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_80_1 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_81_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_81_1 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_82_0 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_82_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_83_0 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_83_1 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_84_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_84_1 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_85_0 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_85_1 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_86_0 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_86_1 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_87_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_87_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_88_0 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_88_1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_89_0 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_89_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_90_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_90_1 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_91_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_91_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_92_0 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_92_1 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_93_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_93_1 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_94_0 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_94_1 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_95_0 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_95_1 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_96_0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_96_1 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_97_0 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_97_1 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_98_0 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_98_1 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_99_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_99_1 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_100_0 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_100_1 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_101_0 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_101_1 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_102_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_102_1 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_103_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_103_1 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_104_0 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_104_1 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_105_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_105_1 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_106_0 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_106_1 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_107_0 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_107_1 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_108_0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_108_1 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_109_0 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_109_1 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_110_0 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_110_1 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_111_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_111_1 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_112_0 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_112_1 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_113_0 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_113_1 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_114_0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_114_1 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_115_0 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_115_1 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_116_0 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_116_1 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_117_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_117_1 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_118_0 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_118_1 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_119_0 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_119_1 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_120_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_120_1 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_121_0 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_121_1 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_122_0 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_122_1 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_123_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_123_1 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_124_0 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_124_1 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_125_0 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_125_1 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_126_0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_126_1 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_127_0 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_127_1 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_128_0 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_128_1 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_129_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_129_1 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_130_0 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_130_1 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_131_0 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_131_1 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_132_0 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_132_1 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_133_0 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_133_1 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_134_0 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_134_1 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_135_0 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_135_1 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_136_0 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_136_1 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_137_0 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_137_1 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_138_0 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_138_1 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_139_0 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_139_1 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_140_0 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_140_1 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_141_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_141_1 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_142_0 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_142_1 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_143_0 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_143_1 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_144_0 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_144_1 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_145_0 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_145_1 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_146_0 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_146_1 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_147_0 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_147_1 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_148_0 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_148_1 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_149_0 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_149_1 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_150_0 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_150_1 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_151_0 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_151_1 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_152_0 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_152_1 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_153_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_153_1 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_154_0 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_154_1 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_155_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_155_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_156_0 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_156_1 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_157_0 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_157_1 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_158_0 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_158_1 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_159_0 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_159_1 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_160_0 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_160_1 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_161_0 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_161_1 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_162_0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_162_1 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_163_0 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_163_1 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_164_0 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_164_1 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_165_0 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_165_1 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_166_0 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_166_1 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_167_0 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_167_1 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_168_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_168_1 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_169_0 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_169_1 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_170_0 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_170_1 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_171_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_171_1 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_172_0 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_172_1 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_173_0 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_173_1 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_174_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_174_1 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_175_0 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_175_1 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_176_0 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_176_1 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_177_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_177_1 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_178_0 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_178_1 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_179_0 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_179_1 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_180_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_180_1 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_181_0 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_181_1 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_182_0 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_182_1 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_183_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_183_1 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_184_0 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_184_1 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_185_0 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_185_1 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_186_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_186_1 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_187_0 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_187_1 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_188_0 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_188_1 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_189_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_189_1 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_190_0 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_190_1 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_191_0 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_191_1 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_192_0 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_192_1 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_193_0 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_193_1 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_194_0 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_194_1 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_195_0 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_195_1 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_196_0 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_196_1 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_197_0 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_197_1 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_198_0 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_198_1 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_199_0 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_199_1 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_200_0 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_200_1 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_201_0 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_201_1 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_202_0 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_202_1 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_203_0 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_203_1 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_204_0 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_204_1 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_205_0 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_205_1 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_206_0 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_206_1 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_207_0 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_207_1 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_208_0 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_208_1 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_209_0 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_209_1 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_210_0 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_210_1 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_211_0 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_211_1 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_212_0 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_212_1 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_213_0 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_213_1 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_214_0 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_214_1 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_215_0 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_215_1 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_216_0 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_216_1 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_217_0 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_217_1 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_218_0 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_218_1 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_219_0 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_219_1 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_220_0 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_220_1 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_221_0 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_221_1 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_222_0 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_222_1 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_223_0 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_223_1 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_224_0 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_224_1 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_225_0 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_225_1 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_226_0 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_226_1 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_227_0 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_227_1 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_228_0 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_228_1 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_229_0 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_229_1 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_230_0 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_230_1 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_231_0 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_231_1 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_232_0 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_232_1 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_233_0 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_233_1 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_234_0 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_234_1 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_235_0 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_235_1 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_236_0 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_236_1 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_237_0 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_237_1 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_238_0 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_238_1 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_239_0 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_239_1 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_240_0 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_240_1 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_241_0 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_241_1 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_242_0 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_242_1 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_243_0 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_243_1 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_244_0 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_244_1 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_245_0 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_245_1 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_246_0 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_246_1 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_247_0 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_247_1 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_248_0 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_248_1 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_249_0 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_249_1 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_250_0 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_250_1 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_251_0 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_251_1 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_252_0 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_252_1 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_253_0 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_253_1 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_254_0 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_254_1 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_255_0 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  valid_255_1 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_256_0 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_256_1 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_257_0 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_257_1 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_258_0 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_258_1 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_259_0 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_259_1 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_260_0 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_260_1 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_261_0 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_261_1 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_262_0 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_262_1 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_263_0 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_263_1 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_264_0 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_264_1 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_265_0 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_265_1 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_266_0 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_266_1 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_267_0 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_267_1 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_268_0 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_268_1 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_269_0 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_269_1 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_270_0 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_270_1 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_271_0 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_271_1 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_272_0 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_272_1 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_273_0 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_273_1 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_274_0 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_274_1 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_275_0 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_275_1 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_276_0 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_276_1 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_277_0 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_277_1 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_278_0 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_278_1 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_279_0 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_279_1 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_280_0 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_280_1 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_281_0 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_281_1 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_282_0 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_282_1 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_283_0 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_283_1 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_284_0 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_284_1 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_285_0 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_285_1 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_286_0 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_286_1 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_287_0 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_287_1 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_288_0 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_288_1 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_289_0 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_289_1 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_290_0 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_290_1 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_291_0 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_291_1 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_292_0 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_292_1 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_293_0 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_293_1 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_294_0 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_294_1 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_295_0 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_295_1 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_296_0 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_296_1 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_297_0 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_297_1 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_298_0 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_298_1 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_299_0 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_299_1 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_300_0 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_300_1 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_301_0 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_301_1 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_302_0 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_302_1 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_303_0 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_303_1 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_304_0 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_304_1 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_305_0 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_305_1 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_306_0 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_306_1 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_307_0 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_307_1 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_308_0 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_308_1 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_309_0 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_309_1 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_310_0 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_310_1 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_311_0 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_311_1 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_312_0 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_312_1 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_313_0 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_313_1 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_314_0 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_314_1 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_315_0 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_315_1 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_316_0 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_316_1 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_317_0 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_317_1 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_318_0 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_318_1 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_319_0 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_319_1 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_320_0 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_320_1 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_321_0 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_321_1 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_322_0 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_322_1 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_323_0 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_323_1 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_324_0 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_324_1 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_325_0 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_325_1 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_326_0 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_326_1 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_327_0 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_327_1 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_328_0 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_328_1 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_329_0 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_329_1 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_330_0 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_330_1 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_331_0 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_331_1 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_332_0 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_332_1 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_333_0 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_333_1 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_334_0 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_334_1 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_335_0 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_335_1 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_336_0 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_336_1 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_337_0 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_337_1 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_338_0 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_338_1 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_339_0 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_339_1 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_340_0 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_340_1 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_341_0 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_341_1 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_342_0 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_342_1 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_343_0 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_343_1 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_344_0 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_344_1 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_345_0 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_345_1 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_346_0 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_346_1 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_347_0 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_347_1 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_348_0 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_348_1 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_349_0 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_349_1 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_350_0 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_350_1 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_351_0 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_351_1 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_352_0 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_352_1 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_353_0 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_353_1 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_354_0 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_354_1 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_355_0 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_355_1 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_356_0 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_356_1 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_357_0 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_357_1 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_358_0 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_358_1 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_359_0 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_359_1 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_360_0 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_360_1 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_361_0 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_361_1 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_362_0 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_362_1 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_363_0 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_363_1 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_364_0 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_364_1 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_365_0 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_365_1 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_366_0 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_366_1 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_367_0 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_367_1 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_368_0 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_368_1 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_369_0 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_369_1 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_370_0 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_370_1 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_371_0 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_371_1 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_372_0 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_372_1 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_373_0 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_373_1 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_374_0 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_374_1 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_375_0 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_375_1 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_376_0 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_376_1 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_377_0 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_377_1 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_378_0 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_378_1 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_379_0 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_379_1 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_380_0 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_380_1 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_381_0 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_381_1 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_382_0 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_382_1 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_383_0 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  valid_383_1 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  valid_384_0 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  valid_384_1 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  valid_385_0 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  valid_385_1 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  valid_386_0 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  valid_386_1 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  valid_387_0 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  valid_387_1 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  valid_388_0 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  valid_388_1 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  valid_389_0 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  valid_389_1 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  valid_390_0 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  valid_390_1 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  valid_391_0 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  valid_391_1 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  valid_392_0 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  valid_392_1 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  valid_393_0 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  valid_393_1 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  valid_394_0 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  valid_394_1 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  valid_395_0 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  valid_395_1 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  valid_396_0 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  valid_396_1 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  valid_397_0 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  valid_397_1 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  valid_398_0 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  valid_398_1 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  valid_399_0 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  valid_399_1 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  valid_400_0 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  valid_400_1 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  valid_401_0 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  valid_401_1 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  valid_402_0 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  valid_402_1 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  valid_403_0 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  valid_403_1 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  valid_404_0 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  valid_404_1 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  valid_405_0 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  valid_405_1 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  valid_406_0 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  valid_406_1 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  valid_407_0 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  valid_407_1 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  valid_408_0 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  valid_408_1 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  valid_409_0 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  valid_409_1 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  valid_410_0 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  valid_410_1 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  valid_411_0 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  valid_411_1 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  valid_412_0 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  valid_412_1 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  valid_413_0 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  valid_413_1 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  valid_414_0 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  valid_414_1 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  valid_415_0 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  valid_415_1 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  valid_416_0 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  valid_416_1 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  valid_417_0 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  valid_417_1 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  valid_418_0 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  valid_418_1 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  valid_419_0 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  valid_419_1 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  valid_420_0 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  valid_420_1 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  valid_421_0 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  valid_421_1 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  valid_422_0 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  valid_422_1 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  valid_423_0 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  valid_423_1 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  valid_424_0 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  valid_424_1 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  valid_425_0 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  valid_425_1 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  valid_426_0 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  valid_426_1 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  valid_427_0 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  valid_427_1 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  valid_428_0 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  valid_428_1 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  valid_429_0 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  valid_429_1 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  valid_430_0 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  valid_430_1 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  valid_431_0 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  valid_431_1 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  valid_432_0 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  valid_432_1 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  valid_433_0 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  valid_433_1 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  valid_434_0 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  valid_434_1 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  valid_435_0 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  valid_435_1 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  valid_436_0 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  valid_436_1 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  valid_437_0 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  valid_437_1 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  valid_438_0 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  valid_438_1 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  valid_439_0 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  valid_439_1 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  valid_440_0 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  valid_440_1 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  valid_441_0 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  valid_441_1 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  valid_442_0 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  valid_442_1 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  valid_443_0 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  valid_443_1 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  valid_444_0 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  valid_444_1 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  valid_445_0 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  valid_445_1 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  valid_446_0 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  valid_446_1 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  valid_447_0 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  valid_447_1 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  valid_448_0 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  valid_448_1 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  valid_449_0 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  valid_449_1 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  valid_450_0 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  valid_450_1 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  valid_451_0 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  valid_451_1 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  valid_452_0 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  valid_452_1 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  valid_453_0 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  valid_453_1 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  valid_454_0 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  valid_454_1 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  valid_455_0 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  valid_455_1 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  valid_456_0 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  valid_456_1 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  valid_457_0 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  valid_457_1 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  valid_458_0 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  valid_458_1 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  valid_459_0 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  valid_459_1 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  valid_460_0 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  valid_460_1 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  valid_461_0 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  valid_461_1 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  valid_462_0 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  valid_462_1 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  valid_463_0 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  valid_463_1 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  valid_464_0 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  valid_464_1 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  valid_465_0 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  valid_465_1 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  valid_466_0 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  valid_466_1 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  valid_467_0 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  valid_467_1 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  valid_468_0 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  valid_468_1 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  valid_469_0 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  valid_469_1 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  valid_470_0 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  valid_470_1 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  valid_471_0 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  valid_471_1 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  valid_472_0 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  valid_472_1 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  valid_473_0 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  valid_473_1 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  valid_474_0 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  valid_474_1 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  valid_475_0 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  valid_475_1 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  valid_476_0 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  valid_476_1 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  valid_477_0 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  valid_477_1 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  valid_478_0 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  valid_478_1 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  valid_479_0 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  valid_479_1 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  valid_480_0 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  valid_480_1 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  valid_481_0 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  valid_481_1 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  valid_482_0 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  valid_482_1 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  valid_483_0 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  valid_483_1 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  valid_484_0 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  valid_484_1 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  valid_485_0 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  valid_485_1 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  valid_486_0 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  valid_486_1 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  valid_487_0 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  valid_487_1 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  valid_488_0 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  valid_488_1 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  valid_489_0 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  valid_489_1 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  valid_490_0 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  valid_490_1 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  valid_491_0 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  valid_491_1 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  valid_492_0 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  valid_492_1 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  valid_493_0 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  valid_493_1 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  valid_494_0 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  valid_494_1 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  valid_495_0 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  valid_495_1 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  valid_496_0 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  valid_496_1 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  valid_497_0 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  valid_497_1 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  valid_498_0 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  valid_498_1 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  valid_499_0 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  valid_499_1 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  valid_500_0 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  valid_500_1 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  valid_501_0 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  valid_501_1 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  valid_502_0 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  valid_502_1 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  valid_503_0 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  valid_503_1 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  valid_504_0 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  valid_504_1 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  valid_505_0 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  valid_505_1 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  valid_506_0 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  valid_506_1 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  valid_507_0 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  valid_507_1 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  valid_508_0 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  valid_508_1 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  valid_509_0 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  valid_509_1 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  valid_510_0 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  valid_510_1 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  valid_511_0 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  valid_511_1 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  data_wstrb_0_0 = _RAND_1025[3:0];
  _RAND_1026 = {1{`RANDOM}};
  data_wstrb_0_1 = _RAND_1026[3:0];
  _RAND_1027 = {1{`RANDOM}};
  data_wstrb_1_0 = _RAND_1027[3:0];
  _RAND_1028 = {1{`RANDOM}};
  data_wstrb_1_1 = _RAND_1028[3:0];
  _RAND_1029 = {1{`RANDOM}};
  tag_wstrb_0 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  tag_wstrb_1 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  tag_wdata = _RAND_1031[19:0];
  _RAND_1032 = {1{`RANDOM}};
  lru_0 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  lru_1 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  lru_2 = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  lru_3 = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  lru_4 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  lru_5 = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  lru_6 = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  lru_7 = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  lru_8 = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  lru_9 = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  lru_10 = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  lru_11 = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  lru_12 = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  lru_13 = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  lru_14 = _RAND_1046[0:0];
  _RAND_1047 = {1{`RANDOM}};
  lru_15 = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  lru_16 = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  lru_17 = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  lru_18 = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  lru_19 = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  lru_20 = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  lru_21 = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  lru_22 = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  lru_23 = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  lru_24 = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  lru_25 = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  lru_26 = _RAND_1058[0:0];
  _RAND_1059 = {1{`RANDOM}};
  lru_27 = _RAND_1059[0:0];
  _RAND_1060 = {1{`RANDOM}};
  lru_28 = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  lru_29 = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  lru_30 = _RAND_1062[0:0];
  _RAND_1063 = {1{`RANDOM}};
  lru_31 = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  lru_32 = _RAND_1064[0:0];
  _RAND_1065 = {1{`RANDOM}};
  lru_33 = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  lru_34 = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  lru_35 = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  lru_36 = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  lru_37 = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  lru_38 = _RAND_1070[0:0];
  _RAND_1071 = {1{`RANDOM}};
  lru_39 = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  lru_40 = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  lru_41 = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  lru_42 = _RAND_1074[0:0];
  _RAND_1075 = {1{`RANDOM}};
  lru_43 = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  lru_44 = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  lru_45 = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  lru_46 = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  lru_47 = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  lru_48 = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  lru_49 = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  lru_50 = _RAND_1082[0:0];
  _RAND_1083 = {1{`RANDOM}};
  lru_51 = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  lru_52 = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  lru_53 = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  lru_54 = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  lru_55 = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  lru_56 = _RAND_1088[0:0];
  _RAND_1089 = {1{`RANDOM}};
  lru_57 = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  lru_58 = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  lru_59 = _RAND_1091[0:0];
  _RAND_1092 = {1{`RANDOM}};
  lru_60 = _RAND_1092[0:0];
  _RAND_1093 = {1{`RANDOM}};
  lru_61 = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  lru_62 = _RAND_1094[0:0];
  _RAND_1095 = {1{`RANDOM}};
  lru_63 = _RAND_1095[0:0];
  _RAND_1096 = {1{`RANDOM}};
  lru_64 = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  lru_65 = _RAND_1097[0:0];
  _RAND_1098 = {1{`RANDOM}};
  lru_66 = _RAND_1098[0:0];
  _RAND_1099 = {1{`RANDOM}};
  lru_67 = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  lru_68 = _RAND_1100[0:0];
  _RAND_1101 = {1{`RANDOM}};
  lru_69 = _RAND_1101[0:0];
  _RAND_1102 = {1{`RANDOM}};
  lru_70 = _RAND_1102[0:0];
  _RAND_1103 = {1{`RANDOM}};
  lru_71 = _RAND_1103[0:0];
  _RAND_1104 = {1{`RANDOM}};
  lru_72 = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  lru_73 = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  lru_74 = _RAND_1106[0:0];
  _RAND_1107 = {1{`RANDOM}};
  lru_75 = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  lru_76 = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  lru_77 = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  lru_78 = _RAND_1110[0:0];
  _RAND_1111 = {1{`RANDOM}};
  lru_79 = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  lru_80 = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  lru_81 = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  lru_82 = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  lru_83 = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  lru_84 = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  lru_85 = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  lru_86 = _RAND_1118[0:0];
  _RAND_1119 = {1{`RANDOM}};
  lru_87 = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  lru_88 = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  lru_89 = _RAND_1121[0:0];
  _RAND_1122 = {1{`RANDOM}};
  lru_90 = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  lru_91 = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  lru_92 = _RAND_1124[0:0];
  _RAND_1125 = {1{`RANDOM}};
  lru_93 = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  lru_94 = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  lru_95 = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  lru_96 = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  lru_97 = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  lru_98 = _RAND_1130[0:0];
  _RAND_1131 = {1{`RANDOM}};
  lru_99 = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  lru_100 = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  lru_101 = _RAND_1133[0:0];
  _RAND_1134 = {1{`RANDOM}};
  lru_102 = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  lru_103 = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  lru_104 = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  lru_105 = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  lru_106 = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  lru_107 = _RAND_1139[0:0];
  _RAND_1140 = {1{`RANDOM}};
  lru_108 = _RAND_1140[0:0];
  _RAND_1141 = {1{`RANDOM}};
  lru_109 = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  lru_110 = _RAND_1142[0:0];
  _RAND_1143 = {1{`RANDOM}};
  lru_111 = _RAND_1143[0:0];
  _RAND_1144 = {1{`RANDOM}};
  lru_112 = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  lru_113 = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  lru_114 = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  lru_115 = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  lru_116 = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  lru_117 = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  lru_118 = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  lru_119 = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  lru_120 = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  lru_121 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  lru_122 = _RAND_1154[0:0];
  _RAND_1155 = {1{`RANDOM}};
  lru_123 = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  lru_124 = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  lru_125 = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  lru_126 = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  lru_127 = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  lru_128 = _RAND_1160[0:0];
  _RAND_1161 = {1{`RANDOM}};
  lru_129 = _RAND_1161[0:0];
  _RAND_1162 = {1{`RANDOM}};
  lru_130 = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  lru_131 = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  lru_132 = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  lru_133 = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  lru_134 = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  lru_135 = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  lru_136 = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  lru_137 = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  lru_138 = _RAND_1170[0:0];
  _RAND_1171 = {1{`RANDOM}};
  lru_139 = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  lru_140 = _RAND_1172[0:0];
  _RAND_1173 = {1{`RANDOM}};
  lru_141 = _RAND_1173[0:0];
  _RAND_1174 = {1{`RANDOM}};
  lru_142 = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  lru_143 = _RAND_1175[0:0];
  _RAND_1176 = {1{`RANDOM}};
  lru_144 = _RAND_1176[0:0];
  _RAND_1177 = {1{`RANDOM}};
  lru_145 = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  lru_146 = _RAND_1178[0:0];
  _RAND_1179 = {1{`RANDOM}};
  lru_147 = _RAND_1179[0:0];
  _RAND_1180 = {1{`RANDOM}};
  lru_148 = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  lru_149 = _RAND_1181[0:0];
  _RAND_1182 = {1{`RANDOM}};
  lru_150 = _RAND_1182[0:0];
  _RAND_1183 = {1{`RANDOM}};
  lru_151 = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  lru_152 = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  lru_153 = _RAND_1185[0:0];
  _RAND_1186 = {1{`RANDOM}};
  lru_154 = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  lru_155 = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  lru_156 = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  lru_157 = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  lru_158 = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  lru_159 = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  lru_160 = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  lru_161 = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  lru_162 = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  lru_163 = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  lru_164 = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  lru_165 = _RAND_1197[0:0];
  _RAND_1198 = {1{`RANDOM}};
  lru_166 = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  lru_167 = _RAND_1199[0:0];
  _RAND_1200 = {1{`RANDOM}};
  lru_168 = _RAND_1200[0:0];
  _RAND_1201 = {1{`RANDOM}};
  lru_169 = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  lru_170 = _RAND_1202[0:0];
  _RAND_1203 = {1{`RANDOM}};
  lru_171 = _RAND_1203[0:0];
  _RAND_1204 = {1{`RANDOM}};
  lru_172 = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  lru_173 = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  lru_174 = _RAND_1206[0:0];
  _RAND_1207 = {1{`RANDOM}};
  lru_175 = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  lru_176 = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  lru_177 = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  lru_178 = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  lru_179 = _RAND_1211[0:0];
  _RAND_1212 = {1{`RANDOM}};
  lru_180 = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  lru_181 = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  lru_182 = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  lru_183 = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  lru_184 = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  lru_185 = _RAND_1217[0:0];
  _RAND_1218 = {1{`RANDOM}};
  lru_186 = _RAND_1218[0:0];
  _RAND_1219 = {1{`RANDOM}};
  lru_187 = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  lru_188 = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  lru_189 = _RAND_1221[0:0];
  _RAND_1222 = {1{`RANDOM}};
  lru_190 = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  lru_191 = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  lru_192 = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  lru_193 = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  lru_194 = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  lru_195 = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  lru_196 = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  lru_197 = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  lru_198 = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  lru_199 = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  lru_200 = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  lru_201 = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  lru_202 = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  lru_203 = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  lru_204 = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  lru_205 = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  lru_206 = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  lru_207 = _RAND_1239[0:0];
  _RAND_1240 = {1{`RANDOM}};
  lru_208 = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  lru_209 = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  lru_210 = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  lru_211 = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  lru_212 = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  lru_213 = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  lru_214 = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  lru_215 = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  lru_216 = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  lru_217 = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  lru_218 = _RAND_1250[0:0];
  _RAND_1251 = {1{`RANDOM}};
  lru_219 = _RAND_1251[0:0];
  _RAND_1252 = {1{`RANDOM}};
  lru_220 = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  lru_221 = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  lru_222 = _RAND_1254[0:0];
  _RAND_1255 = {1{`RANDOM}};
  lru_223 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  lru_224 = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  lru_225 = _RAND_1257[0:0];
  _RAND_1258 = {1{`RANDOM}};
  lru_226 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  lru_227 = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  lru_228 = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  lru_229 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  lru_230 = _RAND_1262[0:0];
  _RAND_1263 = {1{`RANDOM}};
  lru_231 = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  lru_232 = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  lru_233 = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  lru_234 = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  lru_235 = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  lru_236 = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  lru_237 = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  lru_238 = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  lru_239 = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  lru_240 = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  lru_241 = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  lru_242 = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  lru_243 = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  lru_244 = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  lru_245 = _RAND_1277[0:0];
  _RAND_1278 = {1{`RANDOM}};
  lru_246 = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  lru_247 = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  lru_248 = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  lru_249 = _RAND_1281[0:0];
  _RAND_1282 = {1{`RANDOM}};
  lru_250 = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  lru_251 = _RAND_1283[0:0];
  _RAND_1284 = {1{`RANDOM}};
  lru_252 = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  lru_253 = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  lru_254 = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  lru_255 = _RAND_1287[0:0];
  _RAND_1288 = {1{`RANDOM}};
  lru_256 = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  lru_257 = _RAND_1289[0:0];
  _RAND_1290 = {1{`RANDOM}};
  lru_258 = _RAND_1290[0:0];
  _RAND_1291 = {1{`RANDOM}};
  lru_259 = _RAND_1291[0:0];
  _RAND_1292 = {1{`RANDOM}};
  lru_260 = _RAND_1292[0:0];
  _RAND_1293 = {1{`RANDOM}};
  lru_261 = _RAND_1293[0:0];
  _RAND_1294 = {1{`RANDOM}};
  lru_262 = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  lru_263 = _RAND_1295[0:0];
  _RAND_1296 = {1{`RANDOM}};
  lru_264 = _RAND_1296[0:0];
  _RAND_1297 = {1{`RANDOM}};
  lru_265 = _RAND_1297[0:0];
  _RAND_1298 = {1{`RANDOM}};
  lru_266 = _RAND_1298[0:0];
  _RAND_1299 = {1{`RANDOM}};
  lru_267 = _RAND_1299[0:0];
  _RAND_1300 = {1{`RANDOM}};
  lru_268 = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  lru_269 = _RAND_1301[0:0];
  _RAND_1302 = {1{`RANDOM}};
  lru_270 = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  lru_271 = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  lru_272 = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  lru_273 = _RAND_1305[0:0];
  _RAND_1306 = {1{`RANDOM}};
  lru_274 = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  lru_275 = _RAND_1307[0:0];
  _RAND_1308 = {1{`RANDOM}};
  lru_276 = _RAND_1308[0:0];
  _RAND_1309 = {1{`RANDOM}};
  lru_277 = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  lru_278 = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  lru_279 = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  lru_280 = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  lru_281 = _RAND_1313[0:0];
  _RAND_1314 = {1{`RANDOM}};
  lru_282 = _RAND_1314[0:0];
  _RAND_1315 = {1{`RANDOM}};
  lru_283 = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  lru_284 = _RAND_1316[0:0];
  _RAND_1317 = {1{`RANDOM}};
  lru_285 = _RAND_1317[0:0];
  _RAND_1318 = {1{`RANDOM}};
  lru_286 = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  lru_287 = _RAND_1319[0:0];
  _RAND_1320 = {1{`RANDOM}};
  lru_288 = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  lru_289 = _RAND_1321[0:0];
  _RAND_1322 = {1{`RANDOM}};
  lru_290 = _RAND_1322[0:0];
  _RAND_1323 = {1{`RANDOM}};
  lru_291 = _RAND_1323[0:0];
  _RAND_1324 = {1{`RANDOM}};
  lru_292 = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  lru_293 = _RAND_1325[0:0];
  _RAND_1326 = {1{`RANDOM}};
  lru_294 = _RAND_1326[0:0];
  _RAND_1327 = {1{`RANDOM}};
  lru_295 = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  lru_296 = _RAND_1328[0:0];
  _RAND_1329 = {1{`RANDOM}};
  lru_297 = _RAND_1329[0:0];
  _RAND_1330 = {1{`RANDOM}};
  lru_298 = _RAND_1330[0:0];
  _RAND_1331 = {1{`RANDOM}};
  lru_299 = _RAND_1331[0:0];
  _RAND_1332 = {1{`RANDOM}};
  lru_300 = _RAND_1332[0:0];
  _RAND_1333 = {1{`RANDOM}};
  lru_301 = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  lru_302 = _RAND_1334[0:0];
  _RAND_1335 = {1{`RANDOM}};
  lru_303 = _RAND_1335[0:0];
  _RAND_1336 = {1{`RANDOM}};
  lru_304 = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  lru_305 = _RAND_1337[0:0];
  _RAND_1338 = {1{`RANDOM}};
  lru_306 = _RAND_1338[0:0];
  _RAND_1339 = {1{`RANDOM}};
  lru_307 = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  lru_308 = _RAND_1340[0:0];
  _RAND_1341 = {1{`RANDOM}};
  lru_309 = _RAND_1341[0:0];
  _RAND_1342 = {1{`RANDOM}};
  lru_310 = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  lru_311 = _RAND_1343[0:0];
  _RAND_1344 = {1{`RANDOM}};
  lru_312 = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  lru_313 = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  lru_314 = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  lru_315 = _RAND_1347[0:0];
  _RAND_1348 = {1{`RANDOM}};
  lru_316 = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  lru_317 = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  lru_318 = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  lru_319 = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  lru_320 = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  lru_321 = _RAND_1353[0:0];
  _RAND_1354 = {1{`RANDOM}};
  lru_322 = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  lru_323 = _RAND_1355[0:0];
  _RAND_1356 = {1{`RANDOM}};
  lru_324 = _RAND_1356[0:0];
  _RAND_1357 = {1{`RANDOM}};
  lru_325 = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  lru_326 = _RAND_1358[0:0];
  _RAND_1359 = {1{`RANDOM}};
  lru_327 = _RAND_1359[0:0];
  _RAND_1360 = {1{`RANDOM}};
  lru_328 = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  lru_329 = _RAND_1361[0:0];
  _RAND_1362 = {1{`RANDOM}};
  lru_330 = _RAND_1362[0:0];
  _RAND_1363 = {1{`RANDOM}};
  lru_331 = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  lru_332 = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  lru_333 = _RAND_1365[0:0];
  _RAND_1366 = {1{`RANDOM}};
  lru_334 = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  lru_335 = _RAND_1367[0:0];
  _RAND_1368 = {1{`RANDOM}};
  lru_336 = _RAND_1368[0:0];
  _RAND_1369 = {1{`RANDOM}};
  lru_337 = _RAND_1369[0:0];
  _RAND_1370 = {1{`RANDOM}};
  lru_338 = _RAND_1370[0:0];
  _RAND_1371 = {1{`RANDOM}};
  lru_339 = _RAND_1371[0:0];
  _RAND_1372 = {1{`RANDOM}};
  lru_340 = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  lru_341 = _RAND_1373[0:0];
  _RAND_1374 = {1{`RANDOM}};
  lru_342 = _RAND_1374[0:0];
  _RAND_1375 = {1{`RANDOM}};
  lru_343 = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  lru_344 = _RAND_1376[0:0];
  _RAND_1377 = {1{`RANDOM}};
  lru_345 = _RAND_1377[0:0];
  _RAND_1378 = {1{`RANDOM}};
  lru_346 = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  lru_347 = _RAND_1379[0:0];
  _RAND_1380 = {1{`RANDOM}};
  lru_348 = _RAND_1380[0:0];
  _RAND_1381 = {1{`RANDOM}};
  lru_349 = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  lru_350 = _RAND_1382[0:0];
  _RAND_1383 = {1{`RANDOM}};
  lru_351 = _RAND_1383[0:0];
  _RAND_1384 = {1{`RANDOM}};
  lru_352 = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  lru_353 = _RAND_1385[0:0];
  _RAND_1386 = {1{`RANDOM}};
  lru_354 = _RAND_1386[0:0];
  _RAND_1387 = {1{`RANDOM}};
  lru_355 = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  lru_356 = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  lru_357 = _RAND_1389[0:0];
  _RAND_1390 = {1{`RANDOM}};
  lru_358 = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  lru_359 = _RAND_1391[0:0];
  _RAND_1392 = {1{`RANDOM}};
  lru_360 = _RAND_1392[0:0];
  _RAND_1393 = {1{`RANDOM}};
  lru_361 = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  lru_362 = _RAND_1394[0:0];
  _RAND_1395 = {1{`RANDOM}};
  lru_363 = _RAND_1395[0:0];
  _RAND_1396 = {1{`RANDOM}};
  lru_364 = _RAND_1396[0:0];
  _RAND_1397 = {1{`RANDOM}};
  lru_365 = _RAND_1397[0:0];
  _RAND_1398 = {1{`RANDOM}};
  lru_366 = _RAND_1398[0:0];
  _RAND_1399 = {1{`RANDOM}};
  lru_367 = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  lru_368 = _RAND_1400[0:0];
  _RAND_1401 = {1{`RANDOM}};
  lru_369 = _RAND_1401[0:0];
  _RAND_1402 = {1{`RANDOM}};
  lru_370 = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  lru_371 = _RAND_1403[0:0];
  _RAND_1404 = {1{`RANDOM}};
  lru_372 = _RAND_1404[0:0];
  _RAND_1405 = {1{`RANDOM}};
  lru_373 = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  lru_374 = _RAND_1406[0:0];
  _RAND_1407 = {1{`RANDOM}};
  lru_375 = _RAND_1407[0:0];
  _RAND_1408 = {1{`RANDOM}};
  lru_376 = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  lru_377 = _RAND_1409[0:0];
  _RAND_1410 = {1{`RANDOM}};
  lru_378 = _RAND_1410[0:0];
  _RAND_1411 = {1{`RANDOM}};
  lru_379 = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  lru_380 = _RAND_1412[0:0];
  _RAND_1413 = {1{`RANDOM}};
  lru_381 = _RAND_1413[0:0];
  _RAND_1414 = {1{`RANDOM}};
  lru_382 = _RAND_1414[0:0];
  _RAND_1415 = {1{`RANDOM}};
  lru_383 = _RAND_1415[0:0];
  _RAND_1416 = {1{`RANDOM}};
  lru_384 = _RAND_1416[0:0];
  _RAND_1417 = {1{`RANDOM}};
  lru_385 = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  lru_386 = _RAND_1418[0:0];
  _RAND_1419 = {1{`RANDOM}};
  lru_387 = _RAND_1419[0:0];
  _RAND_1420 = {1{`RANDOM}};
  lru_388 = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  lru_389 = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  lru_390 = _RAND_1422[0:0];
  _RAND_1423 = {1{`RANDOM}};
  lru_391 = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  lru_392 = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  lru_393 = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  lru_394 = _RAND_1426[0:0];
  _RAND_1427 = {1{`RANDOM}};
  lru_395 = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  lru_396 = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  lru_397 = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  lru_398 = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  lru_399 = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  lru_400 = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  lru_401 = _RAND_1433[0:0];
  _RAND_1434 = {1{`RANDOM}};
  lru_402 = _RAND_1434[0:0];
  _RAND_1435 = {1{`RANDOM}};
  lru_403 = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  lru_404 = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  lru_405 = _RAND_1437[0:0];
  _RAND_1438 = {1{`RANDOM}};
  lru_406 = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  lru_407 = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  lru_408 = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  lru_409 = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  lru_410 = _RAND_1442[0:0];
  _RAND_1443 = {1{`RANDOM}};
  lru_411 = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  lru_412 = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  lru_413 = _RAND_1445[0:0];
  _RAND_1446 = {1{`RANDOM}};
  lru_414 = _RAND_1446[0:0];
  _RAND_1447 = {1{`RANDOM}};
  lru_415 = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  lru_416 = _RAND_1448[0:0];
  _RAND_1449 = {1{`RANDOM}};
  lru_417 = _RAND_1449[0:0];
  _RAND_1450 = {1{`RANDOM}};
  lru_418 = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  lru_419 = _RAND_1451[0:0];
  _RAND_1452 = {1{`RANDOM}};
  lru_420 = _RAND_1452[0:0];
  _RAND_1453 = {1{`RANDOM}};
  lru_421 = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  lru_422 = _RAND_1454[0:0];
  _RAND_1455 = {1{`RANDOM}};
  lru_423 = _RAND_1455[0:0];
  _RAND_1456 = {1{`RANDOM}};
  lru_424 = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  lru_425 = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  lru_426 = _RAND_1458[0:0];
  _RAND_1459 = {1{`RANDOM}};
  lru_427 = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  lru_428 = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  lru_429 = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  lru_430 = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  lru_431 = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  lru_432 = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  lru_433 = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  lru_434 = _RAND_1466[0:0];
  _RAND_1467 = {1{`RANDOM}};
  lru_435 = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  lru_436 = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  lru_437 = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  lru_438 = _RAND_1470[0:0];
  _RAND_1471 = {1{`RANDOM}};
  lru_439 = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  lru_440 = _RAND_1472[0:0];
  _RAND_1473 = {1{`RANDOM}};
  lru_441 = _RAND_1473[0:0];
  _RAND_1474 = {1{`RANDOM}};
  lru_442 = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  lru_443 = _RAND_1475[0:0];
  _RAND_1476 = {1{`RANDOM}};
  lru_444 = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  lru_445 = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  lru_446 = _RAND_1478[0:0];
  _RAND_1479 = {1{`RANDOM}};
  lru_447 = _RAND_1479[0:0];
  _RAND_1480 = {1{`RANDOM}};
  lru_448 = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  lru_449 = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  lru_450 = _RAND_1482[0:0];
  _RAND_1483 = {1{`RANDOM}};
  lru_451 = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  lru_452 = _RAND_1484[0:0];
  _RAND_1485 = {1{`RANDOM}};
  lru_453 = _RAND_1485[0:0];
  _RAND_1486 = {1{`RANDOM}};
  lru_454 = _RAND_1486[0:0];
  _RAND_1487 = {1{`RANDOM}};
  lru_455 = _RAND_1487[0:0];
  _RAND_1488 = {1{`RANDOM}};
  lru_456 = _RAND_1488[0:0];
  _RAND_1489 = {1{`RANDOM}};
  lru_457 = _RAND_1489[0:0];
  _RAND_1490 = {1{`RANDOM}};
  lru_458 = _RAND_1490[0:0];
  _RAND_1491 = {1{`RANDOM}};
  lru_459 = _RAND_1491[0:0];
  _RAND_1492 = {1{`RANDOM}};
  lru_460 = _RAND_1492[0:0];
  _RAND_1493 = {1{`RANDOM}};
  lru_461 = _RAND_1493[0:0];
  _RAND_1494 = {1{`RANDOM}};
  lru_462 = _RAND_1494[0:0];
  _RAND_1495 = {1{`RANDOM}};
  lru_463 = _RAND_1495[0:0];
  _RAND_1496 = {1{`RANDOM}};
  lru_464 = _RAND_1496[0:0];
  _RAND_1497 = {1{`RANDOM}};
  lru_465 = _RAND_1497[0:0];
  _RAND_1498 = {1{`RANDOM}};
  lru_466 = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  lru_467 = _RAND_1499[0:0];
  _RAND_1500 = {1{`RANDOM}};
  lru_468 = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  lru_469 = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  lru_470 = _RAND_1502[0:0];
  _RAND_1503 = {1{`RANDOM}};
  lru_471 = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  lru_472 = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  lru_473 = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  lru_474 = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  lru_475 = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  lru_476 = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  lru_477 = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  lru_478 = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  lru_479 = _RAND_1511[0:0];
  _RAND_1512 = {1{`RANDOM}};
  lru_480 = _RAND_1512[0:0];
  _RAND_1513 = {1{`RANDOM}};
  lru_481 = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  lru_482 = _RAND_1514[0:0];
  _RAND_1515 = {1{`RANDOM}};
  lru_483 = _RAND_1515[0:0];
  _RAND_1516 = {1{`RANDOM}};
  lru_484 = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  lru_485 = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  lru_486 = _RAND_1518[0:0];
  _RAND_1519 = {1{`RANDOM}};
  lru_487 = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  lru_488 = _RAND_1520[0:0];
  _RAND_1521 = {1{`RANDOM}};
  lru_489 = _RAND_1521[0:0];
  _RAND_1522 = {1{`RANDOM}};
  lru_490 = _RAND_1522[0:0];
  _RAND_1523 = {1{`RANDOM}};
  lru_491 = _RAND_1523[0:0];
  _RAND_1524 = {1{`RANDOM}};
  lru_492 = _RAND_1524[0:0];
  _RAND_1525 = {1{`RANDOM}};
  lru_493 = _RAND_1525[0:0];
  _RAND_1526 = {1{`RANDOM}};
  lru_494 = _RAND_1526[0:0];
  _RAND_1527 = {1{`RANDOM}};
  lru_495 = _RAND_1527[0:0];
  _RAND_1528 = {1{`RANDOM}};
  lru_496 = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  lru_497 = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  lru_498 = _RAND_1530[0:0];
  _RAND_1531 = {1{`RANDOM}};
  lru_499 = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  lru_500 = _RAND_1532[0:0];
  _RAND_1533 = {1{`RANDOM}};
  lru_501 = _RAND_1533[0:0];
  _RAND_1534 = {1{`RANDOM}};
  lru_502 = _RAND_1534[0:0];
  _RAND_1535 = {1{`RANDOM}};
  lru_503 = _RAND_1535[0:0];
  _RAND_1536 = {1{`RANDOM}};
  lru_504 = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  lru_505 = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  lru_506 = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  lru_507 = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  lru_508 = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  lru_509 = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  lru_510 = _RAND_1542[0:0];
  _RAND_1543 = {1{`RANDOM}};
  lru_511 = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  tlb_vpn = _RAND_1544[19:0];
  _RAND_1545 = {1{`RANDOM}};
  tlb_ppn = _RAND_1545[19:0];
  _RAND_1546 = {1{`RANDOM}};
  tlb_uncached = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  tlb_valid = _RAND_1547[0:0];
  _RAND_1548 = {1{`RANDOM}};
  rset = _RAND_1548[5:0];
  _RAND_1549 = {1{`RANDOM}};
  saved_0_inst = _RAND_1549[31:0];
  _RAND_1550 = {1{`RANDOM}};
  saved_0_valid = _RAND_1550[0:0];
  _RAND_1551 = {1{`RANDOM}};
  saved_1_inst = _RAND_1551[31:0];
  _RAND_1552 = {1{`RANDOM}};
  saved_1_valid = _RAND_1552[0:0];
  _RAND_1553 = {1{`RANDOM}};
  axi_cnt_value = _RAND_1553[4:0];
  _RAND_1554 = {1{`RANDOM}};
  ar_addr = _RAND_1554[31:0];
  _RAND_1555 = {1{`RANDOM}};
  ar_len = _RAND_1555[7:0];
  _RAND_1556 = {1{`RANDOM}};
  ar_size = _RAND_1556[2:0];
  _RAND_1557 = {1{`RANDOM}};
  arvalid = _RAND_1557[0:0];
  _RAND_1558 = {1{`RANDOM}};
  rready = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  tlb1_invalid = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  io_cpu_tlb2_vpn_r = _RAND_1560[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input  [31:0] io_enq_bits_addr,
  input  [3:0]  io_enq_bits_strb,
  input  [1:0]  io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output [31:0] io_deq_bits_addr,
  output [3:0]  io_deq_bits_strb,
  output [1:0]  io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_data [0:3]; // @[Decoupled.scala 275:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 275:95]
  wire [1:0] ram_data_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 275:95]
  reg [31:0] ram_addr [0:3]; // @[Decoupled.scala 275:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [1:0] ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [31:0] ram_addr_MPORT_data; // @[Decoupled.scala 275:95]
  wire [1:0] ram_addr_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 275:95]
  reg [3:0] ram_strb [0:3]; // @[Decoupled.scala 275:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [1:0] ram_strb_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [3:0] ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [3:0] ram_strb_MPORT_data; // @[Decoupled.scala 275:95]
  wire [1:0] ram_strb_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_strb_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_strb_MPORT_en; // @[Decoupled.scala 275:95]
  reg [1:0] ram_size [0:3]; // @[Decoupled.scala 275:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [1:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 275:95]
  wire [1:0] ram_size_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 275:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = enq_ptr_value;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  assign io_deq_bits_strb = ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_strb[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enq_ptr_value = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  deq_ptr_value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleDualPortRam_8(
  input         clock,
  input         reset,
  input  [9:0]  io_raddr,
  output [31:0] io_rdata,
  input  [9:0]  io_waddr,
  input         io_wen,
  input  [3:0]  io_wstrb,
  input  [31:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] bank_0 [0:1023]; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_0_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  wire [9:0] bank_0_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_0_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_0_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [9:0] bank_0_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_0_MPORT_mask; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_0_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  reg  bank_0_io_rdata_MPORT_en_pipe_0;
  reg [9:0] bank_0_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_1 [0:1023]; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_1_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  wire [9:0] bank_1_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_1_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_1_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [9:0] bank_1_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_1_MPORT_mask; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_1_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  reg  bank_1_io_rdata_MPORT_en_pipe_0;
  reg [9:0] bank_1_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_2 [0:1023]; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_2_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  wire [9:0] bank_2_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_2_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_2_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [9:0] bank_2_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_2_MPORT_mask; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_2_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  reg  bank_2_io_rdata_MPORT_en_pipe_0;
  reg [9:0] bank_2_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_3 [0:1023]; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_3_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  wire [9:0] bank_3_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_3_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [7:0] bank_3_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
  wire [9:0] bank_3_MPORT_addr; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_3_MPORT_mask; // @[SimpleDualPortRam.scala 68:29]
  wire  bank_3_MPORT_en; // @[SimpleDualPortRam.scala 68:29]
  reg  bank_3_io_rdata_MPORT_en_pipe_0;
  reg [9:0] bank_3_io_rdata_MPORT_addr_pipe_0;
  wire  _T_2 = |io_wstrb | ~io_wen; // @[SimpleDualPortRam.scala 64:20]
  wire [15:0] io_rdata_lo = {bank_1_io_rdata_MPORT_data,bank_0_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 70:44]
  wire [15:0] io_rdata_hi = {bank_3_io_rdata_MPORT_data,bank_2_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 70:44]
  assign bank_0_io_rdata_MPORT_en = bank_0_io_rdata_MPORT_en_pipe_0;
  assign bank_0_io_rdata_MPORT_addr = bank_0_io_rdata_MPORT_addr_pipe_0;
  assign bank_0_io_rdata_MPORT_data = bank_0[bank_0_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 68:29]
  assign bank_0_MPORT_data = io_wdata[7:0];
  assign bank_0_MPORT_addr = io_waddr;
  assign bank_0_MPORT_mask = io_wstrb[0];
  assign bank_0_MPORT_en = io_wen;
  assign bank_1_io_rdata_MPORT_en = bank_1_io_rdata_MPORT_en_pipe_0;
  assign bank_1_io_rdata_MPORT_addr = bank_1_io_rdata_MPORT_addr_pipe_0;
  assign bank_1_io_rdata_MPORT_data = bank_1[bank_1_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 68:29]
  assign bank_1_MPORT_data = io_wdata[15:8];
  assign bank_1_MPORT_addr = io_waddr;
  assign bank_1_MPORT_mask = io_wstrb[1];
  assign bank_1_MPORT_en = io_wen;
  assign bank_2_io_rdata_MPORT_en = bank_2_io_rdata_MPORT_en_pipe_0;
  assign bank_2_io_rdata_MPORT_addr = bank_2_io_rdata_MPORT_addr_pipe_0;
  assign bank_2_io_rdata_MPORT_data = bank_2[bank_2_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 68:29]
  assign bank_2_MPORT_data = io_wdata[23:16];
  assign bank_2_MPORT_addr = io_waddr;
  assign bank_2_MPORT_mask = io_wstrb[2];
  assign bank_2_MPORT_en = io_wen;
  assign bank_3_io_rdata_MPORT_en = bank_3_io_rdata_MPORT_en_pipe_0;
  assign bank_3_io_rdata_MPORT_addr = bank_3_io_rdata_MPORT_addr_pipe_0;
  assign bank_3_io_rdata_MPORT_data = bank_3[bank_3_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 68:29]
  assign bank_3_MPORT_data = io_wdata[31:24];
  assign bank_3_MPORT_addr = io_waddr;
  assign bank_3_MPORT_mask = io_wstrb[3];
  assign bank_3_MPORT_en = io_wen;
  assign io_rdata = {io_rdata_hi,io_rdata_lo}; // @[SimpleDualPortRam.scala 70:44]
  always @(posedge clock) begin
    if (bank_0_MPORT_en & bank_0_MPORT_mask) begin
      bank_0[bank_0_MPORT_addr] <= bank_0_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
    end
    bank_0_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_0_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_1_MPORT_en & bank_1_MPORT_mask) begin
      bank_1[bank_1_MPORT_addr] <= bank_1_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
    end
    bank_1_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_1_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_2_MPORT_en & bank_2_MPORT_mask) begin
      bank_2[bank_2_MPORT_addr] <= bank_2_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
    end
    bank_2_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_2_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_3_MPORT_en & bank_3_MPORT_mask) begin
      bank_3[bank_3_MPORT_addr] <= bank_3_MPORT_data; // @[SimpleDualPortRam.scala 68:29]
    end
    bank_3_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_3_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed: when write port enable is high, write vector cannot be all 0\n    at SimpleDualPortRam.scala:63 assert(\n"
            ); // @[SimpleDualPortRam.scala 63:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & ~reset) begin
          $fatal; // @[SimpleDualPortRam.scala 63:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    bank_0[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    bank_1[initvar] = _RAND_3[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    bank_2[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    bank_3[initvar] = _RAND_9[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bank_0_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bank_0_io_rdata_MPORT_addr_pipe_0 = _RAND_2[9:0];
  _RAND_4 = {1{`RANDOM}};
  bank_1_io_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  bank_1_io_rdata_MPORT_addr_pipe_0 = _RAND_5[9:0];
  _RAND_7 = {1{`RANDOM}};
  bank_2_io_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  bank_2_io_rdata_MPORT_addr_pipe_0 = _RAND_8[9:0];
  _RAND_10 = {1{`RANDOM}};
  bank_3_io_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  bank_3_io_rdata_MPORT_addr_pipe_0 = _RAND_11[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleDualPortRam_9(
  input         clock,
  input         reset,
  input  [6:0]  io_raddr,
  output [19:0] io_rdata,
  input  [6:0]  io_waddr,
  input         io_wen,
  input         io_wstrb,
  input  [19:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] bank [0:127]; // @[SimpleDualPortRam.scala 78:29]
  wire  bank_io_rdata_MPORT_en; // @[SimpleDualPortRam.scala 78:29]
  wire [6:0] bank_io_rdata_MPORT_addr; // @[SimpleDualPortRam.scala 78:29]
  wire [19:0] bank_io_rdata_MPORT_data; // @[SimpleDualPortRam.scala 78:29]
  wire [19:0] bank_MPORT_data; // @[SimpleDualPortRam.scala 78:29]
  wire [6:0] bank_MPORT_addr; // @[SimpleDualPortRam.scala 78:29]
  wire  bank_MPORT_mask; // @[SimpleDualPortRam.scala 78:29]
  wire  bank_MPORT_en; // @[SimpleDualPortRam.scala 78:29]
  reg  bank_io_rdata_MPORT_en_pipe_0;
  reg [6:0] bank_io_rdata_MPORT_addr_pipe_0;
  wire  _T_2 = |io_wstrb | ~io_wen; // @[SimpleDualPortRam.scala 64:20]
  wire [31:0] _GEN_7 = {{12'd0}, bank_io_rdata_MPORT_data}; // @[SimpleDualPortRam.scala 80:20 81:18 83:18]
  assign bank_io_rdata_MPORT_en = bank_io_rdata_MPORT_en_pipe_0;
  assign bank_io_rdata_MPORT_addr = bank_io_rdata_MPORT_addr_pipe_0;
  assign bank_io_rdata_MPORT_data = bank[bank_io_rdata_MPORT_addr]; // @[SimpleDualPortRam.scala 78:29]
  assign bank_MPORT_data = io_wdata;
  assign bank_MPORT_addr = io_waddr;
  assign bank_MPORT_mask = 1'h1;
  assign bank_MPORT_en = io_wen;
  assign io_rdata = _GEN_7[19:0];
  always @(posedge clock) begin
    if (bank_MPORT_en & bank_MPORT_mask) begin
      bank[bank_MPORT_addr] <= bank_MPORT_data; // @[SimpleDualPortRam.scala 78:29]
    end
    bank_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed: when write port enable is high, write vector cannot be all 0\n    at SimpleDualPortRam.scala:63 assert(\n"
            ); // @[SimpleDualPortRam.scala 63:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & ~reset) begin
          $fatal; // @[SimpleDualPortRam.scala 63:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    bank[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bank_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bank_io_rdata_MPORT_addr_pipe_0 = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input         clock,
  input         reset,
  input         io_cpu_stallM,
  output        io_cpu_dstall,
  input  [31:0] io_cpu_E_mem_va,
  input  [31:0] io_cpu_M_mem_va,
  input  [31:0] io_cpu_M_fence_addr,
  input         io_cpu_M_fence_d,
  input         io_cpu_M_mem_en,
  input         io_cpu_M_mem_write,
  input  [3:0]  io_cpu_M_wmask,
  input  [1:0]  io_cpu_M_mem_size,
  input  [31:0] io_cpu_M_wdata,
  output [31:0] io_cpu_M_rdata,
  output [18:0] io_cpu_tlb_vpn2,
  input         io_cpu_tlb_found,
  input  [19:0] io_cpu_tlb_entry_pfn_0,
  input  [19:0] io_cpu_tlb_entry_pfn_1,
  input         io_cpu_tlb_entry_c_0,
  input         io_cpu_tlb_entry_c_1,
  input         io_cpu_tlb_entry_d_0,
  input         io_cpu_tlb_entry_d_1,
  input         io_cpu_tlb_entry_v_0,
  input         io_cpu_tlb_entry_v_1,
  input         io_cpu_fence_tlb,
  output        io_cpu_data_tlb_refill,
  output        io_cpu_data_tlb_invalid,
  output        io_cpu_data_tlb_mod,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output [7:0]  io_axi_ar_bits_len,
  output [2:0]  io_axi_ar_bits_size,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [31:0] io_axi_r_bits_data,
  input         io_axi_r_bits_last,
  input         io_axi_aw_ready,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  output [7:0]  io_axi_aw_bits_len,
  output [2:0]  io_axi_aw_bits_size,
  input         io_axi_w_ready,
  output        io_axi_w_valid,
  output [31:0] io_axi_w_bits_data,
  output [3:0]  io_axi_w_bits_strb,
  output        io_axi_w_bits_last,
  output        io_axi_b_ready,
  input         io_axi_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
`endif // RANDOMIZE_REG_INIT
  wire  write_buffer_clock; // @[DCache.scala 82:28]
  wire  write_buffer_reset; // @[DCache.scala 82:28]
  wire  write_buffer_io_enq_ready; // @[DCache.scala 82:28]
  wire  write_buffer_io_enq_valid; // @[DCache.scala 82:28]
  wire [31:0] write_buffer_io_enq_bits_data; // @[DCache.scala 82:28]
  wire [31:0] write_buffer_io_enq_bits_addr; // @[DCache.scala 82:28]
  wire [3:0] write_buffer_io_enq_bits_strb; // @[DCache.scala 82:28]
  wire [1:0] write_buffer_io_enq_bits_size; // @[DCache.scala 82:28]
  wire  write_buffer_io_deq_ready; // @[DCache.scala 82:28]
  wire  write_buffer_io_deq_valid; // @[DCache.scala 82:28]
  wire [31:0] write_buffer_io_deq_bits_data; // @[DCache.scala 82:28]
  wire [31:0] write_buffer_io_deq_bits_addr; // @[DCache.scala 82:28]
  wire [3:0] write_buffer_io_deq_bits_strb; // @[DCache.scala 82:28]
  wire [1:0] write_buffer_io_deq_bits_size; // @[DCache.scala 82:28]
  wire  bank_ram_clock; // @[DCache.scala 153:26]
  wire  bank_ram_reset; // @[DCache.scala 153:26]
  wire [9:0] bank_ram_io_raddr; // @[DCache.scala 153:26]
  wire [31:0] bank_ram_io_rdata; // @[DCache.scala 153:26]
  wire [9:0] bank_ram_io_waddr; // @[DCache.scala 153:26]
  wire  bank_ram_io_wen; // @[DCache.scala 153:26]
  wire [3:0] bank_ram_io_wstrb; // @[DCache.scala 153:26]
  wire [31:0] bank_ram_io_wdata; // @[DCache.scala 153:26]
  wire  tag_ram_clock; // @[DCache.scala 163:25]
  wire  tag_ram_reset; // @[DCache.scala 163:25]
  wire [6:0] tag_ram_io_raddr; // @[DCache.scala 163:25]
  wire [19:0] tag_ram_io_rdata; // @[DCache.scala 163:25]
  wire [6:0] tag_ram_io_waddr; // @[DCache.scala 163:25]
  wire  tag_ram_io_wen; // @[DCache.scala 163:25]
  wire  tag_ram_io_wstrb; // @[DCache.scala 163:25]
  wire [19:0] tag_ram_io_wdata; // @[DCache.scala 163:25]
  wire  bank_ram_1_clock; // @[DCache.scala 153:26]
  wire  bank_ram_1_reset; // @[DCache.scala 153:26]
  wire [9:0] bank_ram_1_io_raddr; // @[DCache.scala 153:26]
  wire [31:0] bank_ram_1_io_rdata; // @[DCache.scala 153:26]
  wire [9:0] bank_ram_1_io_waddr; // @[DCache.scala 153:26]
  wire  bank_ram_1_io_wen; // @[DCache.scala 153:26]
  wire [3:0] bank_ram_1_io_wstrb; // @[DCache.scala 153:26]
  wire [31:0] bank_ram_1_io_wdata; // @[DCache.scala 153:26]
  wire  tag_ram_1_clock; // @[DCache.scala 163:25]
  wire  tag_ram_1_reset; // @[DCache.scala 163:25]
  wire [6:0] tag_ram_1_io_raddr; // @[DCache.scala 163:25]
  wire [19:0] tag_ram_1_io_rdata; // @[DCache.scala 163:25]
  wire [6:0] tag_ram_1_io_waddr; // @[DCache.scala 163:25]
  wire  tag_ram_1_io_wen; // @[DCache.scala 163:25]
  wire  tag_ram_1_io_wstrb; // @[DCache.scala 163:25]
  wire [19:0] tag_ram_1_io_wdata; // @[DCache.scala 163:25]
  reg [19:0] tlb_vpn; // @[DCache.scala 46:20]
  reg [19:0] tlb_ppn; // @[DCache.scala 46:20]
  reg  tlb_uncached; // @[DCache.scala 46:20]
  reg  tlb_dirty; // @[DCache.scala 46:20]
  reg  tlb_valid; // @[DCache.scala 46:20]
  wire  direct_mapped = io_cpu_M_mem_va[31:30] == 2'h2; // @[DCache.scala 54:41]
  wire  M_mem_uncached = direct_mapped ? io_cpu_M_mem_va[29] : tlb_uncached; // @[DCache.scala 55:27]
  wire [19:0] _data_tag_T_1 = {3'h0,io_cpu_M_mem_va[28:12]}; // @[Cat.scala 33:92]
  wire [19:0] data_tag = direct_mapped ? _data_tag_T_1 : tlb_ppn; // @[DCache.scala 56:27]
  wire [19:0] data_vpn = io_cpu_M_mem_va[31:12]; // @[DCache.scala 57:32]
  wire [31:0] M_mem_pa = {data_tag,io_cpu_M_mem_va[11:0]}; // @[Cat.scala 33:92]
  wire  l1tlb_ok = tlb_vpn == data_vpn & tlb_valid; // @[DCache.scala 60:40]
  wire  _translation_ok_T_2 = ~io_cpu_M_mem_write; // @[DCache.scala 62:61]
  wire  translation_ok = direct_mapped | l1tlb_ok & (~io_cpu_M_mem_write | tlb_dirty); // @[DCache.scala 62:19]
  reg [2:0] state; // @[DCache.scala 65:96]
  reg  valid_0_0; // @[DCache.scala 68:22]
  reg  valid_0_1; // @[DCache.scala 68:22]
  reg  valid_1_0; // @[DCache.scala 68:22]
  reg  valid_1_1; // @[DCache.scala 68:22]
  reg  valid_2_0; // @[DCache.scala 68:22]
  reg  valid_2_1; // @[DCache.scala 68:22]
  reg  valid_3_0; // @[DCache.scala 68:22]
  reg  valid_3_1; // @[DCache.scala 68:22]
  reg  valid_4_0; // @[DCache.scala 68:22]
  reg  valid_4_1; // @[DCache.scala 68:22]
  reg  valid_5_0; // @[DCache.scala 68:22]
  reg  valid_5_1; // @[DCache.scala 68:22]
  reg  valid_6_0; // @[DCache.scala 68:22]
  reg  valid_6_1; // @[DCache.scala 68:22]
  reg  valid_7_0; // @[DCache.scala 68:22]
  reg  valid_7_1; // @[DCache.scala 68:22]
  reg  valid_8_0; // @[DCache.scala 68:22]
  reg  valid_8_1; // @[DCache.scala 68:22]
  reg  valid_9_0; // @[DCache.scala 68:22]
  reg  valid_9_1; // @[DCache.scala 68:22]
  reg  valid_10_0; // @[DCache.scala 68:22]
  reg  valid_10_1; // @[DCache.scala 68:22]
  reg  valid_11_0; // @[DCache.scala 68:22]
  reg  valid_11_1; // @[DCache.scala 68:22]
  reg  valid_12_0; // @[DCache.scala 68:22]
  reg  valid_12_1; // @[DCache.scala 68:22]
  reg  valid_13_0; // @[DCache.scala 68:22]
  reg  valid_13_1; // @[DCache.scala 68:22]
  reg  valid_14_0; // @[DCache.scala 68:22]
  reg  valid_14_1; // @[DCache.scala 68:22]
  reg  valid_15_0; // @[DCache.scala 68:22]
  reg  valid_15_1; // @[DCache.scala 68:22]
  reg  valid_16_0; // @[DCache.scala 68:22]
  reg  valid_16_1; // @[DCache.scala 68:22]
  reg  valid_17_0; // @[DCache.scala 68:22]
  reg  valid_17_1; // @[DCache.scala 68:22]
  reg  valid_18_0; // @[DCache.scala 68:22]
  reg  valid_18_1; // @[DCache.scala 68:22]
  reg  valid_19_0; // @[DCache.scala 68:22]
  reg  valid_19_1; // @[DCache.scala 68:22]
  reg  valid_20_0; // @[DCache.scala 68:22]
  reg  valid_20_1; // @[DCache.scala 68:22]
  reg  valid_21_0; // @[DCache.scala 68:22]
  reg  valid_21_1; // @[DCache.scala 68:22]
  reg  valid_22_0; // @[DCache.scala 68:22]
  reg  valid_22_1; // @[DCache.scala 68:22]
  reg  valid_23_0; // @[DCache.scala 68:22]
  reg  valid_23_1; // @[DCache.scala 68:22]
  reg  valid_24_0; // @[DCache.scala 68:22]
  reg  valid_24_1; // @[DCache.scala 68:22]
  reg  valid_25_0; // @[DCache.scala 68:22]
  reg  valid_25_1; // @[DCache.scala 68:22]
  reg  valid_26_0; // @[DCache.scala 68:22]
  reg  valid_26_1; // @[DCache.scala 68:22]
  reg  valid_27_0; // @[DCache.scala 68:22]
  reg  valid_27_1; // @[DCache.scala 68:22]
  reg  valid_28_0; // @[DCache.scala 68:22]
  reg  valid_28_1; // @[DCache.scala 68:22]
  reg  valid_29_0; // @[DCache.scala 68:22]
  reg  valid_29_1; // @[DCache.scala 68:22]
  reg  valid_30_0; // @[DCache.scala 68:22]
  reg  valid_30_1; // @[DCache.scala 68:22]
  reg  valid_31_0; // @[DCache.scala 68:22]
  reg  valid_31_1; // @[DCache.scala 68:22]
  reg  valid_32_0; // @[DCache.scala 68:22]
  reg  valid_32_1; // @[DCache.scala 68:22]
  reg  valid_33_0; // @[DCache.scala 68:22]
  reg  valid_33_1; // @[DCache.scala 68:22]
  reg  valid_34_0; // @[DCache.scala 68:22]
  reg  valid_34_1; // @[DCache.scala 68:22]
  reg  valid_35_0; // @[DCache.scala 68:22]
  reg  valid_35_1; // @[DCache.scala 68:22]
  reg  valid_36_0; // @[DCache.scala 68:22]
  reg  valid_36_1; // @[DCache.scala 68:22]
  reg  valid_37_0; // @[DCache.scala 68:22]
  reg  valid_37_1; // @[DCache.scala 68:22]
  reg  valid_38_0; // @[DCache.scala 68:22]
  reg  valid_38_1; // @[DCache.scala 68:22]
  reg  valid_39_0; // @[DCache.scala 68:22]
  reg  valid_39_1; // @[DCache.scala 68:22]
  reg  valid_40_0; // @[DCache.scala 68:22]
  reg  valid_40_1; // @[DCache.scala 68:22]
  reg  valid_41_0; // @[DCache.scala 68:22]
  reg  valid_41_1; // @[DCache.scala 68:22]
  reg  valid_42_0; // @[DCache.scala 68:22]
  reg  valid_42_1; // @[DCache.scala 68:22]
  reg  valid_43_0; // @[DCache.scala 68:22]
  reg  valid_43_1; // @[DCache.scala 68:22]
  reg  valid_44_0; // @[DCache.scala 68:22]
  reg  valid_44_1; // @[DCache.scala 68:22]
  reg  valid_45_0; // @[DCache.scala 68:22]
  reg  valid_45_1; // @[DCache.scala 68:22]
  reg  valid_46_0; // @[DCache.scala 68:22]
  reg  valid_46_1; // @[DCache.scala 68:22]
  reg  valid_47_0; // @[DCache.scala 68:22]
  reg  valid_47_1; // @[DCache.scala 68:22]
  reg  valid_48_0; // @[DCache.scala 68:22]
  reg  valid_48_1; // @[DCache.scala 68:22]
  reg  valid_49_0; // @[DCache.scala 68:22]
  reg  valid_49_1; // @[DCache.scala 68:22]
  reg  valid_50_0; // @[DCache.scala 68:22]
  reg  valid_50_1; // @[DCache.scala 68:22]
  reg  valid_51_0; // @[DCache.scala 68:22]
  reg  valid_51_1; // @[DCache.scala 68:22]
  reg  valid_52_0; // @[DCache.scala 68:22]
  reg  valid_52_1; // @[DCache.scala 68:22]
  reg  valid_53_0; // @[DCache.scala 68:22]
  reg  valid_53_1; // @[DCache.scala 68:22]
  reg  valid_54_0; // @[DCache.scala 68:22]
  reg  valid_54_1; // @[DCache.scala 68:22]
  reg  valid_55_0; // @[DCache.scala 68:22]
  reg  valid_55_1; // @[DCache.scala 68:22]
  reg  valid_56_0; // @[DCache.scala 68:22]
  reg  valid_56_1; // @[DCache.scala 68:22]
  reg  valid_57_0; // @[DCache.scala 68:22]
  reg  valid_57_1; // @[DCache.scala 68:22]
  reg  valid_58_0; // @[DCache.scala 68:22]
  reg  valid_58_1; // @[DCache.scala 68:22]
  reg  valid_59_0; // @[DCache.scala 68:22]
  reg  valid_59_1; // @[DCache.scala 68:22]
  reg  valid_60_0; // @[DCache.scala 68:22]
  reg  valid_60_1; // @[DCache.scala 68:22]
  reg  valid_61_0; // @[DCache.scala 68:22]
  reg  valid_61_1; // @[DCache.scala 68:22]
  reg  valid_62_0; // @[DCache.scala 68:22]
  reg  valid_62_1; // @[DCache.scala 68:22]
  reg  valid_63_0; // @[DCache.scala 68:22]
  reg  valid_63_1; // @[DCache.scala 68:22]
  reg  valid_64_0; // @[DCache.scala 68:22]
  reg  valid_64_1; // @[DCache.scala 68:22]
  reg  valid_65_0; // @[DCache.scala 68:22]
  reg  valid_65_1; // @[DCache.scala 68:22]
  reg  valid_66_0; // @[DCache.scala 68:22]
  reg  valid_66_1; // @[DCache.scala 68:22]
  reg  valid_67_0; // @[DCache.scala 68:22]
  reg  valid_67_1; // @[DCache.scala 68:22]
  reg  valid_68_0; // @[DCache.scala 68:22]
  reg  valid_68_1; // @[DCache.scala 68:22]
  reg  valid_69_0; // @[DCache.scala 68:22]
  reg  valid_69_1; // @[DCache.scala 68:22]
  reg  valid_70_0; // @[DCache.scala 68:22]
  reg  valid_70_1; // @[DCache.scala 68:22]
  reg  valid_71_0; // @[DCache.scala 68:22]
  reg  valid_71_1; // @[DCache.scala 68:22]
  reg  valid_72_0; // @[DCache.scala 68:22]
  reg  valid_72_1; // @[DCache.scala 68:22]
  reg  valid_73_0; // @[DCache.scala 68:22]
  reg  valid_73_1; // @[DCache.scala 68:22]
  reg  valid_74_0; // @[DCache.scala 68:22]
  reg  valid_74_1; // @[DCache.scala 68:22]
  reg  valid_75_0; // @[DCache.scala 68:22]
  reg  valid_75_1; // @[DCache.scala 68:22]
  reg  valid_76_0; // @[DCache.scala 68:22]
  reg  valid_76_1; // @[DCache.scala 68:22]
  reg  valid_77_0; // @[DCache.scala 68:22]
  reg  valid_77_1; // @[DCache.scala 68:22]
  reg  valid_78_0; // @[DCache.scala 68:22]
  reg  valid_78_1; // @[DCache.scala 68:22]
  reg  valid_79_0; // @[DCache.scala 68:22]
  reg  valid_79_1; // @[DCache.scala 68:22]
  reg  valid_80_0; // @[DCache.scala 68:22]
  reg  valid_80_1; // @[DCache.scala 68:22]
  reg  valid_81_0; // @[DCache.scala 68:22]
  reg  valid_81_1; // @[DCache.scala 68:22]
  reg  valid_82_0; // @[DCache.scala 68:22]
  reg  valid_82_1; // @[DCache.scala 68:22]
  reg  valid_83_0; // @[DCache.scala 68:22]
  reg  valid_83_1; // @[DCache.scala 68:22]
  reg  valid_84_0; // @[DCache.scala 68:22]
  reg  valid_84_1; // @[DCache.scala 68:22]
  reg  valid_85_0; // @[DCache.scala 68:22]
  reg  valid_85_1; // @[DCache.scala 68:22]
  reg  valid_86_0; // @[DCache.scala 68:22]
  reg  valid_86_1; // @[DCache.scala 68:22]
  reg  valid_87_0; // @[DCache.scala 68:22]
  reg  valid_87_1; // @[DCache.scala 68:22]
  reg  valid_88_0; // @[DCache.scala 68:22]
  reg  valid_88_1; // @[DCache.scala 68:22]
  reg  valid_89_0; // @[DCache.scala 68:22]
  reg  valid_89_1; // @[DCache.scala 68:22]
  reg  valid_90_0; // @[DCache.scala 68:22]
  reg  valid_90_1; // @[DCache.scala 68:22]
  reg  valid_91_0; // @[DCache.scala 68:22]
  reg  valid_91_1; // @[DCache.scala 68:22]
  reg  valid_92_0; // @[DCache.scala 68:22]
  reg  valid_92_1; // @[DCache.scala 68:22]
  reg  valid_93_0; // @[DCache.scala 68:22]
  reg  valid_93_1; // @[DCache.scala 68:22]
  reg  valid_94_0; // @[DCache.scala 68:22]
  reg  valid_94_1; // @[DCache.scala 68:22]
  reg  valid_95_0; // @[DCache.scala 68:22]
  reg  valid_95_1; // @[DCache.scala 68:22]
  reg  valid_96_0; // @[DCache.scala 68:22]
  reg  valid_96_1; // @[DCache.scala 68:22]
  reg  valid_97_0; // @[DCache.scala 68:22]
  reg  valid_97_1; // @[DCache.scala 68:22]
  reg  valid_98_0; // @[DCache.scala 68:22]
  reg  valid_98_1; // @[DCache.scala 68:22]
  reg  valid_99_0; // @[DCache.scala 68:22]
  reg  valid_99_1; // @[DCache.scala 68:22]
  reg  valid_100_0; // @[DCache.scala 68:22]
  reg  valid_100_1; // @[DCache.scala 68:22]
  reg  valid_101_0; // @[DCache.scala 68:22]
  reg  valid_101_1; // @[DCache.scala 68:22]
  reg  valid_102_0; // @[DCache.scala 68:22]
  reg  valid_102_1; // @[DCache.scala 68:22]
  reg  valid_103_0; // @[DCache.scala 68:22]
  reg  valid_103_1; // @[DCache.scala 68:22]
  reg  valid_104_0; // @[DCache.scala 68:22]
  reg  valid_104_1; // @[DCache.scala 68:22]
  reg  valid_105_0; // @[DCache.scala 68:22]
  reg  valid_105_1; // @[DCache.scala 68:22]
  reg  valid_106_0; // @[DCache.scala 68:22]
  reg  valid_106_1; // @[DCache.scala 68:22]
  reg  valid_107_0; // @[DCache.scala 68:22]
  reg  valid_107_1; // @[DCache.scala 68:22]
  reg  valid_108_0; // @[DCache.scala 68:22]
  reg  valid_108_1; // @[DCache.scala 68:22]
  reg  valid_109_0; // @[DCache.scala 68:22]
  reg  valid_109_1; // @[DCache.scala 68:22]
  reg  valid_110_0; // @[DCache.scala 68:22]
  reg  valid_110_1; // @[DCache.scala 68:22]
  reg  valid_111_0; // @[DCache.scala 68:22]
  reg  valid_111_1; // @[DCache.scala 68:22]
  reg  valid_112_0; // @[DCache.scala 68:22]
  reg  valid_112_1; // @[DCache.scala 68:22]
  reg  valid_113_0; // @[DCache.scala 68:22]
  reg  valid_113_1; // @[DCache.scala 68:22]
  reg  valid_114_0; // @[DCache.scala 68:22]
  reg  valid_114_1; // @[DCache.scala 68:22]
  reg  valid_115_0; // @[DCache.scala 68:22]
  reg  valid_115_1; // @[DCache.scala 68:22]
  reg  valid_116_0; // @[DCache.scala 68:22]
  reg  valid_116_1; // @[DCache.scala 68:22]
  reg  valid_117_0; // @[DCache.scala 68:22]
  reg  valid_117_1; // @[DCache.scala 68:22]
  reg  valid_118_0; // @[DCache.scala 68:22]
  reg  valid_118_1; // @[DCache.scala 68:22]
  reg  valid_119_0; // @[DCache.scala 68:22]
  reg  valid_119_1; // @[DCache.scala 68:22]
  reg  valid_120_0; // @[DCache.scala 68:22]
  reg  valid_120_1; // @[DCache.scala 68:22]
  reg  valid_121_0; // @[DCache.scala 68:22]
  reg  valid_121_1; // @[DCache.scala 68:22]
  reg  valid_122_0; // @[DCache.scala 68:22]
  reg  valid_122_1; // @[DCache.scala 68:22]
  reg  valid_123_0; // @[DCache.scala 68:22]
  reg  valid_123_1; // @[DCache.scala 68:22]
  reg  valid_124_0; // @[DCache.scala 68:22]
  reg  valid_124_1; // @[DCache.scala 68:22]
  reg  valid_125_0; // @[DCache.scala 68:22]
  reg  valid_125_1; // @[DCache.scala 68:22]
  reg  valid_126_0; // @[DCache.scala 68:22]
  reg  valid_126_1; // @[DCache.scala 68:22]
  reg  valid_127_0; // @[DCache.scala 68:22]
  reg  valid_127_1; // @[DCache.scala 68:22]
  reg  dirty_0_0; // @[DCache.scala 69:22]
  reg  dirty_0_1; // @[DCache.scala 69:22]
  reg  dirty_1_0; // @[DCache.scala 69:22]
  reg  dirty_1_1; // @[DCache.scala 69:22]
  reg  dirty_2_0; // @[DCache.scala 69:22]
  reg  dirty_2_1; // @[DCache.scala 69:22]
  reg  dirty_3_0; // @[DCache.scala 69:22]
  reg  dirty_3_1; // @[DCache.scala 69:22]
  reg  dirty_4_0; // @[DCache.scala 69:22]
  reg  dirty_4_1; // @[DCache.scala 69:22]
  reg  dirty_5_0; // @[DCache.scala 69:22]
  reg  dirty_5_1; // @[DCache.scala 69:22]
  reg  dirty_6_0; // @[DCache.scala 69:22]
  reg  dirty_6_1; // @[DCache.scala 69:22]
  reg  dirty_7_0; // @[DCache.scala 69:22]
  reg  dirty_7_1; // @[DCache.scala 69:22]
  reg  dirty_8_0; // @[DCache.scala 69:22]
  reg  dirty_8_1; // @[DCache.scala 69:22]
  reg  dirty_9_0; // @[DCache.scala 69:22]
  reg  dirty_9_1; // @[DCache.scala 69:22]
  reg  dirty_10_0; // @[DCache.scala 69:22]
  reg  dirty_10_1; // @[DCache.scala 69:22]
  reg  dirty_11_0; // @[DCache.scala 69:22]
  reg  dirty_11_1; // @[DCache.scala 69:22]
  reg  dirty_12_0; // @[DCache.scala 69:22]
  reg  dirty_12_1; // @[DCache.scala 69:22]
  reg  dirty_13_0; // @[DCache.scala 69:22]
  reg  dirty_13_1; // @[DCache.scala 69:22]
  reg  dirty_14_0; // @[DCache.scala 69:22]
  reg  dirty_14_1; // @[DCache.scala 69:22]
  reg  dirty_15_0; // @[DCache.scala 69:22]
  reg  dirty_15_1; // @[DCache.scala 69:22]
  reg  dirty_16_0; // @[DCache.scala 69:22]
  reg  dirty_16_1; // @[DCache.scala 69:22]
  reg  dirty_17_0; // @[DCache.scala 69:22]
  reg  dirty_17_1; // @[DCache.scala 69:22]
  reg  dirty_18_0; // @[DCache.scala 69:22]
  reg  dirty_18_1; // @[DCache.scala 69:22]
  reg  dirty_19_0; // @[DCache.scala 69:22]
  reg  dirty_19_1; // @[DCache.scala 69:22]
  reg  dirty_20_0; // @[DCache.scala 69:22]
  reg  dirty_20_1; // @[DCache.scala 69:22]
  reg  dirty_21_0; // @[DCache.scala 69:22]
  reg  dirty_21_1; // @[DCache.scala 69:22]
  reg  dirty_22_0; // @[DCache.scala 69:22]
  reg  dirty_22_1; // @[DCache.scala 69:22]
  reg  dirty_23_0; // @[DCache.scala 69:22]
  reg  dirty_23_1; // @[DCache.scala 69:22]
  reg  dirty_24_0; // @[DCache.scala 69:22]
  reg  dirty_24_1; // @[DCache.scala 69:22]
  reg  dirty_25_0; // @[DCache.scala 69:22]
  reg  dirty_25_1; // @[DCache.scala 69:22]
  reg  dirty_26_0; // @[DCache.scala 69:22]
  reg  dirty_26_1; // @[DCache.scala 69:22]
  reg  dirty_27_0; // @[DCache.scala 69:22]
  reg  dirty_27_1; // @[DCache.scala 69:22]
  reg  dirty_28_0; // @[DCache.scala 69:22]
  reg  dirty_28_1; // @[DCache.scala 69:22]
  reg  dirty_29_0; // @[DCache.scala 69:22]
  reg  dirty_29_1; // @[DCache.scala 69:22]
  reg  dirty_30_0; // @[DCache.scala 69:22]
  reg  dirty_30_1; // @[DCache.scala 69:22]
  reg  dirty_31_0; // @[DCache.scala 69:22]
  reg  dirty_31_1; // @[DCache.scala 69:22]
  reg  dirty_32_0; // @[DCache.scala 69:22]
  reg  dirty_32_1; // @[DCache.scala 69:22]
  reg  dirty_33_0; // @[DCache.scala 69:22]
  reg  dirty_33_1; // @[DCache.scala 69:22]
  reg  dirty_34_0; // @[DCache.scala 69:22]
  reg  dirty_34_1; // @[DCache.scala 69:22]
  reg  dirty_35_0; // @[DCache.scala 69:22]
  reg  dirty_35_1; // @[DCache.scala 69:22]
  reg  dirty_36_0; // @[DCache.scala 69:22]
  reg  dirty_36_1; // @[DCache.scala 69:22]
  reg  dirty_37_0; // @[DCache.scala 69:22]
  reg  dirty_37_1; // @[DCache.scala 69:22]
  reg  dirty_38_0; // @[DCache.scala 69:22]
  reg  dirty_38_1; // @[DCache.scala 69:22]
  reg  dirty_39_0; // @[DCache.scala 69:22]
  reg  dirty_39_1; // @[DCache.scala 69:22]
  reg  dirty_40_0; // @[DCache.scala 69:22]
  reg  dirty_40_1; // @[DCache.scala 69:22]
  reg  dirty_41_0; // @[DCache.scala 69:22]
  reg  dirty_41_1; // @[DCache.scala 69:22]
  reg  dirty_42_0; // @[DCache.scala 69:22]
  reg  dirty_42_1; // @[DCache.scala 69:22]
  reg  dirty_43_0; // @[DCache.scala 69:22]
  reg  dirty_43_1; // @[DCache.scala 69:22]
  reg  dirty_44_0; // @[DCache.scala 69:22]
  reg  dirty_44_1; // @[DCache.scala 69:22]
  reg  dirty_45_0; // @[DCache.scala 69:22]
  reg  dirty_45_1; // @[DCache.scala 69:22]
  reg  dirty_46_0; // @[DCache.scala 69:22]
  reg  dirty_46_1; // @[DCache.scala 69:22]
  reg  dirty_47_0; // @[DCache.scala 69:22]
  reg  dirty_47_1; // @[DCache.scala 69:22]
  reg  dirty_48_0; // @[DCache.scala 69:22]
  reg  dirty_48_1; // @[DCache.scala 69:22]
  reg  dirty_49_0; // @[DCache.scala 69:22]
  reg  dirty_49_1; // @[DCache.scala 69:22]
  reg  dirty_50_0; // @[DCache.scala 69:22]
  reg  dirty_50_1; // @[DCache.scala 69:22]
  reg  dirty_51_0; // @[DCache.scala 69:22]
  reg  dirty_51_1; // @[DCache.scala 69:22]
  reg  dirty_52_0; // @[DCache.scala 69:22]
  reg  dirty_52_1; // @[DCache.scala 69:22]
  reg  dirty_53_0; // @[DCache.scala 69:22]
  reg  dirty_53_1; // @[DCache.scala 69:22]
  reg  dirty_54_0; // @[DCache.scala 69:22]
  reg  dirty_54_1; // @[DCache.scala 69:22]
  reg  dirty_55_0; // @[DCache.scala 69:22]
  reg  dirty_55_1; // @[DCache.scala 69:22]
  reg  dirty_56_0; // @[DCache.scala 69:22]
  reg  dirty_56_1; // @[DCache.scala 69:22]
  reg  dirty_57_0; // @[DCache.scala 69:22]
  reg  dirty_57_1; // @[DCache.scala 69:22]
  reg  dirty_58_0; // @[DCache.scala 69:22]
  reg  dirty_58_1; // @[DCache.scala 69:22]
  reg  dirty_59_0; // @[DCache.scala 69:22]
  reg  dirty_59_1; // @[DCache.scala 69:22]
  reg  dirty_60_0; // @[DCache.scala 69:22]
  reg  dirty_60_1; // @[DCache.scala 69:22]
  reg  dirty_61_0; // @[DCache.scala 69:22]
  reg  dirty_61_1; // @[DCache.scala 69:22]
  reg  dirty_62_0; // @[DCache.scala 69:22]
  reg  dirty_62_1; // @[DCache.scala 69:22]
  reg  dirty_63_0; // @[DCache.scala 69:22]
  reg  dirty_63_1; // @[DCache.scala 69:22]
  reg  dirty_64_0; // @[DCache.scala 69:22]
  reg  dirty_64_1; // @[DCache.scala 69:22]
  reg  dirty_65_0; // @[DCache.scala 69:22]
  reg  dirty_65_1; // @[DCache.scala 69:22]
  reg  dirty_66_0; // @[DCache.scala 69:22]
  reg  dirty_66_1; // @[DCache.scala 69:22]
  reg  dirty_67_0; // @[DCache.scala 69:22]
  reg  dirty_67_1; // @[DCache.scala 69:22]
  reg  dirty_68_0; // @[DCache.scala 69:22]
  reg  dirty_68_1; // @[DCache.scala 69:22]
  reg  dirty_69_0; // @[DCache.scala 69:22]
  reg  dirty_69_1; // @[DCache.scala 69:22]
  reg  dirty_70_0; // @[DCache.scala 69:22]
  reg  dirty_70_1; // @[DCache.scala 69:22]
  reg  dirty_71_0; // @[DCache.scala 69:22]
  reg  dirty_71_1; // @[DCache.scala 69:22]
  reg  dirty_72_0; // @[DCache.scala 69:22]
  reg  dirty_72_1; // @[DCache.scala 69:22]
  reg  dirty_73_0; // @[DCache.scala 69:22]
  reg  dirty_73_1; // @[DCache.scala 69:22]
  reg  dirty_74_0; // @[DCache.scala 69:22]
  reg  dirty_74_1; // @[DCache.scala 69:22]
  reg  dirty_75_0; // @[DCache.scala 69:22]
  reg  dirty_75_1; // @[DCache.scala 69:22]
  reg  dirty_76_0; // @[DCache.scala 69:22]
  reg  dirty_76_1; // @[DCache.scala 69:22]
  reg  dirty_77_0; // @[DCache.scala 69:22]
  reg  dirty_77_1; // @[DCache.scala 69:22]
  reg  dirty_78_0; // @[DCache.scala 69:22]
  reg  dirty_78_1; // @[DCache.scala 69:22]
  reg  dirty_79_0; // @[DCache.scala 69:22]
  reg  dirty_79_1; // @[DCache.scala 69:22]
  reg  dirty_80_0; // @[DCache.scala 69:22]
  reg  dirty_80_1; // @[DCache.scala 69:22]
  reg  dirty_81_0; // @[DCache.scala 69:22]
  reg  dirty_81_1; // @[DCache.scala 69:22]
  reg  dirty_82_0; // @[DCache.scala 69:22]
  reg  dirty_82_1; // @[DCache.scala 69:22]
  reg  dirty_83_0; // @[DCache.scala 69:22]
  reg  dirty_83_1; // @[DCache.scala 69:22]
  reg  dirty_84_0; // @[DCache.scala 69:22]
  reg  dirty_84_1; // @[DCache.scala 69:22]
  reg  dirty_85_0; // @[DCache.scala 69:22]
  reg  dirty_85_1; // @[DCache.scala 69:22]
  reg  dirty_86_0; // @[DCache.scala 69:22]
  reg  dirty_86_1; // @[DCache.scala 69:22]
  reg  dirty_87_0; // @[DCache.scala 69:22]
  reg  dirty_87_1; // @[DCache.scala 69:22]
  reg  dirty_88_0; // @[DCache.scala 69:22]
  reg  dirty_88_1; // @[DCache.scala 69:22]
  reg  dirty_89_0; // @[DCache.scala 69:22]
  reg  dirty_89_1; // @[DCache.scala 69:22]
  reg  dirty_90_0; // @[DCache.scala 69:22]
  reg  dirty_90_1; // @[DCache.scala 69:22]
  reg  dirty_91_0; // @[DCache.scala 69:22]
  reg  dirty_91_1; // @[DCache.scala 69:22]
  reg  dirty_92_0; // @[DCache.scala 69:22]
  reg  dirty_92_1; // @[DCache.scala 69:22]
  reg  dirty_93_0; // @[DCache.scala 69:22]
  reg  dirty_93_1; // @[DCache.scala 69:22]
  reg  dirty_94_0; // @[DCache.scala 69:22]
  reg  dirty_94_1; // @[DCache.scala 69:22]
  reg  dirty_95_0; // @[DCache.scala 69:22]
  reg  dirty_95_1; // @[DCache.scala 69:22]
  reg  dirty_96_0; // @[DCache.scala 69:22]
  reg  dirty_96_1; // @[DCache.scala 69:22]
  reg  dirty_97_0; // @[DCache.scala 69:22]
  reg  dirty_97_1; // @[DCache.scala 69:22]
  reg  dirty_98_0; // @[DCache.scala 69:22]
  reg  dirty_98_1; // @[DCache.scala 69:22]
  reg  dirty_99_0; // @[DCache.scala 69:22]
  reg  dirty_99_1; // @[DCache.scala 69:22]
  reg  dirty_100_0; // @[DCache.scala 69:22]
  reg  dirty_100_1; // @[DCache.scala 69:22]
  reg  dirty_101_0; // @[DCache.scala 69:22]
  reg  dirty_101_1; // @[DCache.scala 69:22]
  reg  dirty_102_0; // @[DCache.scala 69:22]
  reg  dirty_102_1; // @[DCache.scala 69:22]
  reg  dirty_103_0; // @[DCache.scala 69:22]
  reg  dirty_103_1; // @[DCache.scala 69:22]
  reg  dirty_104_0; // @[DCache.scala 69:22]
  reg  dirty_104_1; // @[DCache.scala 69:22]
  reg  dirty_105_0; // @[DCache.scala 69:22]
  reg  dirty_105_1; // @[DCache.scala 69:22]
  reg  dirty_106_0; // @[DCache.scala 69:22]
  reg  dirty_106_1; // @[DCache.scala 69:22]
  reg  dirty_107_0; // @[DCache.scala 69:22]
  reg  dirty_107_1; // @[DCache.scala 69:22]
  reg  dirty_108_0; // @[DCache.scala 69:22]
  reg  dirty_108_1; // @[DCache.scala 69:22]
  reg  dirty_109_0; // @[DCache.scala 69:22]
  reg  dirty_109_1; // @[DCache.scala 69:22]
  reg  dirty_110_0; // @[DCache.scala 69:22]
  reg  dirty_110_1; // @[DCache.scala 69:22]
  reg  dirty_111_0; // @[DCache.scala 69:22]
  reg  dirty_111_1; // @[DCache.scala 69:22]
  reg  dirty_112_0; // @[DCache.scala 69:22]
  reg  dirty_112_1; // @[DCache.scala 69:22]
  reg  dirty_113_0; // @[DCache.scala 69:22]
  reg  dirty_113_1; // @[DCache.scala 69:22]
  reg  dirty_114_0; // @[DCache.scala 69:22]
  reg  dirty_114_1; // @[DCache.scala 69:22]
  reg  dirty_115_0; // @[DCache.scala 69:22]
  reg  dirty_115_1; // @[DCache.scala 69:22]
  reg  dirty_116_0; // @[DCache.scala 69:22]
  reg  dirty_116_1; // @[DCache.scala 69:22]
  reg  dirty_117_0; // @[DCache.scala 69:22]
  reg  dirty_117_1; // @[DCache.scala 69:22]
  reg  dirty_118_0; // @[DCache.scala 69:22]
  reg  dirty_118_1; // @[DCache.scala 69:22]
  reg  dirty_119_0; // @[DCache.scala 69:22]
  reg  dirty_119_1; // @[DCache.scala 69:22]
  reg  dirty_120_0; // @[DCache.scala 69:22]
  reg  dirty_120_1; // @[DCache.scala 69:22]
  reg  dirty_121_0; // @[DCache.scala 69:22]
  reg  dirty_121_1; // @[DCache.scala 69:22]
  reg  dirty_122_0; // @[DCache.scala 69:22]
  reg  dirty_122_1; // @[DCache.scala 69:22]
  reg  dirty_123_0; // @[DCache.scala 69:22]
  reg  dirty_123_1; // @[DCache.scala 69:22]
  reg  dirty_124_0; // @[DCache.scala 69:22]
  reg  dirty_124_1; // @[DCache.scala 69:22]
  reg  dirty_125_0; // @[DCache.scala 69:22]
  reg  dirty_125_1; // @[DCache.scala 69:22]
  reg  dirty_126_0; // @[DCache.scala 69:22]
  reg  dirty_126_1; // @[DCache.scala 69:22]
  reg  dirty_127_0; // @[DCache.scala 69:22]
  reg  dirty_127_1; // @[DCache.scala 69:22]
  reg  lru_0; // @[DCache.scala 70:22]
  reg  lru_1; // @[DCache.scala 70:22]
  reg  lru_2; // @[DCache.scala 70:22]
  reg  lru_3; // @[DCache.scala 70:22]
  reg  lru_4; // @[DCache.scala 70:22]
  reg  lru_5; // @[DCache.scala 70:22]
  reg  lru_6; // @[DCache.scala 70:22]
  reg  lru_7; // @[DCache.scala 70:22]
  reg  lru_8; // @[DCache.scala 70:22]
  reg  lru_9; // @[DCache.scala 70:22]
  reg  lru_10; // @[DCache.scala 70:22]
  reg  lru_11; // @[DCache.scala 70:22]
  reg  lru_12; // @[DCache.scala 70:22]
  reg  lru_13; // @[DCache.scala 70:22]
  reg  lru_14; // @[DCache.scala 70:22]
  reg  lru_15; // @[DCache.scala 70:22]
  reg  lru_16; // @[DCache.scala 70:22]
  reg  lru_17; // @[DCache.scala 70:22]
  reg  lru_18; // @[DCache.scala 70:22]
  reg  lru_19; // @[DCache.scala 70:22]
  reg  lru_20; // @[DCache.scala 70:22]
  reg  lru_21; // @[DCache.scala 70:22]
  reg  lru_22; // @[DCache.scala 70:22]
  reg  lru_23; // @[DCache.scala 70:22]
  reg  lru_24; // @[DCache.scala 70:22]
  reg  lru_25; // @[DCache.scala 70:22]
  reg  lru_26; // @[DCache.scala 70:22]
  reg  lru_27; // @[DCache.scala 70:22]
  reg  lru_28; // @[DCache.scala 70:22]
  reg  lru_29; // @[DCache.scala 70:22]
  reg  lru_30; // @[DCache.scala 70:22]
  reg  lru_31; // @[DCache.scala 70:22]
  reg  lru_32; // @[DCache.scala 70:22]
  reg  lru_33; // @[DCache.scala 70:22]
  reg  lru_34; // @[DCache.scala 70:22]
  reg  lru_35; // @[DCache.scala 70:22]
  reg  lru_36; // @[DCache.scala 70:22]
  reg  lru_37; // @[DCache.scala 70:22]
  reg  lru_38; // @[DCache.scala 70:22]
  reg  lru_39; // @[DCache.scala 70:22]
  reg  lru_40; // @[DCache.scala 70:22]
  reg  lru_41; // @[DCache.scala 70:22]
  reg  lru_42; // @[DCache.scala 70:22]
  reg  lru_43; // @[DCache.scala 70:22]
  reg  lru_44; // @[DCache.scala 70:22]
  reg  lru_45; // @[DCache.scala 70:22]
  reg  lru_46; // @[DCache.scala 70:22]
  reg  lru_47; // @[DCache.scala 70:22]
  reg  lru_48; // @[DCache.scala 70:22]
  reg  lru_49; // @[DCache.scala 70:22]
  reg  lru_50; // @[DCache.scala 70:22]
  reg  lru_51; // @[DCache.scala 70:22]
  reg  lru_52; // @[DCache.scala 70:22]
  reg  lru_53; // @[DCache.scala 70:22]
  reg  lru_54; // @[DCache.scala 70:22]
  reg  lru_55; // @[DCache.scala 70:22]
  reg  lru_56; // @[DCache.scala 70:22]
  reg  lru_57; // @[DCache.scala 70:22]
  reg  lru_58; // @[DCache.scala 70:22]
  reg  lru_59; // @[DCache.scala 70:22]
  reg  lru_60; // @[DCache.scala 70:22]
  reg  lru_61; // @[DCache.scala 70:22]
  reg  lru_62; // @[DCache.scala 70:22]
  reg  lru_63; // @[DCache.scala 70:22]
  reg  lru_64; // @[DCache.scala 70:22]
  reg  lru_65; // @[DCache.scala 70:22]
  reg  lru_66; // @[DCache.scala 70:22]
  reg  lru_67; // @[DCache.scala 70:22]
  reg  lru_68; // @[DCache.scala 70:22]
  reg  lru_69; // @[DCache.scala 70:22]
  reg  lru_70; // @[DCache.scala 70:22]
  reg  lru_71; // @[DCache.scala 70:22]
  reg  lru_72; // @[DCache.scala 70:22]
  reg  lru_73; // @[DCache.scala 70:22]
  reg  lru_74; // @[DCache.scala 70:22]
  reg  lru_75; // @[DCache.scala 70:22]
  reg  lru_76; // @[DCache.scala 70:22]
  reg  lru_77; // @[DCache.scala 70:22]
  reg  lru_78; // @[DCache.scala 70:22]
  reg  lru_79; // @[DCache.scala 70:22]
  reg  lru_80; // @[DCache.scala 70:22]
  reg  lru_81; // @[DCache.scala 70:22]
  reg  lru_82; // @[DCache.scala 70:22]
  reg  lru_83; // @[DCache.scala 70:22]
  reg  lru_84; // @[DCache.scala 70:22]
  reg  lru_85; // @[DCache.scala 70:22]
  reg  lru_86; // @[DCache.scala 70:22]
  reg  lru_87; // @[DCache.scala 70:22]
  reg  lru_88; // @[DCache.scala 70:22]
  reg  lru_89; // @[DCache.scala 70:22]
  reg  lru_90; // @[DCache.scala 70:22]
  reg  lru_91; // @[DCache.scala 70:22]
  reg  lru_92; // @[DCache.scala 70:22]
  reg  lru_93; // @[DCache.scala 70:22]
  reg  lru_94; // @[DCache.scala 70:22]
  reg  lru_95; // @[DCache.scala 70:22]
  reg  lru_96; // @[DCache.scala 70:22]
  reg  lru_97; // @[DCache.scala 70:22]
  reg  lru_98; // @[DCache.scala 70:22]
  reg  lru_99; // @[DCache.scala 70:22]
  reg  lru_100; // @[DCache.scala 70:22]
  reg  lru_101; // @[DCache.scala 70:22]
  reg  lru_102; // @[DCache.scala 70:22]
  reg  lru_103; // @[DCache.scala 70:22]
  reg  lru_104; // @[DCache.scala 70:22]
  reg  lru_105; // @[DCache.scala 70:22]
  reg  lru_106; // @[DCache.scala 70:22]
  reg  lru_107; // @[DCache.scala 70:22]
  reg  lru_108; // @[DCache.scala 70:22]
  reg  lru_109; // @[DCache.scala 70:22]
  reg  lru_110; // @[DCache.scala 70:22]
  reg  lru_111; // @[DCache.scala 70:22]
  reg  lru_112; // @[DCache.scala 70:22]
  reg  lru_113; // @[DCache.scala 70:22]
  reg  lru_114; // @[DCache.scala 70:22]
  reg  lru_115; // @[DCache.scala 70:22]
  reg  lru_116; // @[DCache.scala 70:22]
  reg  lru_117; // @[DCache.scala 70:22]
  reg  lru_118; // @[DCache.scala 70:22]
  reg  lru_119; // @[DCache.scala 70:22]
  reg  lru_120; // @[DCache.scala 70:22]
  reg  lru_121; // @[DCache.scala 70:22]
  reg  lru_122; // @[DCache.scala 70:22]
  reg  lru_123; // @[DCache.scala 70:22]
  reg  lru_124; // @[DCache.scala 70:22]
  reg  lru_125; // @[DCache.scala 70:22]
  reg  lru_126; // @[DCache.scala 70:22]
  reg  lru_127; // @[DCache.scala 70:22]
  reg  tag_wstrb_0; // @[DCache.scala 72:33]
  reg  tag_wstrb_1; // @[DCache.scala 72:33]
  reg [3:0] bram_replace_wea_0; // @[DCache.scala 73:33]
  reg [3:0] bram_replace_wea_1; // @[DCache.scala 73:33]
  reg [19:0] tag_wdata; // @[DCache.scala 77:26]
  wire  _bram_addr_choose_T_1 = state != 3'h5; // @[DCache.scala 80:55]
  wire  bram_addr_choose = state != 3'h0 & state != 3'h5; // @[DCache.scala 80:45]
  wire [5:0] fence_line_addr = io_cpu_M_fence_addr[11:6]; // @[DCache.scala 88:45]
  reg [3:0] axi_wcnt; // @[DCache.scala 89:40]
  reg [9:0] bram_replace_addr; // @[DCache.scala 90:40]
  reg [9:0] bram_read_ready_addr; // @[DCache.scala 91:40]
  reg [9:0] bram_replace_write_addr; // @[DCache.scala 92:40]
  reg [31:0] bram_r_buffer_0; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_1; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_2; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_3; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_4; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_5; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_6; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_7; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_8; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_9; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_10; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_11; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_12; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_13; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_14; // @[DCache.scala 94:40]
  reg [31:0] bram_r_buffer_15; // @[DCache.scala 94:40]
  reg  bram_use_replace_addr; // @[DCache.scala 95:40]
  reg  fence_working; // @[DCache.scala 97:40]
  reg  replace_working; // @[DCache.scala 98:40]
  reg  ar_handshake; // @[DCache.scala 99:40]
  reg  aw_handshake; // @[DCache.scala 100:40]
  reg  replace_writeback; // @[DCache.scala 101:40]
  wire [9:0] _data_raddr_T_2 = bram_addr_choose ? io_cpu_M_mem_va[11:2] : io_cpu_E_mem_va[11:2]; // @[DCache.scala 107:8]
  wire [5:0] _tag_raddr_T_3 = bram_addr_choose ? io_cpu_M_mem_va[11:6] : io_cpu_E_mem_va[11:6]; // @[DCache.scala 112:8]
  wire [5:0] tag_raddr = bram_use_replace_addr ? bram_replace_addr[9:4] : _tag_raddr_T_3; // @[DCache.scala 109:22]
  wire  data_bram_wdata_sel = state == 3'h4; // @[DCache.scala 116:35]
  wire [19:0] cache_tag_0 = tag_ram_io_rdata; // @[DCache.scala 120:24 166:22]
  wire  _GEN_3 = 6'h1 == io_cpu_M_mem_va[11:6] ? valid_1_0 : valid_0_0; // @[DCache.scala 173:{55,55}]
  wire  _GEN_4 = 6'h2 == io_cpu_M_mem_va[11:6] ? valid_2_0 : _GEN_3; // @[DCache.scala 173:{55,55}]
  wire  _GEN_5 = 6'h3 == io_cpu_M_mem_va[11:6] ? valid_3_0 : _GEN_4; // @[DCache.scala 173:{55,55}]
  wire  _GEN_6 = 6'h4 == io_cpu_M_mem_va[11:6] ? valid_4_0 : _GEN_5; // @[DCache.scala 173:{55,55}]
  wire  _GEN_7 = 6'h5 == io_cpu_M_mem_va[11:6] ? valid_5_0 : _GEN_6; // @[DCache.scala 173:{55,55}]
  wire  _GEN_8 = 6'h6 == io_cpu_M_mem_va[11:6] ? valid_6_0 : _GEN_7; // @[DCache.scala 173:{55,55}]
  wire  _GEN_9 = 6'h7 == io_cpu_M_mem_va[11:6] ? valid_7_0 : _GEN_8; // @[DCache.scala 173:{55,55}]
  wire  _GEN_10 = 6'h8 == io_cpu_M_mem_va[11:6] ? valid_8_0 : _GEN_9; // @[DCache.scala 173:{55,55}]
  wire  _GEN_11 = 6'h9 == io_cpu_M_mem_va[11:6] ? valid_9_0 : _GEN_10; // @[DCache.scala 173:{55,55}]
  wire  _GEN_12 = 6'ha == io_cpu_M_mem_va[11:6] ? valid_10_0 : _GEN_11; // @[DCache.scala 173:{55,55}]
  wire  _GEN_13 = 6'hb == io_cpu_M_mem_va[11:6] ? valid_11_0 : _GEN_12; // @[DCache.scala 173:{55,55}]
  wire  _GEN_14 = 6'hc == io_cpu_M_mem_va[11:6] ? valid_12_0 : _GEN_13; // @[DCache.scala 173:{55,55}]
  wire  _GEN_15 = 6'hd == io_cpu_M_mem_va[11:6] ? valid_13_0 : _GEN_14; // @[DCache.scala 173:{55,55}]
  wire  _GEN_16 = 6'he == io_cpu_M_mem_va[11:6] ? valid_14_0 : _GEN_15; // @[DCache.scala 173:{55,55}]
  wire  _GEN_17 = 6'hf == io_cpu_M_mem_va[11:6] ? valid_15_0 : _GEN_16; // @[DCache.scala 173:{55,55}]
  wire  _GEN_18 = 6'h10 == io_cpu_M_mem_va[11:6] ? valid_16_0 : _GEN_17; // @[DCache.scala 173:{55,55}]
  wire  _GEN_19 = 6'h11 == io_cpu_M_mem_va[11:6] ? valid_17_0 : _GEN_18; // @[DCache.scala 173:{55,55}]
  wire  _GEN_20 = 6'h12 == io_cpu_M_mem_va[11:6] ? valid_18_0 : _GEN_19; // @[DCache.scala 173:{55,55}]
  wire  _GEN_21 = 6'h13 == io_cpu_M_mem_va[11:6] ? valid_19_0 : _GEN_20; // @[DCache.scala 173:{55,55}]
  wire  _GEN_22 = 6'h14 == io_cpu_M_mem_va[11:6] ? valid_20_0 : _GEN_21; // @[DCache.scala 173:{55,55}]
  wire  _GEN_23 = 6'h15 == io_cpu_M_mem_va[11:6] ? valid_21_0 : _GEN_22; // @[DCache.scala 173:{55,55}]
  wire  _GEN_24 = 6'h16 == io_cpu_M_mem_va[11:6] ? valid_22_0 : _GEN_23; // @[DCache.scala 173:{55,55}]
  wire  _GEN_25 = 6'h17 == io_cpu_M_mem_va[11:6] ? valid_23_0 : _GEN_24; // @[DCache.scala 173:{55,55}]
  wire  _GEN_26 = 6'h18 == io_cpu_M_mem_va[11:6] ? valid_24_0 : _GEN_25; // @[DCache.scala 173:{55,55}]
  wire  _GEN_27 = 6'h19 == io_cpu_M_mem_va[11:6] ? valid_25_0 : _GEN_26; // @[DCache.scala 173:{55,55}]
  wire  _GEN_28 = 6'h1a == io_cpu_M_mem_va[11:6] ? valid_26_0 : _GEN_27; // @[DCache.scala 173:{55,55}]
  wire  _GEN_29 = 6'h1b == io_cpu_M_mem_va[11:6] ? valid_27_0 : _GEN_28; // @[DCache.scala 173:{55,55}]
  wire  _GEN_30 = 6'h1c == io_cpu_M_mem_va[11:6] ? valid_28_0 : _GEN_29; // @[DCache.scala 173:{55,55}]
  wire  _GEN_31 = 6'h1d == io_cpu_M_mem_va[11:6] ? valid_29_0 : _GEN_30; // @[DCache.scala 173:{55,55}]
  wire  _GEN_32 = 6'h1e == io_cpu_M_mem_va[11:6] ? valid_30_0 : _GEN_31; // @[DCache.scala 173:{55,55}]
  wire  _GEN_33 = 6'h1f == io_cpu_M_mem_va[11:6] ? valid_31_0 : _GEN_32; // @[DCache.scala 173:{55,55}]
  wire  _GEN_34 = 6'h20 == io_cpu_M_mem_va[11:6] ? valid_32_0 : _GEN_33; // @[DCache.scala 173:{55,55}]
  wire  _GEN_35 = 6'h21 == io_cpu_M_mem_va[11:6] ? valid_33_0 : _GEN_34; // @[DCache.scala 173:{55,55}]
  wire  _GEN_36 = 6'h22 == io_cpu_M_mem_va[11:6] ? valid_34_0 : _GEN_35; // @[DCache.scala 173:{55,55}]
  wire  _GEN_37 = 6'h23 == io_cpu_M_mem_va[11:6] ? valid_35_0 : _GEN_36; // @[DCache.scala 173:{55,55}]
  wire  _GEN_38 = 6'h24 == io_cpu_M_mem_va[11:6] ? valid_36_0 : _GEN_37; // @[DCache.scala 173:{55,55}]
  wire  _GEN_39 = 6'h25 == io_cpu_M_mem_va[11:6] ? valid_37_0 : _GEN_38; // @[DCache.scala 173:{55,55}]
  wire  _GEN_40 = 6'h26 == io_cpu_M_mem_va[11:6] ? valid_38_0 : _GEN_39; // @[DCache.scala 173:{55,55}]
  wire  _GEN_41 = 6'h27 == io_cpu_M_mem_va[11:6] ? valid_39_0 : _GEN_40; // @[DCache.scala 173:{55,55}]
  wire  _GEN_42 = 6'h28 == io_cpu_M_mem_va[11:6] ? valid_40_0 : _GEN_41; // @[DCache.scala 173:{55,55}]
  wire  _GEN_43 = 6'h29 == io_cpu_M_mem_va[11:6] ? valid_41_0 : _GEN_42; // @[DCache.scala 173:{55,55}]
  wire  _GEN_44 = 6'h2a == io_cpu_M_mem_va[11:6] ? valid_42_0 : _GEN_43; // @[DCache.scala 173:{55,55}]
  wire  _GEN_45 = 6'h2b == io_cpu_M_mem_va[11:6] ? valid_43_0 : _GEN_44; // @[DCache.scala 173:{55,55}]
  wire  _GEN_46 = 6'h2c == io_cpu_M_mem_va[11:6] ? valid_44_0 : _GEN_45; // @[DCache.scala 173:{55,55}]
  wire  _GEN_47 = 6'h2d == io_cpu_M_mem_va[11:6] ? valid_45_0 : _GEN_46; // @[DCache.scala 173:{55,55}]
  wire  _GEN_48 = 6'h2e == io_cpu_M_mem_va[11:6] ? valid_46_0 : _GEN_47; // @[DCache.scala 173:{55,55}]
  wire  _GEN_49 = 6'h2f == io_cpu_M_mem_va[11:6] ? valid_47_0 : _GEN_48; // @[DCache.scala 173:{55,55}]
  wire  _GEN_50 = 6'h30 == io_cpu_M_mem_va[11:6] ? valid_48_0 : _GEN_49; // @[DCache.scala 173:{55,55}]
  wire  _GEN_51 = 6'h31 == io_cpu_M_mem_va[11:6] ? valid_49_0 : _GEN_50; // @[DCache.scala 173:{55,55}]
  wire  _GEN_52 = 6'h32 == io_cpu_M_mem_va[11:6] ? valid_50_0 : _GEN_51; // @[DCache.scala 173:{55,55}]
  wire  _GEN_53 = 6'h33 == io_cpu_M_mem_va[11:6] ? valid_51_0 : _GEN_52; // @[DCache.scala 173:{55,55}]
  wire  _GEN_54 = 6'h34 == io_cpu_M_mem_va[11:6] ? valid_52_0 : _GEN_53; // @[DCache.scala 173:{55,55}]
  wire  _GEN_55 = 6'h35 == io_cpu_M_mem_va[11:6] ? valid_53_0 : _GEN_54; // @[DCache.scala 173:{55,55}]
  wire  _GEN_56 = 6'h36 == io_cpu_M_mem_va[11:6] ? valid_54_0 : _GEN_55; // @[DCache.scala 173:{55,55}]
  wire  _GEN_57 = 6'h37 == io_cpu_M_mem_va[11:6] ? valid_55_0 : _GEN_56; // @[DCache.scala 173:{55,55}]
  wire  _GEN_58 = 6'h38 == io_cpu_M_mem_va[11:6] ? valid_56_0 : _GEN_57; // @[DCache.scala 173:{55,55}]
  wire  _GEN_59 = 6'h39 == io_cpu_M_mem_va[11:6] ? valid_57_0 : _GEN_58; // @[DCache.scala 173:{55,55}]
  wire  _GEN_60 = 6'h3a == io_cpu_M_mem_va[11:6] ? valid_58_0 : _GEN_59; // @[DCache.scala 173:{55,55}]
  wire  _GEN_61 = 6'h3b == io_cpu_M_mem_va[11:6] ? valid_59_0 : _GEN_60; // @[DCache.scala 173:{55,55}]
  wire  _GEN_62 = 6'h3c == io_cpu_M_mem_va[11:6] ? valid_60_0 : _GEN_61; // @[DCache.scala 173:{55,55}]
  wire  _GEN_63 = 6'h3d == io_cpu_M_mem_va[11:6] ? valid_61_0 : _GEN_62; // @[DCache.scala 173:{55,55}]
  wire  _GEN_64 = 6'h3e == io_cpu_M_mem_va[11:6] ? valid_62_0 : _GEN_63; // @[DCache.scala 173:{55,55}]
  wire  _GEN_65 = 6'h3f == io_cpu_M_mem_va[11:6] ? valid_63_0 : _GEN_64; // @[DCache.scala 173:{55,55}]
  wire [6:0] _GEN_1731 = {{1'd0}, io_cpu_M_mem_va[11:6]}; // @[DCache.scala 173:{55,55}]
  wire  _GEN_66 = 7'h40 == _GEN_1731 ? valid_64_0 : _GEN_65; // @[DCache.scala 173:{55,55}]
  wire  _GEN_67 = 7'h41 == _GEN_1731 ? valid_65_0 : _GEN_66; // @[DCache.scala 173:{55,55}]
  wire  _GEN_68 = 7'h42 == _GEN_1731 ? valid_66_0 : _GEN_67; // @[DCache.scala 173:{55,55}]
  wire  _GEN_69 = 7'h43 == _GEN_1731 ? valid_67_0 : _GEN_68; // @[DCache.scala 173:{55,55}]
  wire  _GEN_70 = 7'h44 == _GEN_1731 ? valid_68_0 : _GEN_69; // @[DCache.scala 173:{55,55}]
  wire  _GEN_71 = 7'h45 == _GEN_1731 ? valid_69_0 : _GEN_70; // @[DCache.scala 173:{55,55}]
  wire  _GEN_72 = 7'h46 == _GEN_1731 ? valid_70_0 : _GEN_71; // @[DCache.scala 173:{55,55}]
  wire  _GEN_73 = 7'h47 == _GEN_1731 ? valid_71_0 : _GEN_72; // @[DCache.scala 173:{55,55}]
  wire  _GEN_74 = 7'h48 == _GEN_1731 ? valid_72_0 : _GEN_73; // @[DCache.scala 173:{55,55}]
  wire  _GEN_75 = 7'h49 == _GEN_1731 ? valid_73_0 : _GEN_74; // @[DCache.scala 173:{55,55}]
  wire  _GEN_76 = 7'h4a == _GEN_1731 ? valid_74_0 : _GEN_75; // @[DCache.scala 173:{55,55}]
  wire  _GEN_77 = 7'h4b == _GEN_1731 ? valid_75_0 : _GEN_76; // @[DCache.scala 173:{55,55}]
  wire  _GEN_78 = 7'h4c == _GEN_1731 ? valid_76_0 : _GEN_77; // @[DCache.scala 173:{55,55}]
  wire  _GEN_79 = 7'h4d == _GEN_1731 ? valid_77_0 : _GEN_78; // @[DCache.scala 173:{55,55}]
  wire  _GEN_80 = 7'h4e == _GEN_1731 ? valid_78_0 : _GEN_79; // @[DCache.scala 173:{55,55}]
  wire  _GEN_81 = 7'h4f == _GEN_1731 ? valid_79_0 : _GEN_80; // @[DCache.scala 173:{55,55}]
  wire  _GEN_82 = 7'h50 == _GEN_1731 ? valid_80_0 : _GEN_81; // @[DCache.scala 173:{55,55}]
  wire  _GEN_83 = 7'h51 == _GEN_1731 ? valid_81_0 : _GEN_82; // @[DCache.scala 173:{55,55}]
  wire  _GEN_84 = 7'h52 == _GEN_1731 ? valid_82_0 : _GEN_83; // @[DCache.scala 173:{55,55}]
  wire  _GEN_85 = 7'h53 == _GEN_1731 ? valid_83_0 : _GEN_84; // @[DCache.scala 173:{55,55}]
  wire  _GEN_86 = 7'h54 == _GEN_1731 ? valid_84_0 : _GEN_85; // @[DCache.scala 173:{55,55}]
  wire  _GEN_87 = 7'h55 == _GEN_1731 ? valid_85_0 : _GEN_86; // @[DCache.scala 173:{55,55}]
  wire  _GEN_88 = 7'h56 == _GEN_1731 ? valid_86_0 : _GEN_87; // @[DCache.scala 173:{55,55}]
  wire  _GEN_89 = 7'h57 == _GEN_1731 ? valid_87_0 : _GEN_88; // @[DCache.scala 173:{55,55}]
  wire  _GEN_90 = 7'h58 == _GEN_1731 ? valid_88_0 : _GEN_89; // @[DCache.scala 173:{55,55}]
  wire  _GEN_91 = 7'h59 == _GEN_1731 ? valid_89_0 : _GEN_90; // @[DCache.scala 173:{55,55}]
  wire  _GEN_92 = 7'h5a == _GEN_1731 ? valid_90_0 : _GEN_91; // @[DCache.scala 173:{55,55}]
  wire  _GEN_93 = 7'h5b == _GEN_1731 ? valid_91_0 : _GEN_92; // @[DCache.scala 173:{55,55}]
  wire  _GEN_94 = 7'h5c == _GEN_1731 ? valid_92_0 : _GEN_93; // @[DCache.scala 173:{55,55}]
  wire  _GEN_95 = 7'h5d == _GEN_1731 ? valid_93_0 : _GEN_94; // @[DCache.scala 173:{55,55}]
  wire  _GEN_96 = 7'h5e == _GEN_1731 ? valid_94_0 : _GEN_95; // @[DCache.scala 173:{55,55}]
  wire  _GEN_97 = 7'h5f == _GEN_1731 ? valid_95_0 : _GEN_96; // @[DCache.scala 173:{55,55}]
  wire  _GEN_98 = 7'h60 == _GEN_1731 ? valid_96_0 : _GEN_97; // @[DCache.scala 173:{55,55}]
  wire  _GEN_99 = 7'h61 == _GEN_1731 ? valid_97_0 : _GEN_98; // @[DCache.scala 173:{55,55}]
  wire  _GEN_100 = 7'h62 == _GEN_1731 ? valid_98_0 : _GEN_99; // @[DCache.scala 173:{55,55}]
  wire  _GEN_101 = 7'h63 == _GEN_1731 ? valid_99_0 : _GEN_100; // @[DCache.scala 173:{55,55}]
  wire  _GEN_102 = 7'h64 == _GEN_1731 ? valid_100_0 : _GEN_101; // @[DCache.scala 173:{55,55}]
  wire  _GEN_103 = 7'h65 == _GEN_1731 ? valid_101_0 : _GEN_102; // @[DCache.scala 173:{55,55}]
  wire  _GEN_104 = 7'h66 == _GEN_1731 ? valid_102_0 : _GEN_103; // @[DCache.scala 173:{55,55}]
  wire  _GEN_105 = 7'h67 == _GEN_1731 ? valid_103_0 : _GEN_104; // @[DCache.scala 173:{55,55}]
  wire  _GEN_106 = 7'h68 == _GEN_1731 ? valid_104_0 : _GEN_105; // @[DCache.scala 173:{55,55}]
  wire  _GEN_107 = 7'h69 == _GEN_1731 ? valid_105_0 : _GEN_106; // @[DCache.scala 173:{55,55}]
  wire  _GEN_108 = 7'h6a == _GEN_1731 ? valid_106_0 : _GEN_107; // @[DCache.scala 173:{55,55}]
  wire  _GEN_109 = 7'h6b == _GEN_1731 ? valid_107_0 : _GEN_108; // @[DCache.scala 173:{55,55}]
  wire  _GEN_110 = 7'h6c == _GEN_1731 ? valid_108_0 : _GEN_109; // @[DCache.scala 173:{55,55}]
  wire  _GEN_111 = 7'h6d == _GEN_1731 ? valid_109_0 : _GEN_110; // @[DCache.scala 173:{55,55}]
  wire  _GEN_112 = 7'h6e == _GEN_1731 ? valid_110_0 : _GEN_111; // @[DCache.scala 173:{55,55}]
  wire  _GEN_113 = 7'h6f == _GEN_1731 ? valid_111_0 : _GEN_112; // @[DCache.scala 173:{55,55}]
  wire  _GEN_114 = 7'h70 == _GEN_1731 ? valid_112_0 : _GEN_113; // @[DCache.scala 173:{55,55}]
  wire  _GEN_115 = 7'h71 == _GEN_1731 ? valid_113_0 : _GEN_114; // @[DCache.scala 173:{55,55}]
  wire  _GEN_116 = 7'h72 == _GEN_1731 ? valid_114_0 : _GEN_115; // @[DCache.scala 173:{55,55}]
  wire  _GEN_117 = 7'h73 == _GEN_1731 ? valid_115_0 : _GEN_116; // @[DCache.scala 173:{55,55}]
  wire  _GEN_118 = 7'h74 == _GEN_1731 ? valid_116_0 : _GEN_117; // @[DCache.scala 173:{55,55}]
  wire  _GEN_119 = 7'h75 == _GEN_1731 ? valid_117_0 : _GEN_118; // @[DCache.scala 173:{55,55}]
  wire  _GEN_120 = 7'h76 == _GEN_1731 ? valid_118_0 : _GEN_119; // @[DCache.scala 173:{55,55}]
  wire  _GEN_121 = 7'h77 == _GEN_1731 ? valid_119_0 : _GEN_120; // @[DCache.scala 173:{55,55}]
  wire  _GEN_122 = 7'h78 == _GEN_1731 ? valid_120_0 : _GEN_121; // @[DCache.scala 173:{55,55}]
  wire  _GEN_123 = 7'h79 == _GEN_1731 ? valid_121_0 : _GEN_122; // @[DCache.scala 173:{55,55}]
  wire  _GEN_124 = 7'h7a == _GEN_1731 ? valid_122_0 : _GEN_123; // @[DCache.scala 173:{55,55}]
  wire  _GEN_125 = 7'h7b == _GEN_1731 ? valid_123_0 : _GEN_124; // @[DCache.scala 173:{55,55}]
  wire  _GEN_126 = 7'h7c == _GEN_1731 ? valid_124_0 : _GEN_125; // @[DCache.scala 173:{55,55}]
  wire  _GEN_127 = 7'h7d == _GEN_1731 ? valid_125_0 : _GEN_126; // @[DCache.scala 173:{55,55}]
  wire  _GEN_128 = 7'h7e == _GEN_1731 ? valid_126_0 : _GEN_127; // @[DCache.scala 173:{55,55}]
  wire  _GEN_129 = 7'h7f == _GEN_1731 ? valid_127_0 : _GEN_128; // @[DCache.scala 173:{55,55}]
  wire  tag_compare_valid_0 = cache_tag_0 == data_tag & _GEN_129 & translation_ok; // @[DCache.scala 173:81]
  wire [19:0] cache_tag_1 = tag_ram_1_io_rdata; // @[DCache.scala 120:24 166:22]
  wire  _GEN_131 = 6'h1 == io_cpu_M_mem_va[11:6] ? valid_1_1 : valid_0_1; // @[DCache.scala 173:{55,55}]
  wire  _GEN_132 = 6'h2 == io_cpu_M_mem_va[11:6] ? valid_2_1 : _GEN_131; // @[DCache.scala 173:{55,55}]
  wire  _GEN_133 = 6'h3 == io_cpu_M_mem_va[11:6] ? valid_3_1 : _GEN_132; // @[DCache.scala 173:{55,55}]
  wire  _GEN_134 = 6'h4 == io_cpu_M_mem_va[11:6] ? valid_4_1 : _GEN_133; // @[DCache.scala 173:{55,55}]
  wire  _GEN_135 = 6'h5 == io_cpu_M_mem_va[11:6] ? valid_5_1 : _GEN_134; // @[DCache.scala 173:{55,55}]
  wire  _GEN_136 = 6'h6 == io_cpu_M_mem_va[11:6] ? valid_6_1 : _GEN_135; // @[DCache.scala 173:{55,55}]
  wire  _GEN_137 = 6'h7 == io_cpu_M_mem_va[11:6] ? valid_7_1 : _GEN_136; // @[DCache.scala 173:{55,55}]
  wire  _GEN_138 = 6'h8 == io_cpu_M_mem_va[11:6] ? valid_8_1 : _GEN_137; // @[DCache.scala 173:{55,55}]
  wire  _GEN_139 = 6'h9 == io_cpu_M_mem_va[11:6] ? valid_9_1 : _GEN_138; // @[DCache.scala 173:{55,55}]
  wire  _GEN_140 = 6'ha == io_cpu_M_mem_va[11:6] ? valid_10_1 : _GEN_139; // @[DCache.scala 173:{55,55}]
  wire  _GEN_141 = 6'hb == io_cpu_M_mem_va[11:6] ? valid_11_1 : _GEN_140; // @[DCache.scala 173:{55,55}]
  wire  _GEN_142 = 6'hc == io_cpu_M_mem_va[11:6] ? valid_12_1 : _GEN_141; // @[DCache.scala 173:{55,55}]
  wire  _GEN_143 = 6'hd == io_cpu_M_mem_va[11:6] ? valid_13_1 : _GEN_142; // @[DCache.scala 173:{55,55}]
  wire  _GEN_144 = 6'he == io_cpu_M_mem_va[11:6] ? valid_14_1 : _GEN_143; // @[DCache.scala 173:{55,55}]
  wire  _GEN_145 = 6'hf == io_cpu_M_mem_va[11:6] ? valid_15_1 : _GEN_144; // @[DCache.scala 173:{55,55}]
  wire  _GEN_146 = 6'h10 == io_cpu_M_mem_va[11:6] ? valid_16_1 : _GEN_145; // @[DCache.scala 173:{55,55}]
  wire  _GEN_147 = 6'h11 == io_cpu_M_mem_va[11:6] ? valid_17_1 : _GEN_146; // @[DCache.scala 173:{55,55}]
  wire  _GEN_148 = 6'h12 == io_cpu_M_mem_va[11:6] ? valid_18_1 : _GEN_147; // @[DCache.scala 173:{55,55}]
  wire  _GEN_149 = 6'h13 == io_cpu_M_mem_va[11:6] ? valid_19_1 : _GEN_148; // @[DCache.scala 173:{55,55}]
  wire  _GEN_150 = 6'h14 == io_cpu_M_mem_va[11:6] ? valid_20_1 : _GEN_149; // @[DCache.scala 173:{55,55}]
  wire  _GEN_151 = 6'h15 == io_cpu_M_mem_va[11:6] ? valid_21_1 : _GEN_150; // @[DCache.scala 173:{55,55}]
  wire  _GEN_152 = 6'h16 == io_cpu_M_mem_va[11:6] ? valid_22_1 : _GEN_151; // @[DCache.scala 173:{55,55}]
  wire  _GEN_153 = 6'h17 == io_cpu_M_mem_va[11:6] ? valid_23_1 : _GEN_152; // @[DCache.scala 173:{55,55}]
  wire  _GEN_154 = 6'h18 == io_cpu_M_mem_va[11:6] ? valid_24_1 : _GEN_153; // @[DCache.scala 173:{55,55}]
  wire  _GEN_155 = 6'h19 == io_cpu_M_mem_va[11:6] ? valid_25_1 : _GEN_154; // @[DCache.scala 173:{55,55}]
  wire  _GEN_156 = 6'h1a == io_cpu_M_mem_va[11:6] ? valid_26_1 : _GEN_155; // @[DCache.scala 173:{55,55}]
  wire  _GEN_157 = 6'h1b == io_cpu_M_mem_va[11:6] ? valid_27_1 : _GEN_156; // @[DCache.scala 173:{55,55}]
  wire  _GEN_158 = 6'h1c == io_cpu_M_mem_va[11:6] ? valid_28_1 : _GEN_157; // @[DCache.scala 173:{55,55}]
  wire  _GEN_159 = 6'h1d == io_cpu_M_mem_va[11:6] ? valid_29_1 : _GEN_158; // @[DCache.scala 173:{55,55}]
  wire  _GEN_160 = 6'h1e == io_cpu_M_mem_va[11:6] ? valid_30_1 : _GEN_159; // @[DCache.scala 173:{55,55}]
  wire  _GEN_161 = 6'h1f == io_cpu_M_mem_va[11:6] ? valid_31_1 : _GEN_160; // @[DCache.scala 173:{55,55}]
  wire  _GEN_162 = 6'h20 == io_cpu_M_mem_va[11:6] ? valid_32_1 : _GEN_161; // @[DCache.scala 173:{55,55}]
  wire  _GEN_163 = 6'h21 == io_cpu_M_mem_va[11:6] ? valid_33_1 : _GEN_162; // @[DCache.scala 173:{55,55}]
  wire  _GEN_164 = 6'h22 == io_cpu_M_mem_va[11:6] ? valid_34_1 : _GEN_163; // @[DCache.scala 173:{55,55}]
  wire  _GEN_165 = 6'h23 == io_cpu_M_mem_va[11:6] ? valid_35_1 : _GEN_164; // @[DCache.scala 173:{55,55}]
  wire  _GEN_166 = 6'h24 == io_cpu_M_mem_va[11:6] ? valid_36_1 : _GEN_165; // @[DCache.scala 173:{55,55}]
  wire  _GEN_167 = 6'h25 == io_cpu_M_mem_va[11:6] ? valid_37_1 : _GEN_166; // @[DCache.scala 173:{55,55}]
  wire  _GEN_168 = 6'h26 == io_cpu_M_mem_va[11:6] ? valid_38_1 : _GEN_167; // @[DCache.scala 173:{55,55}]
  wire  _GEN_169 = 6'h27 == io_cpu_M_mem_va[11:6] ? valid_39_1 : _GEN_168; // @[DCache.scala 173:{55,55}]
  wire  _GEN_170 = 6'h28 == io_cpu_M_mem_va[11:6] ? valid_40_1 : _GEN_169; // @[DCache.scala 173:{55,55}]
  wire  _GEN_171 = 6'h29 == io_cpu_M_mem_va[11:6] ? valid_41_1 : _GEN_170; // @[DCache.scala 173:{55,55}]
  wire  _GEN_172 = 6'h2a == io_cpu_M_mem_va[11:6] ? valid_42_1 : _GEN_171; // @[DCache.scala 173:{55,55}]
  wire  _GEN_173 = 6'h2b == io_cpu_M_mem_va[11:6] ? valid_43_1 : _GEN_172; // @[DCache.scala 173:{55,55}]
  wire  _GEN_174 = 6'h2c == io_cpu_M_mem_va[11:6] ? valid_44_1 : _GEN_173; // @[DCache.scala 173:{55,55}]
  wire  _GEN_175 = 6'h2d == io_cpu_M_mem_va[11:6] ? valid_45_1 : _GEN_174; // @[DCache.scala 173:{55,55}]
  wire  _GEN_176 = 6'h2e == io_cpu_M_mem_va[11:6] ? valid_46_1 : _GEN_175; // @[DCache.scala 173:{55,55}]
  wire  _GEN_177 = 6'h2f == io_cpu_M_mem_va[11:6] ? valid_47_1 : _GEN_176; // @[DCache.scala 173:{55,55}]
  wire  _GEN_178 = 6'h30 == io_cpu_M_mem_va[11:6] ? valid_48_1 : _GEN_177; // @[DCache.scala 173:{55,55}]
  wire  _GEN_179 = 6'h31 == io_cpu_M_mem_va[11:6] ? valid_49_1 : _GEN_178; // @[DCache.scala 173:{55,55}]
  wire  _GEN_180 = 6'h32 == io_cpu_M_mem_va[11:6] ? valid_50_1 : _GEN_179; // @[DCache.scala 173:{55,55}]
  wire  _GEN_181 = 6'h33 == io_cpu_M_mem_va[11:6] ? valid_51_1 : _GEN_180; // @[DCache.scala 173:{55,55}]
  wire  _GEN_182 = 6'h34 == io_cpu_M_mem_va[11:6] ? valid_52_1 : _GEN_181; // @[DCache.scala 173:{55,55}]
  wire  _GEN_183 = 6'h35 == io_cpu_M_mem_va[11:6] ? valid_53_1 : _GEN_182; // @[DCache.scala 173:{55,55}]
  wire  _GEN_184 = 6'h36 == io_cpu_M_mem_va[11:6] ? valid_54_1 : _GEN_183; // @[DCache.scala 173:{55,55}]
  wire  _GEN_185 = 6'h37 == io_cpu_M_mem_va[11:6] ? valid_55_1 : _GEN_184; // @[DCache.scala 173:{55,55}]
  wire  _GEN_186 = 6'h38 == io_cpu_M_mem_va[11:6] ? valid_56_1 : _GEN_185; // @[DCache.scala 173:{55,55}]
  wire  _GEN_187 = 6'h39 == io_cpu_M_mem_va[11:6] ? valid_57_1 : _GEN_186; // @[DCache.scala 173:{55,55}]
  wire  _GEN_188 = 6'h3a == io_cpu_M_mem_va[11:6] ? valid_58_1 : _GEN_187; // @[DCache.scala 173:{55,55}]
  wire  _GEN_189 = 6'h3b == io_cpu_M_mem_va[11:6] ? valid_59_1 : _GEN_188; // @[DCache.scala 173:{55,55}]
  wire  _GEN_190 = 6'h3c == io_cpu_M_mem_va[11:6] ? valid_60_1 : _GEN_189; // @[DCache.scala 173:{55,55}]
  wire  _GEN_191 = 6'h3d == io_cpu_M_mem_va[11:6] ? valid_61_1 : _GEN_190; // @[DCache.scala 173:{55,55}]
  wire  _GEN_192 = 6'h3e == io_cpu_M_mem_va[11:6] ? valid_62_1 : _GEN_191; // @[DCache.scala 173:{55,55}]
  wire  _GEN_193 = 6'h3f == io_cpu_M_mem_va[11:6] ? valid_63_1 : _GEN_192; // @[DCache.scala 173:{55,55}]
  wire  _GEN_194 = 7'h40 == _GEN_1731 ? valid_64_1 : _GEN_193; // @[DCache.scala 173:{55,55}]
  wire  _GEN_195 = 7'h41 == _GEN_1731 ? valid_65_1 : _GEN_194; // @[DCache.scala 173:{55,55}]
  wire  _GEN_196 = 7'h42 == _GEN_1731 ? valid_66_1 : _GEN_195; // @[DCache.scala 173:{55,55}]
  wire  _GEN_197 = 7'h43 == _GEN_1731 ? valid_67_1 : _GEN_196; // @[DCache.scala 173:{55,55}]
  wire  _GEN_198 = 7'h44 == _GEN_1731 ? valid_68_1 : _GEN_197; // @[DCache.scala 173:{55,55}]
  wire  _GEN_199 = 7'h45 == _GEN_1731 ? valid_69_1 : _GEN_198; // @[DCache.scala 173:{55,55}]
  wire  _GEN_200 = 7'h46 == _GEN_1731 ? valid_70_1 : _GEN_199; // @[DCache.scala 173:{55,55}]
  wire  _GEN_201 = 7'h47 == _GEN_1731 ? valid_71_1 : _GEN_200; // @[DCache.scala 173:{55,55}]
  wire  _GEN_202 = 7'h48 == _GEN_1731 ? valid_72_1 : _GEN_201; // @[DCache.scala 173:{55,55}]
  wire  _GEN_203 = 7'h49 == _GEN_1731 ? valid_73_1 : _GEN_202; // @[DCache.scala 173:{55,55}]
  wire  _GEN_204 = 7'h4a == _GEN_1731 ? valid_74_1 : _GEN_203; // @[DCache.scala 173:{55,55}]
  wire  _GEN_205 = 7'h4b == _GEN_1731 ? valid_75_1 : _GEN_204; // @[DCache.scala 173:{55,55}]
  wire  _GEN_206 = 7'h4c == _GEN_1731 ? valid_76_1 : _GEN_205; // @[DCache.scala 173:{55,55}]
  wire  _GEN_207 = 7'h4d == _GEN_1731 ? valid_77_1 : _GEN_206; // @[DCache.scala 173:{55,55}]
  wire  _GEN_208 = 7'h4e == _GEN_1731 ? valid_78_1 : _GEN_207; // @[DCache.scala 173:{55,55}]
  wire  _GEN_209 = 7'h4f == _GEN_1731 ? valid_79_1 : _GEN_208; // @[DCache.scala 173:{55,55}]
  wire  _GEN_210 = 7'h50 == _GEN_1731 ? valid_80_1 : _GEN_209; // @[DCache.scala 173:{55,55}]
  wire  _GEN_211 = 7'h51 == _GEN_1731 ? valid_81_1 : _GEN_210; // @[DCache.scala 173:{55,55}]
  wire  _GEN_212 = 7'h52 == _GEN_1731 ? valid_82_1 : _GEN_211; // @[DCache.scala 173:{55,55}]
  wire  _GEN_213 = 7'h53 == _GEN_1731 ? valid_83_1 : _GEN_212; // @[DCache.scala 173:{55,55}]
  wire  _GEN_214 = 7'h54 == _GEN_1731 ? valid_84_1 : _GEN_213; // @[DCache.scala 173:{55,55}]
  wire  _GEN_215 = 7'h55 == _GEN_1731 ? valid_85_1 : _GEN_214; // @[DCache.scala 173:{55,55}]
  wire  _GEN_216 = 7'h56 == _GEN_1731 ? valid_86_1 : _GEN_215; // @[DCache.scala 173:{55,55}]
  wire  _GEN_217 = 7'h57 == _GEN_1731 ? valid_87_1 : _GEN_216; // @[DCache.scala 173:{55,55}]
  wire  _GEN_218 = 7'h58 == _GEN_1731 ? valid_88_1 : _GEN_217; // @[DCache.scala 173:{55,55}]
  wire  _GEN_219 = 7'h59 == _GEN_1731 ? valid_89_1 : _GEN_218; // @[DCache.scala 173:{55,55}]
  wire  _GEN_220 = 7'h5a == _GEN_1731 ? valid_90_1 : _GEN_219; // @[DCache.scala 173:{55,55}]
  wire  _GEN_221 = 7'h5b == _GEN_1731 ? valid_91_1 : _GEN_220; // @[DCache.scala 173:{55,55}]
  wire  _GEN_222 = 7'h5c == _GEN_1731 ? valid_92_1 : _GEN_221; // @[DCache.scala 173:{55,55}]
  wire  _GEN_223 = 7'h5d == _GEN_1731 ? valid_93_1 : _GEN_222; // @[DCache.scala 173:{55,55}]
  wire  _GEN_224 = 7'h5e == _GEN_1731 ? valid_94_1 : _GEN_223; // @[DCache.scala 173:{55,55}]
  wire  _GEN_225 = 7'h5f == _GEN_1731 ? valid_95_1 : _GEN_224; // @[DCache.scala 173:{55,55}]
  wire  _GEN_226 = 7'h60 == _GEN_1731 ? valid_96_1 : _GEN_225; // @[DCache.scala 173:{55,55}]
  wire  _GEN_227 = 7'h61 == _GEN_1731 ? valid_97_1 : _GEN_226; // @[DCache.scala 173:{55,55}]
  wire  _GEN_228 = 7'h62 == _GEN_1731 ? valid_98_1 : _GEN_227; // @[DCache.scala 173:{55,55}]
  wire  _GEN_229 = 7'h63 == _GEN_1731 ? valid_99_1 : _GEN_228; // @[DCache.scala 173:{55,55}]
  wire  _GEN_230 = 7'h64 == _GEN_1731 ? valid_100_1 : _GEN_229; // @[DCache.scala 173:{55,55}]
  wire  _GEN_231 = 7'h65 == _GEN_1731 ? valid_101_1 : _GEN_230; // @[DCache.scala 173:{55,55}]
  wire  _GEN_232 = 7'h66 == _GEN_1731 ? valid_102_1 : _GEN_231; // @[DCache.scala 173:{55,55}]
  wire  _GEN_233 = 7'h67 == _GEN_1731 ? valid_103_1 : _GEN_232; // @[DCache.scala 173:{55,55}]
  wire  _GEN_234 = 7'h68 == _GEN_1731 ? valid_104_1 : _GEN_233; // @[DCache.scala 173:{55,55}]
  wire  _GEN_235 = 7'h69 == _GEN_1731 ? valid_105_1 : _GEN_234; // @[DCache.scala 173:{55,55}]
  wire  _GEN_236 = 7'h6a == _GEN_1731 ? valid_106_1 : _GEN_235; // @[DCache.scala 173:{55,55}]
  wire  _GEN_237 = 7'h6b == _GEN_1731 ? valid_107_1 : _GEN_236; // @[DCache.scala 173:{55,55}]
  wire  _GEN_238 = 7'h6c == _GEN_1731 ? valid_108_1 : _GEN_237; // @[DCache.scala 173:{55,55}]
  wire  _GEN_239 = 7'h6d == _GEN_1731 ? valid_109_1 : _GEN_238; // @[DCache.scala 173:{55,55}]
  wire  _GEN_240 = 7'h6e == _GEN_1731 ? valid_110_1 : _GEN_239; // @[DCache.scala 173:{55,55}]
  wire  _GEN_241 = 7'h6f == _GEN_1731 ? valid_111_1 : _GEN_240; // @[DCache.scala 173:{55,55}]
  wire  _GEN_242 = 7'h70 == _GEN_1731 ? valid_112_1 : _GEN_241; // @[DCache.scala 173:{55,55}]
  wire  _GEN_243 = 7'h71 == _GEN_1731 ? valid_113_1 : _GEN_242; // @[DCache.scala 173:{55,55}]
  wire  _GEN_244 = 7'h72 == _GEN_1731 ? valid_114_1 : _GEN_243; // @[DCache.scala 173:{55,55}]
  wire  _GEN_245 = 7'h73 == _GEN_1731 ? valid_115_1 : _GEN_244; // @[DCache.scala 173:{55,55}]
  wire  _GEN_246 = 7'h74 == _GEN_1731 ? valid_116_1 : _GEN_245; // @[DCache.scala 173:{55,55}]
  wire  _GEN_247 = 7'h75 == _GEN_1731 ? valid_117_1 : _GEN_246; // @[DCache.scala 173:{55,55}]
  wire  _GEN_248 = 7'h76 == _GEN_1731 ? valid_118_1 : _GEN_247; // @[DCache.scala 173:{55,55}]
  wire  _GEN_249 = 7'h77 == _GEN_1731 ? valid_119_1 : _GEN_248; // @[DCache.scala 173:{55,55}]
  wire  _GEN_250 = 7'h78 == _GEN_1731 ? valid_120_1 : _GEN_249; // @[DCache.scala 173:{55,55}]
  wire  _GEN_251 = 7'h79 == _GEN_1731 ? valid_121_1 : _GEN_250; // @[DCache.scala 173:{55,55}]
  wire  _GEN_252 = 7'h7a == _GEN_1731 ? valid_122_1 : _GEN_251; // @[DCache.scala 173:{55,55}]
  wire  _GEN_253 = 7'h7b == _GEN_1731 ? valid_123_1 : _GEN_252; // @[DCache.scala 173:{55,55}]
  wire  _GEN_254 = 7'h7c == _GEN_1731 ? valid_124_1 : _GEN_253; // @[DCache.scala 173:{55,55}]
  wire  _GEN_255 = 7'h7d == _GEN_1731 ? valid_125_1 : _GEN_254; // @[DCache.scala 173:{55,55}]
  wire  _GEN_256 = 7'h7e == _GEN_1731 ? valid_126_1 : _GEN_255; // @[DCache.scala 173:{55,55}]
  wire  _GEN_257 = 7'h7f == _GEN_1731 ? valid_127_1 : _GEN_256; // @[DCache.scala 173:{55,55}]
  wire  tag_compare_valid_1 = cache_tag_1 == data_tag & _GEN_257 & translation_ok; // @[DCache.scala 173:81]
  wire  cache_hit = tag_compare_valid_0 | tag_compare_valid_1; // @[DCache.scala 123:53]
  wire  mmio_read_stall = M_mem_uncached & _translation_ok_T_2; // @[DCache.scala 125:41]
  wire  mmio_write_stall = M_mem_uncached & io_cpu_M_mem_write & ~write_buffer_io_enq_ready; // @[DCache.scala 126:56]
  wire  _cached_stall_T = ~M_mem_uncached; // @[DCache.scala 127:26]
  wire  _cached_stall_T_1 = ~cache_hit; // @[DCache.scala 127:45]
  wire  cached_stall = ~M_mem_uncached & ~cache_hit; // @[DCache.scala 127:42]
  wire  tlb_stall = ~translation_ok; // @[DCache.scala 128:26]
  wire  _io_cpu_dstall_T = state == 3'h0; // @[DCache.scala 136:11]
  wire  _io_cpu_dstall_T_4 = io_cpu_M_mem_en ? cached_stall | mmio_read_stall | mmio_write_stall | tlb_stall :
    io_cpu_M_fence_d; // @[DCache.scala 137:8]
  reg [31:0] saved_rdata; // @[DCache.scala 141:28]
  reg [9:0] last_line_addr; // @[DCache.scala 144:35]
  reg [31:0] last_wea_0; // @[DCache.scala 145:35]
  reg [31:0] last_wea_1; // @[DCache.scala 145:35]
  reg [31:0] last_wdata; // @[DCache.scala 146:35]
  wire  _cache_data_forward_0_T_1 = last_line_addr == io_cpu_M_mem_va[11:2]; // @[DCache.scala 175:22]
  wire [31:0] _cache_data_forward_0_T_2 = last_wea_0 & last_wdata; // @[DCache.scala 176:21]
  wire [31:0] cache_data_0 = bank_ram_io_rdata; // @[DCache.scala 119:24 156:23]
  wire [31:0] _cache_data_forward_0_T_3 = ~last_wea_0; // @[DCache.scala 176:55]
  wire [31:0] _cache_data_forward_0_T_4 = cache_data_0 & _cache_data_forward_0_T_3; // @[DCache.scala 176:52]
  wire [31:0] _cache_data_forward_0_T_5 = _cache_data_forward_0_T_2 | _cache_data_forward_0_T_4; // @[DCache.scala 176:35]
  wire [31:0] cache_data_forward_0 = _cache_data_forward_0_T_1 ? _cache_data_forward_0_T_5 : cache_data_0; // @[DCache.scala 174:33]
  wire [31:0] _cache_data_forward_1_T_2 = last_wea_1 & last_wdata; // @[DCache.scala 176:21]
  wire [31:0] cache_data_1 = bank_ram_1_io_rdata; // @[DCache.scala 119:24 156:23]
  wire [31:0] _cache_data_forward_1_T_3 = ~last_wea_1; // @[DCache.scala 176:55]
  wire [31:0] _cache_data_forward_1_T_4 = cache_data_1 & _cache_data_forward_1_T_3; // @[DCache.scala 176:52]
  wire [31:0] _cache_data_forward_1_T_5 = _cache_data_forward_1_T_2 | _cache_data_forward_1_T_4; // @[DCache.scala 176:35]
  wire [31:0] cache_data_forward_1 = _cache_data_forward_0_T_1 ? _cache_data_forward_1_T_5 : cache_data_1; // @[DCache.scala 174:33]
  wire [31:0] _GEN_1 = tag_compare_valid_1 ? cache_data_forward_1 : cache_data_forward_0; // @[DCache.scala 149:{24,24}]
  wire  _data_wstrb_0_T_5 = tag_compare_valid_0 & io_cpu_M_mem_en & io_cpu_M_mem_write & _cached_stall_T &
    _io_cpu_dstall_T; // @[DCache.scala 181:74]
  wire [3:0] data_wstrb_0 = _data_wstrb_0_T_5 ? io_cpu_M_wmask : bram_replace_wea_0; // @[DCache.scala 180:25]
  wire [7:0] _last_wea_0_T_2 = data_wstrb_0[3] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _last_wea_0_T_5 = data_wstrb_0[2] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _last_wea_0_T_8 = data_wstrb_0[1] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _last_wea_0_T_11 = data_wstrb_0[0] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _last_wea_0_T_12 = {_last_wea_0_T_2,_last_wea_0_T_5,_last_wea_0_T_8,_last_wea_0_T_11}; // @[Cat.scala 33:92]
  wire  _data_wstrb_1_T_5 = tag_compare_valid_1 & io_cpu_M_mem_en & io_cpu_M_mem_write & _cached_stall_T &
    _io_cpu_dstall_T; // @[DCache.scala 181:74]
  wire [3:0] data_wstrb_1 = _data_wstrb_1_T_5 ? io_cpu_M_wmask : bram_replace_wea_1; // @[DCache.scala 180:25]
  wire [7:0] _last_wea_1_T_2 = data_wstrb_1[3] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _last_wea_1_T_5 = data_wstrb_1[2] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _last_wea_1_T_8 = data_wstrb_1[1] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _last_wea_1_T_11 = data_wstrb_1[0] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _last_wea_1_T_12 = {_last_wea_1_T_2,_last_wea_1_T_5,_last_wea_1_T_8,_last_wea_1_T_11}; // @[Cat.scala 33:92]
  reg  write_buffer_axi_busy; // @[DCache.scala 197:38]
  reg [31:0] ar_addr; // @[DCache.scala 199:24]
  reg [7:0] ar_len; // @[DCache.scala 199:24]
  reg [2:0] ar_size; // @[DCache.scala 199:24]
  reg  arvalid; // @[DCache.scala 200:24]
  reg  rready; // @[DCache.scala 203:23]
  reg [31:0] aw_addr; // @[DCache.scala 205:24]
  reg [7:0] aw_len; // @[DCache.scala 205:24]
  reg [2:0] aw_size; // @[DCache.scala 205:24]
  reg  awvalid; // @[DCache.scala 206:24]
  reg [31:0] w_data; // @[DCache.scala 209:23]
  reg [3:0] w_strb; // @[DCache.scala 209:23]
  reg  w_last; // @[DCache.scala 209:23]
  reg  wvalid; // @[DCache.scala 210:23]
  reg  current_mmio_write_saved; // @[DCache.scala 216:41]
  wire  _T = io_axi_aw_ready & io_axi_aw_valid; // @[Decoupled.scala 52:35]
  wire  _GEN_258 = _T ? 1'h0 : awvalid; // @[DCache.scala 220:26 221:15 206:24]
  wire  _T_1 = io_axi_w_ready & io_axi_w_valid; // @[Decoupled.scala 52:35]
  wire  _GEN_259 = _T_1 ? 1'h0 : wvalid; // @[DCache.scala 223:25 224:14 210:23]
  wire  _GEN_260 = _T_1 ? 1'h0 : w_last; // @[DCache.scala 223:25 225:14 209:23]
  wire  _T_2 = io_axi_b_ready & io_axi_b_valid; // @[Decoupled.scala 52:35]
  wire  _T_3 = write_buffer_io_deq_ready & write_buffer_io_deq_valid; // @[Decoupled.scala 52:35]
  wire [2:0] _aw_size_T = {1'h0,write_buffer_io_deq_bits_size}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_262 = _T_3 ? write_buffer_io_deq_bits_addr : aw_addr; // @[DCache.scala 232:36 233:15 205:24]
  wire [2:0] _GEN_263 = _T_3 ? _aw_size_T : aw_size; // @[DCache.scala 232:36 234:15 205:24]
  wire [31:0] _GEN_264 = _T_3 ? write_buffer_io_deq_bits_data : w_data; // @[DCache.scala 232:36 235:15 209:23]
  wire [3:0] _GEN_265 = _T_3 ? write_buffer_io_deq_bits_strb : w_strb; // @[DCache.scala 232:36 236:15 209:23]
  wire  _GEN_266 = write_buffer_io_deq_valid; // @[DCache.scala 230:41 231:31 85:29]
  wire [31:0] _GEN_267 = write_buffer_io_deq_valid ? _GEN_262 : aw_addr; // @[DCache.scala 205:24 230:41]
  wire [2:0] _GEN_268 = write_buffer_io_deq_valid ? _GEN_263 : aw_size; // @[DCache.scala 205:24 230:41]
  wire [31:0] _GEN_269 = write_buffer_io_deq_valid ? _GEN_264 : w_data; // @[DCache.scala 209:23 230:41]
  wire [3:0] _GEN_270 = write_buffer_io_deq_valid ? _GEN_265 : w_strb; // @[DCache.scala 209:23 230:41]
  wire [7:0] _GEN_271 = write_buffer_io_deq_valid ? 8'h0 : aw_len; // @[DCache.scala 205:24 230:41 238:27]
  wire  _GEN_272 = write_buffer_io_deq_valid | awvalid; // @[DCache.scala 206:24 230:41 239:27]
  wire  _GEN_273 = write_buffer_io_deq_valid | w_last; // @[DCache.scala 209:23 230:41 240:27]
  wire  _GEN_274 = write_buffer_io_deq_valid | wvalid; // @[DCache.scala 210:23 230:41 241:27]
  wire  _GEN_275 = write_buffer_io_deq_valid | write_buffer_axi_busy; // @[DCache.scala 230:41 242:27 197:38]
  wire  _GEN_276 = write_buffer_axi_busy ? _GEN_258 : _GEN_272; // @[DCache.scala 219:31]
  wire  _GEN_277 = write_buffer_axi_busy ? _GEN_259 : _GEN_274; // @[DCache.scala 219:31]
  wire  _GEN_278 = write_buffer_axi_busy ? _GEN_260 : _GEN_273; // @[DCache.scala 219:31]
  wire [31:0] _GEN_281 = write_buffer_axi_busy ? aw_addr : _GEN_267; // @[DCache.scala 205:24 219:31]
  wire [2:0] _GEN_282 = write_buffer_axi_busy ? aw_size : _GEN_268; // @[DCache.scala 205:24 219:31]
  wire [31:0] _GEN_283 = write_buffer_axi_busy ? w_data : _GEN_269; // @[DCache.scala 209:23 219:31]
  wire [3:0] _GEN_284 = write_buffer_axi_busy ? w_strb : _GEN_270; // @[DCache.scala 209:23 219:31]
  wire [7:0] _GEN_285 = write_buffer_axi_busy ? aw_len : _GEN_271; // @[DCache.scala 205:24 219:31]
  reg [18:0] tlb2_vpn; // @[DCache.scala 245:21]
  reg  data_tlb_refill; // @[DCache.scala 250:25]
  reg  data_tlb_invalid; // @[DCache.scala 250:25]
  reg  data_tlb_mod; // @[DCache.scala 250:25]
  wire [2:0] _GEN_286 = l1tlb_ok ? 3'h5 : 3'h1; // @[DCache.scala 264:26 265:26 268:22]
  wire  _GEN_287 = l1tlb_ok | data_tlb_mod; // @[DCache.scala 250:25 264:26 266:26]
  wire [19:0] _GEN_288 = l1tlb_ok ? {{1'd0}, tlb2_vpn} : data_vpn; // @[DCache.scala 245:21 264:26 269:22]
  wire  _T_7 = write_buffer_io_enq_ready & ~current_mmio_write_saved; // @[DCache.scala 273:44]
  wire  _write_buffer_io_enq_bits_addr_T = io_cpu_M_mem_size == 2'h2; // @[DCache.scala 276:28]
  wire [31:0] _write_buffer_io_enq_bits_addr_T_2 = {M_mem_pa[31:2],2'h0}; // @[Cat.scala 33:92]
  wire [31:0] _write_buffer_io_enq_bits_addr_T_3 = _write_buffer_io_enq_bits_addr_T ? _write_buffer_io_enq_bits_addr_T_2
     : M_mem_pa; // @[DCache.scala 275:51]
  wire [31:0] _GEN_290 = write_buffer_io_enq_ready & ~current_mmio_write_saved ? _write_buffer_io_enq_bits_addr_T_3 : 32'h0
    ; // @[DCache.scala 273:74 275:45 84:29]
  wire [1:0] _GEN_291 = write_buffer_io_enq_ready & ~current_mmio_write_saved ? io_cpu_M_mem_size : 2'h0; // @[DCache.scala 273:74 280:45 84:29]
  wire [3:0] _GEN_292 = write_buffer_io_enq_ready & ~current_mmio_write_saved ? io_cpu_M_wmask : 4'h0; // @[DCache.scala 273:74 281:45 84:29]
  wire [31:0] _GEN_293 = write_buffer_io_enq_ready & ~current_mmio_write_saved ? io_cpu_M_wdata : 32'h0; // @[DCache.scala 273:74 282:45 84:29]
  wire  _GEN_294 = write_buffer_io_enq_ready & ~current_mmio_write_saved | current_mmio_write_saved; // @[DCache.scala 273:74 284:40 216:41]
  wire  _T_8 = ~io_cpu_dstall; // @[DCache.scala 286:18]
  wire  _T_10 = ~io_cpu_dstall & ~io_cpu_stallM; // @[DCache.scala 286:33]
  wire  _GEN_295 = ~io_cpu_dstall & ~io_cpu_stallM ? 1'h0 : _GEN_294; // @[DCache.scala 286:45 287:40]
  wire  _T_12 = ~_GEN_275; // @[DCache.scala 289:22]
  wire [2:0] _ar_size_T = {1'h0,io_cpu_M_mem_size}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_296 = ~_GEN_275 ? _write_buffer_io_enq_bits_addr_T_3 : ar_addr; // @[DCache.scala 289:77 290:21 199:24]
  wire [7:0] _GEN_297 = ~_GEN_275 ? 8'h0 : ar_len; // @[DCache.scala 289:77 291:21 199:24]
  wire [2:0] _GEN_298 = ~_GEN_275 ? _ar_size_T : ar_size; // @[DCache.scala 289:77 292:21 199:24]
  wire  _GEN_299 = ~_GEN_275 | arvalid; // @[DCache.scala 289:77 293:21 200:24]
  wire [2:0] _GEN_300 = ~_GEN_275 ? 3'h2 : state; // @[DCache.scala 289:77 294:21 65:96]
  wire  _GEN_301 = ~_GEN_275 | rready; // @[DCache.scala 289:77 295:21 203:23]
  wire  _GEN_302 = io_cpu_M_mem_write & _T_7; // @[DCache.scala 272:29 83:29]
  wire [31:0] _GEN_303 = io_cpu_M_mem_write ? _GEN_290 : 32'h0; // @[DCache.scala 272:29 84:29]
  wire [1:0] _GEN_304 = io_cpu_M_mem_write ? _GEN_291 : 2'h0; // @[DCache.scala 272:29 84:29]
  wire [3:0] _GEN_305 = io_cpu_M_mem_write ? _GEN_292 : 4'h0; // @[DCache.scala 272:29 84:29]
  wire [31:0] _GEN_306 = io_cpu_M_mem_write ? _GEN_293 : 32'h0; // @[DCache.scala 272:29 84:29]
  wire  _GEN_307 = io_cpu_M_mem_write ? _GEN_295 : current_mmio_write_saved; // @[DCache.scala 272:29 216:41]
  wire [31:0] _GEN_308 = io_cpu_M_mem_write ? ar_addr : _GEN_296; // @[DCache.scala 199:24 272:29]
  wire [7:0] _GEN_309 = io_cpu_M_mem_write ? ar_len : _GEN_297; // @[DCache.scala 199:24 272:29]
  wire [2:0] _GEN_310 = io_cpu_M_mem_write ? ar_size : _GEN_298; // @[DCache.scala 199:24 272:29]
  wire  _GEN_311 = io_cpu_M_mem_write ? arvalid : _GEN_299; // @[DCache.scala 200:24 272:29]
  wire [2:0] _GEN_312 = io_cpu_M_mem_write ? state : _GEN_300; // @[DCache.scala 272:29 65:96]
  wire  _GEN_313 = io_cpu_M_mem_write ? rready : _GEN_301; // @[DCache.scala 203:23 272:29]
  wire [9:0] _bram_replace_addr_T = {io_cpu_M_mem_va[11:6],4'h0}; // @[Cat.scala 33:92]
  wire  _GEN_315 = 6'h1 == io_cpu_M_mem_va[11:6] ? lru_1 : lru_0; // @[DCache.scala 307:{37,37}]
  wire  _GEN_316 = 6'h2 == io_cpu_M_mem_va[11:6] ? lru_2 : _GEN_315; // @[DCache.scala 307:{37,37}]
  wire  _GEN_317 = 6'h3 == io_cpu_M_mem_va[11:6] ? lru_3 : _GEN_316; // @[DCache.scala 307:{37,37}]
  wire  _GEN_318 = 6'h4 == io_cpu_M_mem_va[11:6] ? lru_4 : _GEN_317; // @[DCache.scala 307:{37,37}]
  wire  _GEN_319 = 6'h5 == io_cpu_M_mem_va[11:6] ? lru_5 : _GEN_318; // @[DCache.scala 307:{37,37}]
  wire  _GEN_320 = 6'h6 == io_cpu_M_mem_va[11:6] ? lru_6 : _GEN_319; // @[DCache.scala 307:{37,37}]
  wire  _GEN_321 = 6'h7 == io_cpu_M_mem_va[11:6] ? lru_7 : _GEN_320; // @[DCache.scala 307:{37,37}]
  wire  _GEN_322 = 6'h8 == io_cpu_M_mem_va[11:6] ? lru_8 : _GEN_321; // @[DCache.scala 307:{37,37}]
  wire  _GEN_323 = 6'h9 == io_cpu_M_mem_va[11:6] ? lru_9 : _GEN_322; // @[DCache.scala 307:{37,37}]
  wire  _GEN_324 = 6'ha == io_cpu_M_mem_va[11:6] ? lru_10 : _GEN_323; // @[DCache.scala 307:{37,37}]
  wire  _GEN_325 = 6'hb == io_cpu_M_mem_va[11:6] ? lru_11 : _GEN_324; // @[DCache.scala 307:{37,37}]
  wire  _GEN_326 = 6'hc == io_cpu_M_mem_va[11:6] ? lru_12 : _GEN_325; // @[DCache.scala 307:{37,37}]
  wire  _GEN_327 = 6'hd == io_cpu_M_mem_va[11:6] ? lru_13 : _GEN_326; // @[DCache.scala 307:{37,37}]
  wire  _GEN_328 = 6'he == io_cpu_M_mem_va[11:6] ? lru_14 : _GEN_327; // @[DCache.scala 307:{37,37}]
  wire  _GEN_329 = 6'hf == io_cpu_M_mem_va[11:6] ? lru_15 : _GEN_328; // @[DCache.scala 307:{37,37}]
  wire  _GEN_330 = 6'h10 == io_cpu_M_mem_va[11:6] ? lru_16 : _GEN_329; // @[DCache.scala 307:{37,37}]
  wire  _GEN_331 = 6'h11 == io_cpu_M_mem_va[11:6] ? lru_17 : _GEN_330; // @[DCache.scala 307:{37,37}]
  wire  _GEN_332 = 6'h12 == io_cpu_M_mem_va[11:6] ? lru_18 : _GEN_331; // @[DCache.scala 307:{37,37}]
  wire  _GEN_333 = 6'h13 == io_cpu_M_mem_va[11:6] ? lru_19 : _GEN_332; // @[DCache.scala 307:{37,37}]
  wire  _GEN_334 = 6'h14 == io_cpu_M_mem_va[11:6] ? lru_20 : _GEN_333; // @[DCache.scala 307:{37,37}]
  wire  _GEN_335 = 6'h15 == io_cpu_M_mem_va[11:6] ? lru_21 : _GEN_334; // @[DCache.scala 307:{37,37}]
  wire  _GEN_336 = 6'h16 == io_cpu_M_mem_va[11:6] ? lru_22 : _GEN_335; // @[DCache.scala 307:{37,37}]
  wire  _GEN_337 = 6'h17 == io_cpu_M_mem_va[11:6] ? lru_23 : _GEN_336; // @[DCache.scala 307:{37,37}]
  wire  _GEN_338 = 6'h18 == io_cpu_M_mem_va[11:6] ? lru_24 : _GEN_337; // @[DCache.scala 307:{37,37}]
  wire  _GEN_339 = 6'h19 == io_cpu_M_mem_va[11:6] ? lru_25 : _GEN_338; // @[DCache.scala 307:{37,37}]
  wire  _GEN_340 = 6'h1a == io_cpu_M_mem_va[11:6] ? lru_26 : _GEN_339; // @[DCache.scala 307:{37,37}]
  wire  _GEN_341 = 6'h1b == io_cpu_M_mem_va[11:6] ? lru_27 : _GEN_340; // @[DCache.scala 307:{37,37}]
  wire  _GEN_342 = 6'h1c == io_cpu_M_mem_va[11:6] ? lru_28 : _GEN_341; // @[DCache.scala 307:{37,37}]
  wire  _GEN_343 = 6'h1d == io_cpu_M_mem_va[11:6] ? lru_29 : _GEN_342; // @[DCache.scala 307:{37,37}]
  wire  _GEN_344 = 6'h1e == io_cpu_M_mem_va[11:6] ? lru_30 : _GEN_343; // @[DCache.scala 307:{37,37}]
  wire  _GEN_345 = 6'h1f == io_cpu_M_mem_va[11:6] ? lru_31 : _GEN_344; // @[DCache.scala 307:{37,37}]
  wire  _GEN_346 = 6'h20 == io_cpu_M_mem_va[11:6] ? lru_32 : _GEN_345; // @[DCache.scala 307:{37,37}]
  wire  _GEN_347 = 6'h21 == io_cpu_M_mem_va[11:6] ? lru_33 : _GEN_346; // @[DCache.scala 307:{37,37}]
  wire  _GEN_348 = 6'h22 == io_cpu_M_mem_va[11:6] ? lru_34 : _GEN_347; // @[DCache.scala 307:{37,37}]
  wire  _GEN_349 = 6'h23 == io_cpu_M_mem_va[11:6] ? lru_35 : _GEN_348; // @[DCache.scala 307:{37,37}]
  wire  _GEN_350 = 6'h24 == io_cpu_M_mem_va[11:6] ? lru_36 : _GEN_349; // @[DCache.scala 307:{37,37}]
  wire  _GEN_351 = 6'h25 == io_cpu_M_mem_va[11:6] ? lru_37 : _GEN_350; // @[DCache.scala 307:{37,37}]
  wire  _GEN_352 = 6'h26 == io_cpu_M_mem_va[11:6] ? lru_38 : _GEN_351; // @[DCache.scala 307:{37,37}]
  wire  _GEN_353 = 6'h27 == io_cpu_M_mem_va[11:6] ? lru_39 : _GEN_352; // @[DCache.scala 307:{37,37}]
  wire  _GEN_354 = 6'h28 == io_cpu_M_mem_va[11:6] ? lru_40 : _GEN_353; // @[DCache.scala 307:{37,37}]
  wire  _GEN_355 = 6'h29 == io_cpu_M_mem_va[11:6] ? lru_41 : _GEN_354; // @[DCache.scala 307:{37,37}]
  wire  _GEN_356 = 6'h2a == io_cpu_M_mem_va[11:6] ? lru_42 : _GEN_355; // @[DCache.scala 307:{37,37}]
  wire  _GEN_357 = 6'h2b == io_cpu_M_mem_va[11:6] ? lru_43 : _GEN_356; // @[DCache.scala 307:{37,37}]
  wire  _GEN_358 = 6'h2c == io_cpu_M_mem_va[11:6] ? lru_44 : _GEN_357; // @[DCache.scala 307:{37,37}]
  wire  _GEN_359 = 6'h2d == io_cpu_M_mem_va[11:6] ? lru_45 : _GEN_358; // @[DCache.scala 307:{37,37}]
  wire  _GEN_360 = 6'h2e == io_cpu_M_mem_va[11:6] ? lru_46 : _GEN_359; // @[DCache.scala 307:{37,37}]
  wire  _GEN_361 = 6'h2f == io_cpu_M_mem_va[11:6] ? lru_47 : _GEN_360; // @[DCache.scala 307:{37,37}]
  wire  _GEN_362 = 6'h30 == io_cpu_M_mem_va[11:6] ? lru_48 : _GEN_361; // @[DCache.scala 307:{37,37}]
  wire  _GEN_363 = 6'h31 == io_cpu_M_mem_va[11:6] ? lru_49 : _GEN_362; // @[DCache.scala 307:{37,37}]
  wire  _GEN_364 = 6'h32 == io_cpu_M_mem_va[11:6] ? lru_50 : _GEN_363; // @[DCache.scala 307:{37,37}]
  wire  _GEN_365 = 6'h33 == io_cpu_M_mem_va[11:6] ? lru_51 : _GEN_364; // @[DCache.scala 307:{37,37}]
  wire  _GEN_366 = 6'h34 == io_cpu_M_mem_va[11:6] ? lru_52 : _GEN_365; // @[DCache.scala 307:{37,37}]
  wire  _GEN_367 = 6'h35 == io_cpu_M_mem_va[11:6] ? lru_53 : _GEN_366; // @[DCache.scala 307:{37,37}]
  wire  _GEN_368 = 6'h36 == io_cpu_M_mem_va[11:6] ? lru_54 : _GEN_367; // @[DCache.scala 307:{37,37}]
  wire  _GEN_369 = 6'h37 == io_cpu_M_mem_va[11:6] ? lru_55 : _GEN_368; // @[DCache.scala 307:{37,37}]
  wire  _GEN_370 = 6'h38 == io_cpu_M_mem_va[11:6] ? lru_56 : _GEN_369; // @[DCache.scala 307:{37,37}]
  wire  _GEN_371 = 6'h39 == io_cpu_M_mem_va[11:6] ? lru_57 : _GEN_370; // @[DCache.scala 307:{37,37}]
  wire  _GEN_372 = 6'h3a == io_cpu_M_mem_va[11:6] ? lru_58 : _GEN_371; // @[DCache.scala 307:{37,37}]
  wire  _GEN_373 = 6'h3b == io_cpu_M_mem_va[11:6] ? lru_59 : _GEN_372; // @[DCache.scala 307:{37,37}]
  wire  _GEN_374 = 6'h3c == io_cpu_M_mem_va[11:6] ? lru_60 : _GEN_373; // @[DCache.scala 307:{37,37}]
  wire  _GEN_375 = 6'h3d == io_cpu_M_mem_va[11:6] ? lru_61 : _GEN_374; // @[DCache.scala 307:{37,37}]
  wire  _GEN_376 = 6'h3e == io_cpu_M_mem_va[11:6] ? lru_62 : _GEN_375; // @[DCache.scala 307:{37,37}]
  wire  _GEN_377 = 6'h3f == io_cpu_M_mem_va[11:6] ? lru_63 : _GEN_376; // @[DCache.scala 307:{37,37}]
  wire  _GEN_378 = 7'h40 == _GEN_1731 ? lru_64 : _GEN_377; // @[DCache.scala 307:{37,37}]
  wire  _GEN_379 = 7'h41 == _GEN_1731 ? lru_65 : _GEN_378; // @[DCache.scala 307:{37,37}]
  wire  _GEN_380 = 7'h42 == _GEN_1731 ? lru_66 : _GEN_379; // @[DCache.scala 307:{37,37}]
  wire  _GEN_381 = 7'h43 == _GEN_1731 ? lru_67 : _GEN_380; // @[DCache.scala 307:{37,37}]
  wire  _GEN_382 = 7'h44 == _GEN_1731 ? lru_68 : _GEN_381; // @[DCache.scala 307:{37,37}]
  wire  _GEN_383 = 7'h45 == _GEN_1731 ? lru_69 : _GEN_382; // @[DCache.scala 307:{37,37}]
  wire  _GEN_384 = 7'h46 == _GEN_1731 ? lru_70 : _GEN_383; // @[DCache.scala 307:{37,37}]
  wire  _GEN_385 = 7'h47 == _GEN_1731 ? lru_71 : _GEN_384; // @[DCache.scala 307:{37,37}]
  wire  _GEN_386 = 7'h48 == _GEN_1731 ? lru_72 : _GEN_385; // @[DCache.scala 307:{37,37}]
  wire  _GEN_387 = 7'h49 == _GEN_1731 ? lru_73 : _GEN_386; // @[DCache.scala 307:{37,37}]
  wire  _GEN_388 = 7'h4a == _GEN_1731 ? lru_74 : _GEN_387; // @[DCache.scala 307:{37,37}]
  wire  _GEN_389 = 7'h4b == _GEN_1731 ? lru_75 : _GEN_388; // @[DCache.scala 307:{37,37}]
  wire  _GEN_390 = 7'h4c == _GEN_1731 ? lru_76 : _GEN_389; // @[DCache.scala 307:{37,37}]
  wire  _GEN_391 = 7'h4d == _GEN_1731 ? lru_77 : _GEN_390; // @[DCache.scala 307:{37,37}]
  wire  _GEN_392 = 7'h4e == _GEN_1731 ? lru_78 : _GEN_391; // @[DCache.scala 307:{37,37}]
  wire  _GEN_393 = 7'h4f == _GEN_1731 ? lru_79 : _GEN_392; // @[DCache.scala 307:{37,37}]
  wire  _GEN_394 = 7'h50 == _GEN_1731 ? lru_80 : _GEN_393; // @[DCache.scala 307:{37,37}]
  wire  _GEN_395 = 7'h51 == _GEN_1731 ? lru_81 : _GEN_394; // @[DCache.scala 307:{37,37}]
  wire  _GEN_396 = 7'h52 == _GEN_1731 ? lru_82 : _GEN_395; // @[DCache.scala 307:{37,37}]
  wire  _GEN_397 = 7'h53 == _GEN_1731 ? lru_83 : _GEN_396; // @[DCache.scala 307:{37,37}]
  wire  _GEN_398 = 7'h54 == _GEN_1731 ? lru_84 : _GEN_397; // @[DCache.scala 307:{37,37}]
  wire  _GEN_399 = 7'h55 == _GEN_1731 ? lru_85 : _GEN_398; // @[DCache.scala 307:{37,37}]
  wire  _GEN_400 = 7'h56 == _GEN_1731 ? lru_86 : _GEN_399; // @[DCache.scala 307:{37,37}]
  wire  _GEN_401 = 7'h57 == _GEN_1731 ? lru_87 : _GEN_400; // @[DCache.scala 307:{37,37}]
  wire  _GEN_402 = 7'h58 == _GEN_1731 ? lru_88 : _GEN_401; // @[DCache.scala 307:{37,37}]
  wire  _GEN_403 = 7'h59 == _GEN_1731 ? lru_89 : _GEN_402; // @[DCache.scala 307:{37,37}]
  wire  _GEN_404 = 7'h5a == _GEN_1731 ? lru_90 : _GEN_403; // @[DCache.scala 307:{37,37}]
  wire  _GEN_405 = 7'h5b == _GEN_1731 ? lru_91 : _GEN_404; // @[DCache.scala 307:{37,37}]
  wire  _GEN_406 = 7'h5c == _GEN_1731 ? lru_92 : _GEN_405; // @[DCache.scala 307:{37,37}]
  wire  _GEN_407 = 7'h5d == _GEN_1731 ? lru_93 : _GEN_406; // @[DCache.scala 307:{37,37}]
  wire  _GEN_408 = 7'h5e == _GEN_1731 ? lru_94 : _GEN_407; // @[DCache.scala 307:{37,37}]
  wire  _GEN_409 = 7'h5f == _GEN_1731 ? lru_95 : _GEN_408; // @[DCache.scala 307:{37,37}]
  wire  _GEN_410 = 7'h60 == _GEN_1731 ? lru_96 : _GEN_409; // @[DCache.scala 307:{37,37}]
  wire  _GEN_411 = 7'h61 == _GEN_1731 ? lru_97 : _GEN_410; // @[DCache.scala 307:{37,37}]
  wire  _GEN_412 = 7'h62 == _GEN_1731 ? lru_98 : _GEN_411; // @[DCache.scala 307:{37,37}]
  wire  _GEN_413 = 7'h63 == _GEN_1731 ? lru_99 : _GEN_412; // @[DCache.scala 307:{37,37}]
  wire  _GEN_414 = 7'h64 == _GEN_1731 ? lru_100 : _GEN_413; // @[DCache.scala 307:{37,37}]
  wire  _GEN_415 = 7'h65 == _GEN_1731 ? lru_101 : _GEN_414; // @[DCache.scala 307:{37,37}]
  wire  _GEN_416 = 7'h66 == _GEN_1731 ? lru_102 : _GEN_415; // @[DCache.scala 307:{37,37}]
  wire  _GEN_417 = 7'h67 == _GEN_1731 ? lru_103 : _GEN_416; // @[DCache.scala 307:{37,37}]
  wire  _GEN_418 = 7'h68 == _GEN_1731 ? lru_104 : _GEN_417; // @[DCache.scala 307:{37,37}]
  wire  _GEN_419 = 7'h69 == _GEN_1731 ? lru_105 : _GEN_418; // @[DCache.scala 307:{37,37}]
  wire  _GEN_420 = 7'h6a == _GEN_1731 ? lru_106 : _GEN_419; // @[DCache.scala 307:{37,37}]
  wire  _GEN_421 = 7'h6b == _GEN_1731 ? lru_107 : _GEN_420; // @[DCache.scala 307:{37,37}]
  wire  _GEN_422 = 7'h6c == _GEN_1731 ? lru_108 : _GEN_421; // @[DCache.scala 307:{37,37}]
  wire  _GEN_423 = 7'h6d == _GEN_1731 ? lru_109 : _GEN_422; // @[DCache.scala 307:{37,37}]
  wire  _GEN_424 = 7'h6e == _GEN_1731 ? lru_110 : _GEN_423; // @[DCache.scala 307:{37,37}]
  wire  _GEN_425 = 7'h6f == _GEN_1731 ? lru_111 : _GEN_424; // @[DCache.scala 307:{37,37}]
  wire  _GEN_426 = 7'h70 == _GEN_1731 ? lru_112 : _GEN_425; // @[DCache.scala 307:{37,37}]
  wire  _GEN_427 = 7'h71 == _GEN_1731 ? lru_113 : _GEN_426; // @[DCache.scala 307:{37,37}]
  wire  _GEN_428 = 7'h72 == _GEN_1731 ? lru_114 : _GEN_427; // @[DCache.scala 307:{37,37}]
  wire  _GEN_429 = 7'h73 == _GEN_1731 ? lru_115 : _GEN_428; // @[DCache.scala 307:{37,37}]
  wire  _GEN_430 = 7'h74 == _GEN_1731 ? lru_116 : _GEN_429; // @[DCache.scala 307:{37,37}]
  wire  _GEN_431 = 7'h75 == _GEN_1731 ? lru_117 : _GEN_430; // @[DCache.scala 307:{37,37}]
  wire  _GEN_432 = 7'h76 == _GEN_1731 ? lru_118 : _GEN_431; // @[DCache.scala 307:{37,37}]
  wire  _GEN_433 = 7'h77 == _GEN_1731 ? lru_119 : _GEN_432; // @[DCache.scala 307:{37,37}]
  wire  _GEN_434 = 7'h78 == _GEN_1731 ? lru_120 : _GEN_433; // @[DCache.scala 307:{37,37}]
  wire  _GEN_435 = 7'h79 == _GEN_1731 ? lru_121 : _GEN_434; // @[DCache.scala 307:{37,37}]
  wire  _GEN_436 = 7'h7a == _GEN_1731 ? lru_122 : _GEN_435; // @[DCache.scala 307:{37,37}]
  wire  _GEN_437 = 7'h7b == _GEN_1731 ? lru_123 : _GEN_436; // @[DCache.scala 307:{37,37}]
  wire  _GEN_438 = 7'h7c == _GEN_1731 ? lru_124 : _GEN_437; // @[DCache.scala 307:{37,37}]
  wire  _GEN_439 = 7'h7d == _GEN_1731 ? lru_125 : _GEN_438; // @[DCache.scala 307:{37,37}]
  wire  _GEN_440 = 7'h7e == _GEN_1731 ? lru_126 : _GEN_439; // @[DCache.scala 307:{37,37}]
  wire  _GEN_441 = 7'h7f == _GEN_1731 ? lru_127 : _GEN_440; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11687 = 6'h0 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_443 = 6'h0 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_0_1 : dirty_0_0; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11688 = 6'h1 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11689 = ~_GEN_441; // @[DCache.scala 307:{37,37}]
  wire  _GEN_444 = 6'h1 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_1_0 : _GEN_443; // @[DCache.scala 307:{37,37}]
  wire  _GEN_445 = 6'h1 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_1_1 : _GEN_444; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11691 = 6'h2 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_446 = 6'h2 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_2_0 : _GEN_445; // @[DCache.scala 307:{37,37}]
  wire  _GEN_447 = 6'h2 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_2_1 : _GEN_446; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11694 = 6'h3 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_448 = 6'h3 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_3_0 : _GEN_447; // @[DCache.scala 307:{37,37}]
  wire  _GEN_449 = 6'h3 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_3_1 : _GEN_448; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11697 = 6'h4 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_450 = 6'h4 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_4_0 : _GEN_449; // @[DCache.scala 307:{37,37}]
  wire  _GEN_451 = 6'h4 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_4_1 : _GEN_450; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11700 = 6'h5 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_452 = 6'h5 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_5_0 : _GEN_451; // @[DCache.scala 307:{37,37}]
  wire  _GEN_453 = 6'h5 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_5_1 : _GEN_452; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11703 = 6'h6 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_454 = 6'h6 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_6_0 : _GEN_453; // @[DCache.scala 307:{37,37}]
  wire  _GEN_455 = 6'h6 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_6_1 : _GEN_454; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11706 = 6'h7 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_456 = 6'h7 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_7_0 : _GEN_455; // @[DCache.scala 307:{37,37}]
  wire  _GEN_457 = 6'h7 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_7_1 : _GEN_456; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11709 = 6'h8 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_458 = 6'h8 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_8_0 : _GEN_457; // @[DCache.scala 307:{37,37}]
  wire  _GEN_459 = 6'h8 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_8_1 : _GEN_458; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11712 = 6'h9 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_460 = 6'h9 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_9_0 : _GEN_459; // @[DCache.scala 307:{37,37}]
  wire  _GEN_461 = 6'h9 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_9_1 : _GEN_460; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11715 = 6'ha == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_462 = 6'ha == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_10_0 : _GEN_461; // @[DCache.scala 307:{37,37}]
  wire  _GEN_463 = 6'ha == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_10_1 : _GEN_462; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11718 = 6'hb == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_464 = 6'hb == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_11_0 : _GEN_463; // @[DCache.scala 307:{37,37}]
  wire  _GEN_465 = 6'hb == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_11_1 : _GEN_464; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11721 = 6'hc == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_466 = 6'hc == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_12_0 : _GEN_465; // @[DCache.scala 307:{37,37}]
  wire  _GEN_467 = 6'hc == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_12_1 : _GEN_466; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11724 = 6'hd == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_468 = 6'hd == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_13_0 : _GEN_467; // @[DCache.scala 307:{37,37}]
  wire  _GEN_469 = 6'hd == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_13_1 : _GEN_468; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11727 = 6'he == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_470 = 6'he == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_14_0 : _GEN_469; // @[DCache.scala 307:{37,37}]
  wire  _GEN_471 = 6'he == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_14_1 : _GEN_470; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11730 = 6'hf == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_472 = 6'hf == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_15_0 : _GEN_471; // @[DCache.scala 307:{37,37}]
  wire  _GEN_473 = 6'hf == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_15_1 : _GEN_472; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11733 = 6'h10 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_474 = 6'h10 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_16_0 : _GEN_473; // @[DCache.scala 307:{37,37}]
  wire  _GEN_475 = 6'h10 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_16_1 : _GEN_474; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11736 = 6'h11 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_476 = 6'h11 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_17_0 : _GEN_475; // @[DCache.scala 307:{37,37}]
  wire  _GEN_477 = 6'h11 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_17_1 : _GEN_476; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11739 = 6'h12 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_478 = 6'h12 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_18_0 : _GEN_477; // @[DCache.scala 307:{37,37}]
  wire  _GEN_479 = 6'h12 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_18_1 : _GEN_478; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11742 = 6'h13 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_480 = 6'h13 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_19_0 : _GEN_479; // @[DCache.scala 307:{37,37}]
  wire  _GEN_481 = 6'h13 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_19_1 : _GEN_480; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11745 = 6'h14 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_482 = 6'h14 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_20_0 : _GEN_481; // @[DCache.scala 307:{37,37}]
  wire  _GEN_483 = 6'h14 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_20_1 : _GEN_482; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11748 = 6'h15 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_484 = 6'h15 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_21_0 : _GEN_483; // @[DCache.scala 307:{37,37}]
  wire  _GEN_485 = 6'h15 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_21_1 : _GEN_484; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11751 = 6'h16 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_486 = 6'h16 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_22_0 : _GEN_485; // @[DCache.scala 307:{37,37}]
  wire  _GEN_487 = 6'h16 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_22_1 : _GEN_486; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11754 = 6'h17 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_488 = 6'h17 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_23_0 : _GEN_487; // @[DCache.scala 307:{37,37}]
  wire  _GEN_489 = 6'h17 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_23_1 : _GEN_488; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11757 = 6'h18 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_490 = 6'h18 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_24_0 : _GEN_489; // @[DCache.scala 307:{37,37}]
  wire  _GEN_491 = 6'h18 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_24_1 : _GEN_490; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11760 = 6'h19 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_492 = 6'h19 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_25_0 : _GEN_491; // @[DCache.scala 307:{37,37}]
  wire  _GEN_493 = 6'h19 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_25_1 : _GEN_492; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11763 = 6'h1a == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_494 = 6'h1a == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_26_0 : _GEN_493; // @[DCache.scala 307:{37,37}]
  wire  _GEN_495 = 6'h1a == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_26_1 : _GEN_494; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11766 = 6'h1b == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_496 = 6'h1b == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_27_0 : _GEN_495; // @[DCache.scala 307:{37,37}]
  wire  _GEN_497 = 6'h1b == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_27_1 : _GEN_496; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11769 = 6'h1c == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_498 = 6'h1c == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_28_0 : _GEN_497; // @[DCache.scala 307:{37,37}]
  wire  _GEN_499 = 6'h1c == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_28_1 : _GEN_498; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11772 = 6'h1d == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_500 = 6'h1d == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_29_0 : _GEN_499; // @[DCache.scala 307:{37,37}]
  wire  _GEN_501 = 6'h1d == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_29_1 : _GEN_500; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11775 = 6'h1e == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_502 = 6'h1e == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_30_0 : _GEN_501; // @[DCache.scala 307:{37,37}]
  wire  _GEN_503 = 6'h1e == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_30_1 : _GEN_502; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11778 = 6'h1f == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_504 = 6'h1f == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_31_0 : _GEN_503; // @[DCache.scala 307:{37,37}]
  wire  _GEN_505 = 6'h1f == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_31_1 : _GEN_504; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11781 = 6'h20 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_506 = 6'h20 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_32_0 : _GEN_505; // @[DCache.scala 307:{37,37}]
  wire  _GEN_507 = 6'h20 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_32_1 : _GEN_506; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11784 = 6'h21 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_508 = 6'h21 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_33_0 : _GEN_507; // @[DCache.scala 307:{37,37}]
  wire  _GEN_509 = 6'h21 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_33_1 : _GEN_508; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11787 = 6'h22 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_510 = 6'h22 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_34_0 : _GEN_509; // @[DCache.scala 307:{37,37}]
  wire  _GEN_511 = 6'h22 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_34_1 : _GEN_510; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11790 = 6'h23 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_512 = 6'h23 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_35_0 : _GEN_511; // @[DCache.scala 307:{37,37}]
  wire  _GEN_513 = 6'h23 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_35_1 : _GEN_512; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11793 = 6'h24 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_514 = 6'h24 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_36_0 : _GEN_513; // @[DCache.scala 307:{37,37}]
  wire  _GEN_515 = 6'h24 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_36_1 : _GEN_514; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11796 = 6'h25 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_516 = 6'h25 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_37_0 : _GEN_515; // @[DCache.scala 307:{37,37}]
  wire  _GEN_517 = 6'h25 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_37_1 : _GEN_516; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11799 = 6'h26 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_518 = 6'h26 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_38_0 : _GEN_517; // @[DCache.scala 307:{37,37}]
  wire  _GEN_519 = 6'h26 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_38_1 : _GEN_518; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11802 = 6'h27 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_520 = 6'h27 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_39_0 : _GEN_519; // @[DCache.scala 307:{37,37}]
  wire  _GEN_521 = 6'h27 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_39_1 : _GEN_520; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11805 = 6'h28 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_522 = 6'h28 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_40_0 : _GEN_521; // @[DCache.scala 307:{37,37}]
  wire  _GEN_523 = 6'h28 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_40_1 : _GEN_522; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11808 = 6'h29 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_524 = 6'h29 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_41_0 : _GEN_523; // @[DCache.scala 307:{37,37}]
  wire  _GEN_525 = 6'h29 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_41_1 : _GEN_524; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11811 = 6'h2a == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_526 = 6'h2a == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_42_0 : _GEN_525; // @[DCache.scala 307:{37,37}]
  wire  _GEN_527 = 6'h2a == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_42_1 : _GEN_526; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11814 = 6'h2b == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_528 = 6'h2b == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_43_0 : _GEN_527; // @[DCache.scala 307:{37,37}]
  wire  _GEN_529 = 6'h2b == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_43_1 : _GEN_528; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11817 = 6'h2c == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_530 = 6'h2c == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_44_0 : _GEN_529; // @[DCache.scala 307:{37,37}]
  wire  _GEN_531 = 6'h2c == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_44_1 : _GEN_530; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11820 = 6'h2d == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_532 = 6'h2d == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_45_0 : _GEN_531; // @[DCache.scala 307:{37,37}]
  wire  _GEN_533 = 6'h2d == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_45_1 : _GEN_532; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11823 = 6'h2e == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_534 = 6'h2e == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_46_0 : _GEN_533; // @[DCache.scala 307:{37,37}]
  wire  _GEN_535 = 6'h2e == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_46_1 : _GEN_534; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11826 = 6'h2f == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_536 = 6'h2f == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_47_0 : _GEN_535; // @[DCache.scala 307:{37,37}]
  wire  _GEN_537 = 6'h2f == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_47_1 : _GEN_536; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11829 = 6'h30 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_538 = 6'h30 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_48_0 : _GEN_537; // @[DCache.scala 307:{37,37}]
  wire  _GEN_539 = 6'h30 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_48_1 : _GEN_538; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11832 = 6'h31 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_540 = 6'h31 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_49_0 : _GEN_539; // @[DCache.scala 307:{37,37}]
  wire  _GEN_541 = 6'h31 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_49_1 : _GEN_540; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11835 = 6'h32 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_542 = 6'h32 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_50_0 : _GEN_541; // @[DCache.scala 307:{37,37}]
  wire  _GEN_543 = 6'h32 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_50_1 : _GEN_542; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11838 = 6'h33 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_544 = 6'h33 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_51_0 : _GEN_543; // @[DCache.scala 307:{37,37}]
  wire  _GEN_545 = 6'h33 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_51_1 : _GEN_544; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11841 = 6'h34 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_546 = 6'h34 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_52_0 : _GEN_545; // @[DCache.scala 307:{37,37}]
  wire  _GEN_547 = 6'h34 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_52_1 : _GEN_546; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11844 = 6'h35 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_548 = 6'h35 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_53_0 : _GEN_547; // @[DCache.scala 307:{37,37}]
  wire  _GEN_549 = 6'h35 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_53_1 : _GEN_548; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11847 = 6'h36 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_550 = 6'h36 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_54_0 : _GEN_549; // @[DCache.scala 307:{37,37}]
  wire  _GEN_551 = 6'h36 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_54_1 : _GEN_550; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11850 = 6'h37 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_552 = 6'h37 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_55_0 : _GEN_551; // @[DCache.scala 307:{37,37}]
  wire  _GEN_553 = 6'h37 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_55_1 : _GEN_552; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11853 = 6'h38 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_554 = 6'h38 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_56_0 : _GEN_553; // @[DCache.scala 307:{37,37}]
  wire  _GEN_555 = 6'h38 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_56_1 : _GEN_554; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11856 = 6'h39 == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_556 = 6'h39 == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_57_0 : _GEN_555; // @[DCache.scala 307:{37,37}]
  wire  _GEN_557 = 6'h39 == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_57_1 : _GEN_556; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11859 = 6'h3a == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_558 = 6'h3a == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_58_0 : _GEN_557; // @[DCache.scala 307:{37,37}]
  wire  _GEN_559 = 6'h3a == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_58_1 : _GEN_558; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11862 = 6'h3b == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_560 = 6'h3b == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_59_0 : _GEN_559; // @[DCache.scala 307:{37,37}]
  wire  _GEN_561 = 6'h3b == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_59_1 : _GEN_560; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11865 = 6'h3c == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_562 = 6'h3c == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_60_0 : _GEN_561; // @[DCache.scala 307:{37,37}]
  wire  _GEN_563 = 6'h3c == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_60_1 : _GEN_562; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11868 = 6'h3d == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_564 = 6'h3d == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_61_0 : _GEN_563; // @[DCache.scala 307:{37,37}]
  wire  _GEN_565 = 6'h3d == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_61_1 : _GEN_564; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11871 = 6'h3e == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_566 = 6'h3e == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_62_0 : _GEN_565; // @[DCache.scala 307:{37,37}]
  wire  _GEN_567 = 6'h3e == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_62_1 : _GEN_566; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11874 = 6'h3f == io_cpu_M_mem_va[11:6]; // @[DCache.scala 307:{37,37}]
  wire  _GEN_568 = 6'h3f == io_cpu_M_mem_va[11:6] & ~_GEN_441 ? dirty_63_0 : _GEN_567; // @[DCache.scala 307:{37,37}]
  wire  _GEN_569 = 6'h3f == io_cpu_M_mem_va[11:6] & _GEN_441 ? dirty_63_1 : _GEN_568; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11878 = 7'h40 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_570 = 7'h40 == _GEN_1731 & ~_GEN_441 ? dirty_64_0 : _GEN_569; // @[DCache.scala 307:{37,37}]
  wire  _GEN_571 = 7'h40 == _GEN_1731 & _GEN_441 ? dirty_64_1 : _GEN_570; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11883 = 7'h41 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_572 = 7'h41 == _GEN_1731 & ~_GEN_441 ? dirty_65_0 : _GEN_571; // @[DCache.scala 307:{37,37}]
  wire  _GEN_573 = 7'h41 == _GEN_1731 & _GEN_441 ? dirty_65_1 : _GEN_572; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11888 = 7'h42 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_574 = 7'h42 == _GEN_1731 & ~_GEN_441 ? dirty_66_0 : _GEN_573; // @[DCache.scala 307:{37,37}]
  wire  _GEN_575 = 7'h42 == _GEN_1731 & _GEN_441 ? dirty_66_1 : _GEN_574; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11893 = 7'h43 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_576 = 7'h43 == _GEN_1731 & ~_GEN_441 ? dirty_67_0 : _GEN_575; // @[DCache.scala 307:{37,37}]
  wire  _GEN_577 = 7'h43 == _GEN_1731 & _GEN_441 ? dirty_67_1 : _GEN_576; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11898 = 7'h44 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_578 = 7'h44 == _GEN_1731 & ~_GEN_441 ? dirty_68_0 : _GEN_577; // @[DCache.scala 307:{37,37}]
  wire  _GEN_579 = 7'h44 == _GEN_1731 & _GEN_441 ? dirty_68_1 : _GEN_578; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11903 = 7'h45 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_580 = 7'h45 == _GEN_1731 & ~_GEN_441 ? dirty_69_0 : _GEN_579; // @[DCache.scala 307:{37,37}]
  wire  _GEN_581 = 7'h45 == _GEN_1731 & _GEN_441 ? dirty_69_1 : _GEN_580; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11908 = 7'h46 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_582 = 7'h46 == _GEN_1731 & ~_GEN_441 ? dirty_70_0 : _GEN_581; // @[DCache.scala 307:{37,37}]
  wire  _GEN_583 = 7'h46 == _GEN_1731 & _GEN_441 ? dirty_70_1 : _GEN_582; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11913 = 7'h47 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_584 = 7'h47 == _GEN_1731 & ~_GEN_441 ? dirty_71_0 : _GEN_583; // @[DCache.scala 307:{37,37}]
  wire  _GEN_585 = 7'h47 == _GEN_1731 & _GEN_441 ? dirty_71_1 : _GEN_584; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11918 = 7'h48 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_586 = 7'h48 == _GEN_1731 & ~_GEN_441 ? dirty_72_0 : _GEN_585; // @[DCache.scala 307:{37,37}]
  wire  _GEN_587 = 7'h48 == _GEN_1731 & _GEN_441 ? dirty_72_1 : _GEN_586; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11923 = 7'h49 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_588 = 7'h49 == _GEN_1731 & ~_GEN_441 ? dirty_73_0 : _GEN_587; // @[DCache.scala 307:{37,37}]
  wire  _GEN_589 = 7'h49 == _GEN_1731 & _GEN_441 ? dirty_73_1 : _GEN_588; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11928 = 7'h4a == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_590 = 7'h4a == _GEN_1731 & ~_GEN_441 ? dirty_74_0 : _GEN_589; // @[DCache.scala 307:{37,37}]
  wire  _GEN_591 = 7'h4a == _GEN_1731 & _GEN_441 ? dirty_74_1 : _GEN_590; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11933 = 7'h4b == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_592 = 7'h4b == _GEN_1731 & ~_GEN_441 ? dirty_75_0 : _GEN_591; // @[DCache.scala 307:{37,37}]
  wire  _GEN_593 = 7'h4b == _GEN_1731 & _GEN_441 ? dirty_75_1 : _GEN_592; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11938 = 7'h4c == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_594 = 7'h4c == _GEN_1731 & ~_GEN_441 ? dirty_76_0 : _GEN_593; // @[DCache.scala 307:{37,37}]
  wire  _GEN_595 = 7'h4c == _GEN_1731 & _GEN_441 ? dirty_76_1 : _GEN_594; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11943 = 7'h4d == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_596 = 7'h4d == _GEN_1731 & ~_GEN_441 ? dirty_77_0 : _GEN_595; // @[DCache.scala 307:{37,37}]
  wire  _GEN_597 = 7'h4d == _GEN_1731 & _GEN_441 ? dirty_77_1 : _GEN_596; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11948 = 7'h4e == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_598 = 7'h4e == _GEN_1731 & ~_GEN_441 ? dirty_78_0 : _GEN_597; // @[DCache.scala 307:{37,37}]
  wire  _GEN_599 = 7'h4e == _GEN_1731 & _GEN_441 ? dirty_78_1 : _GEN_598; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11953 = 7'h4f == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_600 = 7'h4f == _GEN_1731 & ~_GEN_441 ? dirty_79_0 : _GEN_599; // @[DCache.scala 307:{37,37}]
  wire  _GEN_601 = 7'h4f == _GEN_1731 & _GEN_441 ? dirty_79_1 : _GEN_600; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11958 = 7'h50 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_602 = 7'h50 == _GEN_1731 & ~_GEN_441 ? dirty_80_0 : _GEN_601; // @[DCache.scala 307:{37,37}]
  wire  _GEN_603 = 7'h50 == _GEN_1731 & _GEN_441 ? dirty_80_1 : _GEN_602; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11963 = 7'h51 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_604 = 7'h51 == _GEN_1731 & ~_GEN_441 ? dirty_81_0 : _GEN_603; // @[DCache.scala 307:{37,37}]
  wire  _GEN_605 = 7'h51 == _GEN_1731 & _GEN_441 ? dirty_81_1 : _GEN_604; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11968 = 7'h52 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_606 = 7'h52 == _GEN_1731 & ~_GEN_441 ? dirty_82_0 : _GEN_605; // @[DCache.scala 307:{37,37}]
  wire  _GEN_607 = 7'h52 == _GEN_1731 & _GEN_441 ? dirty_82_1 : _GEN_606; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11973 = 7'h53 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_608 = 7'h53 == _GEN_1731 & ~_GEN_441 ? dirty_83_0 : _GEN_607; // @[DCache.scala 307:{37,37}]
  wire  _GEN_609 = 7'h53 == _GEN_1731 & _GEN_441 ? dirty_83_1 : _GEN_608; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11978 = 7'h54 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_610 = 7'h54 == _GEN_1731 & ~_GEN_441 ? dirty_84_0 : _GEN_609; // @[DCache.scala 307:{37,37}]
  wire  _GEN_611 = 7'h54 == _GEN_1731 & _GEN_441 ? dirty_84_1 : _GEN_610; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11983 = 7'h55 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_612 = 7'h55 == _GEN_1731 & ~_GEN_441 ? dirty_85_0 : _GEN_611; // @[DCache.scala 307:{37,37}]
  wire  _GEN_613 = 7'h55 == _GEN_1731 & _GEN_441 ? dirty_85_1 : _GEN_612; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11988 = 7'h56 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_614 = 7'h56 == _GEN_1731 & ~_GEN_441 ? dirty_86_0 : _GEN_613; // @[DCache.scala 307:{37,37}]
  wire  _GEN_615 = 7'h56 == _GEN_1731 & _GEN_441 ? dirty_86_1 : _GEN_614; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11993 = 7'h57 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_616 = 7'h57 == _GEN_1731 & ~_GEN_441 ? dirty_87_0 : _GEN_615; // @[DCache.scala 307:{37,37}]
  wire  _GEN_617 = 7'h57 == _GEN_1731 & _GEN_441 ? dirty_87_1 : _GEN_616; // @[DCache.scala 307:{37,37}]
  wire  _GEN_11998 = 7'h58 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_618 = 7'h58 == _GEN_1731 & ~_GEN_441 ? dirty_88_0 : _GEN_617; // @[DCache.scala 307:{37,37}]
  wire  _GEN_619 = 7'h58 == _GEN_1731 & _GEN_441 ? dirty_88_1 : _GEN_618; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12003 = 7'h59 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_620 = 7'h59 == _GEN_1731 & ~_GEN_441 ? dirty_89_0 : _GEN_619; // @[DCache.scala 307:{37,37}]
  wire  _GEN_621 = 7'h59 == _GEN_1731 & _GEN_441 ? dirty_89_1 : _GEN_620; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12008 = 7'h5a == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_622 = 7'h5a == _GEN_1731 & ~_GEN_441 ? dirty_90_0 : _GEN_621; // @[DCache.scala 307:{37,37}]
  wire  _GEN_623 = 7'h5a == _GEN_1731 & _GEN_441 ? dirty_90_1 : _GEN_622; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12013 = 7'h5b == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_624 = 7'h5b == _GEN_1731 & ~_GEN_441 ? dirty_91_0 : _GEN_623; // @[DCache.scala 307:{37,37}]
  wire  _GEN_625 = 7'h5b == _GEN_1731 & _GEN_441 ? dirty_91_1 : _GEN_624; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12018 = 7'h5c == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_626 = 7'h5c == _GEN_1731 & ~_GEN_441 ? dirty_92_0 : _GEN_625; // @[DCache.scala 307:{37,37}]
  wire  _GEN_627 = 7'h5c == _GEN_1731 & _GEN_441 ? dirty_92_1 : _GEN_626; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12023 = 7'h5d == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_628 = 7'h5d == _GEN_1731 & ~_GEN_441 ? dirty_93_0 : _GEN_627; // @[DCache.scala 307:{37,37}]
  wire  _GEN_629 = 7'h5d == _GEN_1731 & _GEN_441 ? dirty_93_1 : _GEN_628; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12028 = 7'h5e == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_630 = 7'h5e == _GEN_1731 & ~_GEN_441 ? dirty_94_0 : _GEN_629; // @[DCache.scala 307:{37,37}]
  wire  _GEN_631 = 7'h5e == _GEN_1731 & _GEN_441 ? dirty_94_1 : _GEN_630; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12033 = 7'h5f == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_632 = 7'h5f == _GEN_1731 & ~_GEN_441 ? dirty_95_0 : _GEN_631; // @[DCache.scala 307:{37,37}]
  wire  _GEN_633 = 7'h5f == _GEN_1731 & _GEN_441 ? dirty_95_1 : _GEN_632; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12038 = 7'h60 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_634 = 7'h60 == _GEN_1731 & ~_GEN_441 ? dirty_96_0 : _GEN_633; // @[DCache.scala 307:{37,37}]
  wire  _GEN_635 = 7'h60 == _GEN_1731 & _GEN_441 ? dirty_96_1 : _GEN_634; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12043 = 7'h61 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_636 = 7'h61 == _GEN_1731 & ~_GEN_441 ? dirty_97_0 : _GEN_635; // @[DCache.scala 307:{37,37}]
  wire  _GEN_637 = 7'h61 == _GEN_1731 & _GEN_441 ? dirty_97_1 : _GEN_636; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12048 = 7'h62 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_638 = 7'h62 == _GEN_1731 & ~_GEN_441 ? dirty_98_0 : _GEN_637; // @[DCache.scala 307:{37,37}]
  wire  _GEN_639 = 7'h62 == _GEN_1731 & _GEN_441 ? dirty_98_1 : _GEN_638; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12053 = 7'h63 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_640 = 7'h63 == _GEN_1731 & ~_GEN_441 ? dirty_99_0 : _GEN_639; // @[DCache.scala 307:{37,37}]
  wire  _GEN_641 = 7'h63 == _GEN_1731 & _GEN_441 ? dirty_99_1 : _GEN_640; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12058 = 7'h64 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_642 = 7'h64 == _GEN_1731 & ~_GEN_441 ? dirty_100_0 : _GEN_641; // @[DCache.scala 307:{37,37}]
  wire  _GEN_643 = 7'h64 == _GEN_1731 & _GEN_441 ? dirty_100_1 : _GEN_642; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12063 = 7'h65 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_644 = 7'h65 == _GEN_1731 & ~_GEN_441 ? dirty_101_0 : _GEN_643; // @[DCache.scala 307:{37,37}]
  wire  _GEN_645 = 7'h65 == _GEN_1731 & _GEN_441 ? dirty_101_1 : _GEN_644; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12068 = 7'h66 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_646 = 7'h66 == _GEN_1731 & ~_GEN_441 ? dirty_102_0 : _GEN_645; // @[DCache.scala 307:{37,37}]
  wire  _GEN_647 = 7'h66 == _GEN_1731 & _GEN_441 ? dirty_102_1 : _GEN_646; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12073 = 7'h67 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_648 = 7'h67 == _GEN_1731 & ~_GEN_441 ? dirty_103_0 : _GEN_647; // @[DCache.scala 307:{37,37}]
  wire  _GEN_649 = 7'h67 == _GEN_1731 & _GEN_441 ? dirty_103_1 : _GEN_648; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12078 = 7'h68 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_650 = 7'h68 == _GEN_1731 & ~_GEN_441 ? dirty_104_0 : _GEN_649; // @[DCache.scala 307:{37,37}]
  wire  _GEN_651 = 7'h68 == _GEN_1731 & _GEN_441 ? dirty_104_1 : _GEN_650; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12083 = 7'h69 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_652 = 7'h69 == _GEN_1731 & ~_GEN_441 ? dirty_105_0 : _GEN_651; // @[DCache.scala 307:{37,37}]
  wire  _GEN_653 = 7'h69 == _GEN_1731 & _GEN_441 ? dirty_105_1 : _GEN_652; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12088 = 7'h6a == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_654 = 7'h6a == _GEN_1731 & ~_GEN_441 ? dirty_106_0 : _GEN_653; // @[DCache.scala 307:{37,37}]
  wire  _GEN_655 = 7'h6a == _GEN_1731 & _GEN_441 ? dirty_106_1 : _GEN_654; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12093 = 7'h6b == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_656 = 7'h6b == _GEN_1731 & ~_GEN_441 ? dirty_107_0 : _GEN_655; // @[DCache.scala 307:{37,37}]
  wire  _GEN_657 = 7'h6b == _GEN_1731 & _GEN_441 ? dirty_107_1 : _GEN_656; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12098 = 7'h6c == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_658 = 7'h6c == _GEN_1731 & ~_GEN_441 ? dirty_108_0 : _GEN_657; // @[DCache.scala 307:{37,37}]
  wire  _GEN_659 = 7'h6c == _GEN_1731 & _GEN_441 ? dirty_108_1 : _GEN_658; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12103 = 7'h6d == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_660 = 7'h6d == _GEN_1731 & ~_GEN_441 ? dirty_109_0 : _GEN_659; // @[DCache.scala 307:{37,37}]
  wire  _GEN_661 = 7'h6d == _GEN_1731 & _GEN_441 ? dirty_109_1 : _GEN_660; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12108 = 7'h6e == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_662 = 7'h6e == _GEN_1731 & ~_GEN_441 ? dirty_110_0 : _GEN_661; // @[DCache.scala 307:{37,37}]
  wire  _GEN_663 = 7'h6e == _GEN_1731 & _GEN_441 ? dirty_110_1 : _GEN_662; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12113 = 7'h6f == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_664 = 7'h6f == _GEN_1731 & ~_GEN_441 ? dirty_111_0 : _GEN_663; // @[DCache.scala 307:{37,37}]
  wire  _GEN_665 = 7'h6f == _GEN_1731 & _GEN_441 ? dirty_111_1 : _GEN_664; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12118 = 7'h70 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_666 = 7'h70 == _GEN_1731 & ~_GEN_441 ? dirty_112_0 : _GEN_665; // @[DCache.scala 307:{37,37}]
  wire  _GEN_667 = 7'h70 == _GEN_1731 & _GEN_441 ? dirty_112_1 : _GEN_666; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12123 = 7'h71 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_668 = 7'h71 == _GEN_1731 & ~_GEN_441 ? dirty_113_0 : _GEN_667; // @[DCache.scala 307:{37,37}]
  wire  _GEN_669 = 7'h71 == _GEN_1731 & _GEN_441 ? dirty_113_1 : _GEN_668; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12128 = 7'h72 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_670 = 7'h72 == _GEN_1731 & ~_GEN_441 ? dirty_114_0 : _GEN_669; // @[DCache.scala 307:{37,37}]
  wire  _GEN_671 = 7'h72 == _GEN_1731 & _GEN_441 ? dirty_114_1 : _GEN_670; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12133 = 7'h73 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_672 = 7'h73 == _GEN_1731 & ~_GEN_441 ? dirty_115_0 : _GEN_671; // @[DCache.scala 307:{37,37}]
  wire  _GEN_673 = 7'h73 == _GEN_1731 & _GEN_441 ? dirty_115_1 : _GEN_672; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12138 = 7'h74 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_674 = 7'h74 == _GEN_1731 & ~_GEN_441 ? dirty_116_0 : _GEN_673; // @[DCache.scala 307:{37,37}]
  wire  _GEN_675 = 7'h74 == _GEN_1731 & _GEN_441 ? dirty_116_1 : _GEN_674; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12143 = 7'h75 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_676 = 7'h75 == _GEN_1731 & ~_GEN_441 ? dirty_117_0 : _GEN_675; // @[DCache.scala 307:{37,37}]
  wire  _GEN_677 = 7'h75 == _GEN_1731 & _GEN_441 ? dirty_117_1 : _GEN_676; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12148 = 7'h76 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_678 = 7'h76 == _GEN_1731 & ~_GEN_441 ? dirty_118_0 : _GEN_677; // @[DCache.scala 307:{37,37}]
  wire  _GEN_679 = 7'h76 == _GEN_1731 & _GEN_441 ? dirty_118_1 : _GEN_678; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12153 = 7'h77 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_680 = 7'h77 == _GEN_1731 & ~_GEN_441 ? dirty_119_0 : _GEN_679; // @[DCache.scala 307:{37,37}]
  wire  _GEN_681 = 7'h77 == _GEN_1731 & _GEN_441 ? dirty_119_1 : _GEN_680; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12158 = 7'h78 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_682 = 7'h78 == _GEN_1731 & ~_GEN_441 ? dirty_120_0 : _GEN_681; // @[DCache.scala 307:{37,37}]
  wire  _GEN_683 = 7'h78 == _GEN_1731 & _GEN_441 ? dirty_120_1 : _GEN_682; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12163 = 7'h79 == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_684 = 7'h79 == _GEN_1731 & ~_GEN_441 ? dirty_121_0 : _GEN_683; // @[DCache.scala 307:{37,37}]
  wire  _GEN_685 = 7'h79 == _GEN_1731 & _GEN_441 ? dirty_121_1 : _GEN_684; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12168 = 7'h7a == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_686 = 7'h7a == _GEN_1731 & ~_GEN_441 ? dirty_122_0 : _GEN_685; // @[DCache.scala 307:{37,37}]
  wire  _GEN_687 = 7'h7a == _GEN_1731 & _GEN_441 ? dirty_122_1 : _GEN_686; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12173 = 7'h7b == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_688 = 7'h7b == _GEN_1731 & ~_GEN_441 ? dirty_123_0 : _GEN_687; // @[DCache.scala 307:{37,37}]
  wire  _GEN_689 = 7'h7b == _GEN_1731 & _GEN_441 ? dirty_123_1 : _GEN_688; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12178 = 7'h7c == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_690 = 7'h7c == _GEN_1731 & ~_GEN_441 ? dirty_124_0 : _GEN_689; // @[DCache.scala 307:{37,37}]
  wire  _GEN_691 = 7'h7c == _GEN_1731 & _GEN_441 ? dirty_124_1 : _GEN_690; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12183 = 7'h7d == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_692 = 7'h7d == _GEN_1731 & ~_GEN_441 ? dirty_125_0 : _GEN_691; // @[DCache.scala 307:{37,37}]
  wire  _GEN_693 = 7'h7d == _GEN_1731 & _GEN_441 ? dirty_125_1 : _GEN_692; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12188 = 7'h7e == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_694 = 7'h7e == _GEN_1731 & ~_GEN_441 ? dirty_126_0 : _GEN_693; // @[DCache.scala 307:{37,37}]
  wire  _GEN_695 = 7'h7e == _GEN_1731 & _GEN_441 ? dirty_126_1 : _GEN_694; // @[DCache.scala 307:{37,37}]
  wire  _GEN_12193 = 7'h7f == _GEN_1731; // @[DCache.scala 307:{37,37}]
  wire  _GEN_696 = 7'h7f == _GEN_1731 & ~_GEN_441 ? dirty_127_0 : _GEN_695; // @[DCache.scala 307:{37,37}]
  wire  _GEN_697 = 7'h7f == _GEN_1731 & _GEN_441 ? dirty_127_1 : _GEN_696; // @[DCache.scala 307:{37,37}]
  wire  _lru_T = ~tag_compare_valid_1; // @[DCache.scala 311:36]
  wire  _GEN_698 = 6'h0 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_0; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_699 = 6'h1 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_1; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_700 = 6'h2 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_2; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_701 = 6'h3 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_3; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_702 = 6'h4 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_4; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_703 = 6'h5 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_5; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_704 = 6'h6 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_6; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_705 = 6'h7 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_7; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_706 = 6'h8 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_8; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_707 = 6'h9 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_9; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_708 = 6'ha == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_10; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_709 = 6'hb == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_11; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_710 = 6'hc == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_12; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_711 = 6'hd == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_13; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_712 = 6'he == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_14; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_713 = 6'hf == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_15; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_714 = 6'h10 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_16; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_715 = 6'h11 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_17; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_716 = 6'h12 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_18; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_717 = 6'h13 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_19; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_718 = 6'h14 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_20; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_719 = 6'h15 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_21; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_720 = 6'h16 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_22; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_721 = 6'h17 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_23; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_722 = 6'h18 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_24; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_723 = 6'h19 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_25; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_724 = 6'h1a == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_26; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_725 = 6'h1b == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_27; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_726 = 6'h1c == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_28; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_727 = 6'h1d == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_29; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_728 = 6'h1e == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_30; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_729 = 6'h1f == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_31; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_730 = 6'h20 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_32; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_731 = 6'h21 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_33; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_732 = 6'h22 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_34; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_733 = 6'h23 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_35; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_734 = 6'h24 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_36; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_735 = 6'h25 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_37; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_736 = 6'h26 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_38; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_737 = 6'h27 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_39; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_738 = 6'h28 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_40; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_739 = 6'h29 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_41; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_740 = 6'h2a == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_42; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_741 = 6'h2b == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_43; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_742 = 6'h2c == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_44; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_743 = 6'h2d == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_45; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_744 = 6'h2e == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_46; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_745 = 6'h2f == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_47; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_746 = 6'h30 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_48; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_747 = 6'h31 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_49; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_748 = 6'h32 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_50; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_749 = 6'h33 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_51; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_750 = 6'h34 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_52; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_751 = 6'h35 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_53; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_752 = 6'h36 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_54; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_753 = 6'h37 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_55; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_754 = 6'h38 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_56; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_755 = 6'h39 == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_57; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_756 = 6'h3a == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_58; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_757 = 6'h3b == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_59; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_758 = 6'h3c == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_60; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_759 = 6'h3d == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_61; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_760 = 6'h3e == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_62; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_761 = 6'h3f == io_cpu_M_mem_va[11:6] ? ~tag_compare_valid_1 : lru_63; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_762 = 7'h40 == _GEN_1731 ? ~tag_compare_valid_1 : lru_64; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_763 = 7'h41 == _GEN_1731 ? ~tag_compare_valid_1 : lru_65; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_764 = 7'h42 == _GEN_1731 ? ~tag_compare_valid_1 : lru_66; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_765 = 7'h43 == _GEN_1731 ? ~tag_compare_valid_1 : lru_67; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_766 = 7'h44 == _GEN_1731 ? ~tag_compare_valid_1 : lru_68; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_767 = 7'h45 == _GEN_1731 ? ~tag_compare_valid_1 : lru_69; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_768 = 7'h46 == _GEN_1731 ? ~tag_compare_valid_1 : lru_70; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_769 = 7'h47 == _GEN_1731 ? ~tag_compare_valid_1 : lru_71; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_770 = 7'h48 == _GEN_1731 ? ~tag_compare_valid_1 : lru_72; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_771 = 7'h49 == _GEN_1731 ? ~tag_compare_valid_1 : lru_73; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_772 = 7'h4a == _GEN_1731 ? ~tag_compare_valid_1 : lru_74; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_773 = 7'h4b == _GEN_1731 ? ~tag_compare_valid_1 : lru_75; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_774 = 7'h4c == _GEN_1731 ? ~tag_compare_valid_1 : lru_76; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_775 = 7'h4d == _GEN_1731 ? ~tag_compare_valid_1 : lru_77; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_776 = 7'h4e == _GEN_1731 ? ~tag_compare_valid_1 : lru_78; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_777 = 7'h4f == _GEN_1731 ? ~tag_compare_valid_1 : lru_79; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_778 = 7'h50 == _GEN_1731 ? ~tag_compare_valid_1 : lru_80; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_779 = 7'h51 == _GEN_1731 ? ~tag_compare_valid_1 : lru_81; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_780 = 7'h52 == _GEN_1731 ? ~tag_compare_valid_1 : lru_82; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_781 = 7'h53 == _GEN_1731 ? ~tag_compare_valid_1 : lru_83; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_782 = 7'h54 == _GEN_1731 ? ~tag_compare_valid_1 : lru_84; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_783 = 7'h55 == _GEN_1731 ? ~tag_compare_valid_1 : lru_85; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_784 = 7'h56 == _GEN_1731 ? ~tag_compare_valid_1 : lru_86; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_785 = 7'h57 == _GEN_1731 ? ~tag_compare_valid_1 : lru_87; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_786 = 7'h58 == _GEN_1731 ? ~tag_compare_valid_1 : lru_88; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_787 = 7'h59 == _GEN_1731 ? ~tag_compare_valid_1 : lru_89; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_788 = 7'h5a == _GEN_1731 ? ~tag_compare_valid_1 : lru_90; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_789 = 7'h5b == _GEN_1731 ? ~tag_compare_valid_1 : lru_91; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_790 = 7'h5c == _GEN_1731 ? ~tag_compare_valid_1 : lru_92; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_791 = 7'h5d == _GEN_1731 ? ~tag_compare_valid_1 : lru_93; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_792 = 7'h5e == _GEN_1731 ? ~tag_compare_valid_1 : lru_94; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_793 = 7'h5f == _GEN_1731 ? ~tag_compare_valid_1 : lru_95; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_794 = 7'h60 == _GEN_1731 ? ~tag_compare_valid_1 : lru_96; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_795 = 7'h61 == _GEN_1731 ? ~tag_compare_valid_1 : lru_97; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_796 = 7'h62 == _GEN_1731 ? ~tag_compare_valid_1 : lru_98; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_797 = 7'h63 == _GEN_1731 ? ~tag_compare_valid_1 : lru_99; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_798 = 7'h64 == _GEN_1731 ? ~tag_compare_valid_1 : lru_100; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_799 = 7'h65 == _GEN_1731 ? ~tag_compare_valid_1 : lru_101; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_800 = 7'h66 == _GEN_1731 ? ~tag_compare_valid_1 : lru_102; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_801 = 7'h67 == _GEN_1731 ? ~tag_compare_valid_1 : lru_103; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_802 = 7'h68 == _GEN_1731 ? ~tag_compare_valid_1 : lru_104; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_803 = 7'h69 == _GEN_1731 ? ~tag_compare_valid_1 : lru_105; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_804 = 7'h6a == _GEN_1731 ? ~tag_compare_valid_1 : lru_106; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_805 = 7'h6b == _GEN_1731 ? ~tag_compare_valid_1 : lru_107; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_806 = 7'h6c == _GEN_1731 ? ~tag_compare_valid_1 : lru_108; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_807 = 7'h6d == _GEN_1731 ? ~tag_compare_valid_1 : lru_109; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_808 = 7'h6e == _GEN_1731 ? ~tag_compare_valid_1 : lru_110; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_809 = 7'h6f == _GEN_1731 ? ~tag_compare_valid_1 : lru_111; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_810 = 7'h70 == _GEN_1731 ? ~tag_compare_valid_1 : lru_112; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_811 = 7'h71 == _GEN_1731 ? ~tag_compare_valid_1 : lru_113; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_812 = 7'h72 == _GEN_1731 ? ~tag_compare_valid_1 : lru_114; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_813 = 7'h73 == _GEN_1731 ? ~tag_compare_valid_1 : lru_115; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_814 = 7'h74 == _GEN_1731 ? ~tag_compare_valid_1 : lru_116; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_815 = 7'h75 == _GEN_1731 ? ~tag_compare_valid_1 : lru_117; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_816 = 7'h76 == _GEN_1731 ? ~tag_compare_valid_1 : lru_118; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_817 = 7'h77 == _GEN_1731 ? ~tag_compare_valid_1 : lru_119; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_818 = 7'h78 == _GEN_1731 ? ~tag_compare_valid_1 : lru_120; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_819 = 7'h79 == _GEN_1731 ? ~tag_compare_valid_1 : lru_121; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_820 = 7'h7a == _GEN_1731 ? ~tag_compare_valid_1 : lru_122; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_821 = 7'h7b == _GEN_1731 ? ~tag_compare_valid_1 : lru_123; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_822 = 7'h7c == _GEN_1731 ? ~tag_compare_valid_1 : lru_124; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_823 = 7'h7d == _GEN_1731 ? ~tag_compare_valid_1 : lru_125; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_824 = 7'h7e == _GEN_1731 ? ~tag_compare_valid_1 : lru_126; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_825 = 7'h7f == _GEN_1731 ? ~tag_compare_valid_1 : lru_127; // @[DCache.scala 311:{33,33} 70:22]
  wire  _GEN_826 = _GEN_11687 & _lru_T | dirty_0_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_827 = _GEN_11687 & tag_compare_valid_1 | dirty_0_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_828 = _GEN_11688 & _lru_T | dirty_1_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_829 = _GEN_11688 & tag_compare_valid_1 | dirty_1_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_830 = _GEN_11691 & _lru_T | dirty_2_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_831 = _GEN_11691 & tag_compare_valid_1 | dirty_2_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_832 = _GEN_11694 & _lru_T | dirty_3_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_833 = _GEN_11694 & tag_compare_valid_1 | dirty_3_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_834 = _GEN_11697 & _lru_T | dirty_4_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_835 = _GEN_11697 & tag_compare_valid_1 | dirty_4_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_836 = _GEN_11700 & _lru_T | dirty_5_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_837 = _GEN_11700 & tag_compare_valid_1 | dirty_5_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_838 = _GEN_11703 & _lru_T | dirty_6_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_839 = _GEN_11703 & tag_compare_valid_1 | dirty_6_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_840 = _GEN_11706 & _lru_T | dirty_7_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_841 = _GEN_11706 & tag_compare_valid_1 | dirty_7_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_842 = _GEN_11709 & _lru_T | dirty_8_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_843 = _GEN_11709 & tag_compare_valid_1 | dirty_8_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_844 = _GEN_11712 & _lru_T | dirty_9_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_845 = _GEN_11712 & tag_compare_valid_1 | dirty_9_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_846 = _GEN_11715 & _lru_T | dirty_10_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_847 = _GEN_11715 & tag_compare_valid_1 | dirty_10_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_848 = _GEN_11718 & _lru_T | dirty_11_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_849 = _GEN_11718 & tag_compare_valid_1 | dirty_11_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_850 = _GEN_11721 & _lru_T | dirty_12_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_851 = _GEN_11721 & tag_compare_valid_1 | dirty_12_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_852 = _GEN_11724 & _lru_T | dirty_13_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_853 = _GEN_11724 & tag_compare_valid_1 | dirty_13_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_854 = _GEN_11727 & _lru_T | dirty_14_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_855 = _GEN_11727 & tag_compare_valid_1 | dirty_14_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_856 = _GEN_11730 & _lru_T | dirty_15_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_857 = _GEN_11730 & tag_compare_valid_1 | dirty_15_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_858 = _GEN_11733 & _lru_T | dirty_16_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_859 = _GEN_11733 & tag_compare_valid_1 | dirty_16_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_860 = _GEN_11736 & _lru_T | dirty_17_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_861 = _GEN_11736 & tag_compare_valid_1 | dirty_17_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_862 = _GEN_11739 & _lru_T | dirty_18_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_863 = _GEN_11739 & tag_compare_valid_1 | dirty_18_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_864 = _GEN_11742 & _lru_T | dirty_19_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_865 = _GEN_11742 & tag_compare_valid_1 | dirty_19_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_866 = _GEN_11745 & _lru_T | dirty_20_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_867 = _GEN_11745 & tag_compare_valid_1 | dirty_20_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_868 = _GEN_11748 & _lru_T | dirty_21_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_869 = _GEN_11748 & tag_compare_valid_1 | dirty_21_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_870 = _GEN_11751 & _lru_T | dirty_22_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_871 = _GEN_11751 & tag_compare_valid_1 | dirty_22_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_872 = _GEN_11754 & _lru_T | dirty_23_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_873 = _GEN_11754 & tag_compare_valid_1 | dirty_23_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_874 = _GEN_11757 & _lru_T | dirty_24_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_875 = _GEN_11757 & tag_compare_valid_1 | dirty_24_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_876 = _GEN_11760 & _lru_T | dirty_25_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_877 = _GEN_11760 & tag_compare_valid_1 | dirty_25_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_878 = _GEN_11763 & _lru_T | dirty_26_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_879 = _GEN_11763 & tag_compare_valid_1 | dirty_26_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_880 = _GEN_11766 & _lru_T | dirty_27_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_881 = _GEN_11766 & tag_compare_valid_1 | dirty_27_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_882 = _GEN_11769 & _lru_T | dirty_28_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_883 = _GEN_11769 & tag_compare_valid_1 | dirty_28_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_884 = _GEN_11772 & _lru_T | dirty_29_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_885 = _GEN_11772 & tag_compare_valid_1 | dirty_29_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_886 = _GEN_11775 & _lru_T | dirty_30_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_887 = _GEN_11775 & tag_compare_valid_1 | dirty_30_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_888 = _GEN_11778 & _lru_T | dirty_31_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_889 = _GEN_11778 & tag_compare_valid_1 | dirty_31_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_890 = _GEN_11781 & _lru_T | dirty_32_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_891 = _GEN_11781 & tag_compare_valid_1 | dirty_32_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_892 = _GEN_11784 & _lru_T | dirty_33_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_893 = _GEN_11784 & tag_compare_valid_1 | dirty_33_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_894 = _GEN_11787 & _lru_T | dirty_34_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_895 = _GEN_11787 & tag_compare_valid_1 | dirty_34_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_896 = _GEN_11790 & _lru_T | dirty_35_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_897 = _GEN_11790 & tag_compare_valid_1 | dirty_35_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_898 = _GEN_11793 & _lru_T | dirty_36_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_899 = _GEN_11793 & tag_compare_valid_1 | dirty_36_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_900 = _GEN_11796 & _lru_T | dirty_37_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_901 = _GEN_11796 & tag_compare_valid_1 | dirty_37_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_902 = _GEN_11799 & _lru_T | dirty_38_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_903 = _GEN_11799 & tag_compare_valid_1 | dirty_38_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_904 = _GEN_11802 & _lru_T | dirty_39_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_905 = _GEN_11802 & tag_compare_valid_1 | dirty_39_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_906 = _GEN_11805 & _lru_T | dirty_40_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_907 = _GEN_11805 & tag_compare_valid_1 | dirty_40_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_908 = _GEN_11808 & _lru_T | dirty_41_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_909 = _GEN_11808 & tag_compare_valid_1 | dirty_41_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_910 = _GEN_11811 & _lru_T | dirty_42_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_911 = _GEN_11811 & tag_compare_valid_1 | dirty_42_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_912 = _GEN_11814 & _lru_T | dirty_43_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_913 = _GEN_11814 & tag_compare_valid_1 | dirty_43_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_914 = _GEN_11817 & _lru_T | dirty_44_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_915 = _GEN_11817 & tag_compare_valid_1 | dirty_44_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_916 = _GEN_11820 & _lru_T | dirty_45_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_917 = _GEN_11820 & tag_compare_valid_1 | dirty_45_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_918 = _GEN_11823 & _lru_T | dirty_46_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_919 = _GEN_11823 & tag_compare_valid_1 | dirty_46_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_920 = _GEN_11826 & _lru_T | dirty_47_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_921 = _GEN_11826 & tag_compare_valid_1 | dirty_47_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_922 = _GEN_11829 & _lru_T | dirty_48_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_923 = _GEN_11829 & tag_compare_valid_1 | dirty_48_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_924 = _GEN_11832 & _lru_T | dirty_49_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_925 = _GEN_11832 & tag_compare_valid_1 | dirty_49_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_926 = _GEN_11835 & _lru_T | dirty_50_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_927 = _GEN_11835 & tag_compare_valid_1 | dirty_50_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_928 = _GEN_11838 & _lru_T | dirty_51_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_929 = _GEN_11838 & tag_compare_valid_1 | dirty_51_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_930 = _GEN_11841 & _lru_T | dirty_52_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_931 = _GEN_11841 & tag_compare_valid_1 | dirty_52_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_932 = _GEN_11844 & _lru_T | dirty_53_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_933 = _GEN_11844 & tag_compare_valid_1 | dirty_53_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_934 = _GEN_11847 & _lru_T | dirty_54_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_935 = _GEN_11847 & tag_compare_valid_1 | dirty_54_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_936 = _GEN_11850 & _lru_T | dirty_55_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_937 = _GEN_11850 & tag_compare_valid_1 | dirty_55_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_938 = _GEN_11853 & _lru_T | dirty_56_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_939 = _GEN_11853 & tag_compare_valid_1 | dirty_56_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_940 = _GEN_11856 & _lru_T | dirty_57_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_941 = _GEN_11856 & tag_compare_valid_1 | dirty_57_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_942 = _GEN_11859 & _lru_T | dirty_58_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_943 = _GEN_11859 & tag_compare_valid_1 | dirty_58_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_944 = _GEN_11862 & _lru_T | dirty_59_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_945 = _GEN_11862 & tag_compare_valid_1 | dirty_59_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_946 = _GEN_11865 & _lru_T | dirty_60_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_947 = _GEN_11865 & tag_compare_valid_1 | dirty_60_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_948 = _GEN_11868 & _lru_T | dirty_61_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_949 = _GEN_11868 & tag_compare_valid_1 | dirty_61_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_950 = _GEN_11871 & _lru_T | dirty_62_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_951 = _GEN_11871 & tag_compare_valid_1 | dirty_62_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_952 = _GEN_11874 & _lru_T | dirty_63_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_953 = _GEN_11874 & tag_compare_valid_1 | dirty_63_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_954 = _GEN_11878 & _lru_T | dirty_64_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_955 = _GEN_11878 & tag_compare_valid_1 | dirty_64_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_956 = _GEN_11883 & _lru_T | dirty_65_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_957 = _GEN_11883 & tag_compare_valid_1 | dirty_65_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_958 = _GEN_11888 & _lru_T | dirty_66_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_959 = _GEN_11888 & tag_compare_valid_1 | dirty_66_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_960 = _GEN_11893 & _lru_T | dirty_67_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_961 = _GEN_11893 & tag_compare_valid_1 | dirty_67_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_962 = _GEN_11898 & _lru_T | dirty_68_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_963 = _GEN_11898 & tag_compare_valid_1 | dirty_68_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_964 = _GEN_11903 & _lru_T | dirty_69_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_965 = _GEN_11903 & tag_compare_valid_1 | dirty_69_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_966 = _GEN_11908 & _lru_T | dirty_70_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_967 = _GEN_11908 & tag_compare_valid_1 | dirty_70_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_968 = _GEN_11913 & _lru_T | dirty_71_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_969 = _GEN_11913 & tag_compare_valid_1 | dirty_71_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_970 = _GEN_11918 & _lru_T | dirty_72_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_971 = _GEN_11918 & tag_compare_valid_1 | dirty_72_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_972 = _GEN_11923 & _lru_T | dirty_73_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_973 = _GEN_11923 & tag_compare_valid_1 | dirty_73_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_974 = _GEN_11928 & _lru_T | dirty_74_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_975 = _GEN_11928 & tag_compare_valid_1 | dirty_74_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_976 = _GEN_11933 & _lru_T | dirty_75_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_977 = _GEN_11933 & tag_compare_valid_1 | dirty_75_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_978 = _GEN_11938 & _lru_T | dirty_76_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_979 = _GEN_11938 & tag_compare_valid_1 | dirty_76_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_980 = _GEN_11943 & _lru_T | dirty_77_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_981 = _GEN_11943 & tag_compare_valid_1 | dirty_77_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_982 = _GEN_11948 & _lru_T | dirty_78_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_983 = _GEN_11948 & tag_compare_valid_1 | dirty_78_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_984 = _GEN_11953 & _lru_T | dirty_79_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_985 = _GEN_11953 & tag_compare_valid_1 | dirty_79_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_986 = _GEN_11958 & _lru_T | dirty_80_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_987 = _GEN_11958 & tag_compare_valid_1 | dirty_80_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_988 = _GEN_11963 & _lru_T | dirty_81_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_989 = _GEN_11963 & tag_compare_valid_1 | dirty_81_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_990 = _GEN_11968 & _lru_T | dirty_82_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_991 = _GEN_11968 & tag_compare_valid_1 | dirty_82_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_992 = _GEN_11973 & _lru_T | dirty_83_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_993 = _GEN_11973 & tag_compare_valid_1 | dirty_83_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_994 = _GEN_11978 & _lru_T | dirty_84_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_995 = _GEN_11978 & tag_compare_valid_1 | dirty_84_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_996 = _GEN_11983 & _lru_T | dirty_85_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_997 = _GEN_11983 & tag_compare_valid_1 | dirty_85_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_998 = _GEN_11988 & _lru_T | dirty_86_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_999 = _GEN_11988 & tag_compare_valid_1 | dirty_86_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1000 = _GEN_11993 & _lru_T | dirty_87_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1001 = _GEN_11993 & tag_compare_valid_1 | dirty_87_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1002 = _GEN_11998 & _lru_T | dirty_88_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1003 = _GEN_11998 & tag_compare_valid_1 | dirty_88_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1004 = _GEN_12003 & _lru_T | dirty_89_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1005 = _GEN_12003 & tag_compare_valid_1 | dirty_89_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1006 = _GEN_12008 & _lru_T | dirty_90_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1007 = _GEN_12008 & tag_compare_valid_1 | dirty_90_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1008 = _GEN_12013 & _lru_T | dirty_91_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1009 = _GEN_12013 & tag_compare_valid_1 | dirty_91_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1010 = _GEN_12018 & _lru_T | dirty_92_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1011 = _GEN_12018 & tag_compare_valid_1 | dirty_92_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1012 = _GEN_12023 & _lru_T | dirty_93_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1013 = _GEN_12023 & tag_compare_valid_1 | dirty_93_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1014 = _GEN_12028 & _lru_T | dirty_94_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1015 = _GEN_12028 & tag_compare_valid_1 | dirty_94_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1016 = _GEN_12033 & _lru_T | dirty_95_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1017 = _GEN_12033 & tag_compare_valid_1 | dirty_95_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1018 = _GEN_12038 & _lru_T | dirty_96_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1019 = _GEN_12038 & tag_compare_valid_1 | dirty_96_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1020 = _GEN_12043 & _lru_T | dirty_97_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1021 = _GEN_12043 & tag_compare_valid_1 | dirty_97_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1022 = _GEN_12048 & _lru_T | dirty_98_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1023 = _GEN_12048 & tag_compare_valid_1 | dirty_98_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1024 = _GEN_12053 & _lru_T | dirty_99_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1025 = _GEN_12053 & tag_compare_valid_1 | dirty_99_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1026 = _GEN_12058 & _lru_T | dirty_100_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1027 = _GEN_12058 & tag_compare_valid_1 | dirty_100_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1028 = _GEN_12063 & _lru_T | dirty_101_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1029 = _GEN_12063 & tag_compare_valid_1 | dirty_101_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1030 = _GEN_12068 & _lru_T | dirty_102_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1031 = _GEN_12068 & tag_compare_valid_1 | dirty_102_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1032 = _GEN_12073 & _lru_T | dirty_103_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1033 = _GEN_12073 & tag_compare_valid_1 | dirty_103_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1034 = _GEN_12078 & _lru_T | dirty_104_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1035 = _GEN_12078 & tag_compare_valid_1 | dirty_104_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1036 = _GEN_12083 & _lru_T | dirty_105_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1037 = _GEN_12083 & tag_compare_valid_1 | dirty_105_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1038 = _GEN_12088 & _lru_T | dirty_106_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1039 = _GEN_12088 & tag_compare_valid_1 | dirty_106_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1040 = _GEN_12093 & _lru_T | dirty_107_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1041 = _GEN_12093 & tag_compare_valid_1 | dirty_107_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1042 = _GEN_12098 & _lru_T | dirty_108_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1043 = _GEN_12098 & tag_compare_valid_1 | dirty_108_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1044 = _GEN_12103 & _lru_T | dirty_109_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1045 = _GEN_12103 & tag_compare_valid_1 | dirty_109_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1046 = _GEN_12108 & _lru_T | dirty_110_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1047 = _GEN_12108 & tag_compare_valid_1 | dirty_110_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1048 = _GEN_12113 & _lru_T | dirty_111_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1049 = _GEN_12113 & tag_compare_valid_1 | dirty_111_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1050 = _GEN_12118 & _lru_T | dirty_112_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1051 = _GEN_12118 & tag_compare_valid_1 | dirty_112_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1052 = _GEN_12123 & _lru_T | dirty_113_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1053 = _GEN_12123 & tag_compare_valid_1 | dirty_113_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1054 = _GEN_12128 & _lru_T | dirty_114_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1055 = _GEN_12128 & tag_compare_valid_1 | dirty_114_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1056 = _GEN_12133 & _lru_T | dirty_115_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1057 = _GEN_12133 & tag_compare_valid_1 | dirty_115_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1058 = _GEN_12138 & _lru_T | dirty_116_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1059 = _GEN_12138 & tag_compare_valid_1 | dirty_116_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1060 = _GEN_12143 & _lru_T | dirty_117_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1061 = _GEN_12143 & tag_compare_valid_1 | dirty_117_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1062 = _GEN_12148 & _lru_T | dirty_118_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1063 = _GEN_12148 & tag_compare_valid_1 | dirty_118_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1064 = _GEN_12153 & _lru_T | dirty_119_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1065 = _GEN_12153 & tag_compare_valid_1 | dirty_119_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1066 = _GEN_12158 & _lru_T | dirty_120_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1067 = _GEN_12158 & tag_compare_valid_1 | dirty_120_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1068 = _GEN_12163 & _lru_T | dirty_121_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1069 = _GEN_12163 & tag_compare_valid_1 | dirty_121_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1070 = _GEN_12168 & _lru_T | dirty_122_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1071 = _GEN_12168 & tag_compare_valid_1 | dirty_122_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1072 = _GEN_12173 & _lru_T | dirty_123_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1073 = _GEN_12173 & tag_compare_valid_1 | dirty_123_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1074 = _GEN_12178 & _lru_T | dirty_124_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1075 = _GEN_12178 & tag_compare_valid_1 | dirty_124_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1076 = _GEN_12183 & _lru_T | dirty_125_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1077 = _GEN_12183 & tag_compare_valid_1 | dirty_125_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1078 = _GEN_12188 & _lru_T | dirty_126_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1079 = _GEN_12188 & tag_compare_valid_1 | dirty_126_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1080 = _GEN_12193 & _lru_T | dirty_127_0; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1081 = _GEN_12193 & tag_compare_valid_1 | dirty_127_1; // @[DCache.scala 313:{50,50} 69:22]
  wire  _GEN_1082 = io_cpu_M_mem_write ? _GEN_826 : dirty_0_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1083 = io_cpu_M_mem_write ? _GEN_827 : dirty_0_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1084 = io_cpu_M_mem_write ? _GEN_828 : dirty_1_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1085 = io_cpu_M_mem_write ? _GEN_829 : dirty_1_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1086 = io_cpu_M_mem_write ? _GEN_830 : dirty_2_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1087 = io_cpu_M_mem_write ? _GEN_831 : dirty_2_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1088 = io_cpu_M_mem_write ? _GEN_832 : dirty_3_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1089 = io_cpu_M_mem_write ? _GEN_833 : dirty_3_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1090 = io_cpu_M_mem_write ? _GEN_834 : dirty_4_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1091 = io_cpu_M_mem_write ? _GEN_835 : dirty_4_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1092 = io_cpu_M_mem_write ? _GEN_836 : dirty_5_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1093 = io_cpu_M_mem_write ? _GEN_837 : dirty_5_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1094 = io_cpu_M_mem_write ? _GEN_838 : dirty_6_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1095 = io_cpu_M_mem_write ? _GEN_839 : dirty_6_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1096 = io_cpu_M_mem_write ? _GEN_840 : dirty_7_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1097 = io_cpu_M_mem_write ? _GEN_841 : dirty_7_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1098 = io_cpu_M_mem_write ? _GEN_842 : dirty_8_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1099 = io_cpu_M_mem_write ? _GEN_843 : dirty_8_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1100 = io_cpu_M_mem_write ? _GEN_844 : dirty_9_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1101 = io_cpu_M_mem_write ? _GEN_845 : dirty_9_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1102 = io_cpu_M_mem_write ? _GEN_846 : dirty_10_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1103 = io_cpu_M_mem_write ? _GEN_847 : dirty_10_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1104 = io_cpu_M_mem_write ? _GEN_848 : dirty_11_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1105 = io_cpu_M_mem_write ? _GEN_849 : dirty_11_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1106 = io_cpu_M_mem_write ? _GEN_850 : dirty_12_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1107 = io_cpu_M_mem_write ? _GEN_851 : dirty_12_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1108 = io_cpu_M_mem_write ? _GEN_852 : dirty_13_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1109 = io_cpu_M_mem_write ? _GEN_853 : dirty_13_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1110 = io_cpu_M_mem_write ? _GEN_854 : dirty_14_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1111 = io_cpu_M_mem_write ? _GEN_855 : dirty_14_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1112 = io_cpu_M_mem_write ? _GEN_856 : dirty_15_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1113 = io_cpu_M_mem_write ? _GEN_857 : dirty_15_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1114 = io_cpu_M_mem_write ? _GEN_858 : dirty_16_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1115 = io_cpu_M_mem_write ? _GEN_859 : dirty_16_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1116 = io_cpu_M_mem_write ? _GEN_860 : dirty_17_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1117 = io_cpu_M_mem_write ? _GEN_861 : dirty_17_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1118 = io_cpu_M_mem_write ? _GEN_862 : dirty_18_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1119 = io_cpu_M_mem_write ? _GEN_863 : dirty_18_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1120 = io_cpu_M_mem_write ? _GEN_864 : dirty_19_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1121 = io_cpu_M_mem_write ? _GEN_865 : dirty_19_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1122 = io_cpu_M_mem_write ? _GEN_866 : dirty_20_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1123 = io_cpu_M_mem_write ? _GEN_867 : dirty_20_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1124 = io_cpu_M_mem_write ? _GEN_868 : dirty_21_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1125 = io_cpu_M_mem_write ? _GEN_869 : dirty_21_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1126 = io_cpu_M_mem_write ? _GEN_870 : dirty_22_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1127 = io_cpu_M_mem_write ? _GEN_871 : dirty_22_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1128 = io_cpu_M_mem_write ? _GEN_872 : dirty_23_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1129 = io_cpu_M_mem_write ? _GEN_873 : dirty_23_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1130 = io_cpu_M_mem_write ? _GEN_874 : dirty_24_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1131 = io_cpu_M_mem_write ? _GEN_875 : dirty_24_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1132 = io_cpu_M_mem_write ? _GEN_876 : dirty_25_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1133 = io_cpu_M_mem_write ? _GEN_877 : dirty_25_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1134 = io_cpu_M_mem_write ? _GEN_878 : dirty_26_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1135 = io_cpu_M_mem_write ? _GEN_879 : dirty_26_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1136 = io_cpu_M_mem_write ? _GEN_880 : dirty_27_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1137 = io_cpu_M_mem_write ? _GEN_881 : dirty_27_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1138 = io_cpu_M_mem_write ? _GEN_882 : dirty_28_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1139 = io_cpu_M_mem_write ? _GEN_883 : dirty_28_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1140 = io_cpu_M_mem_write ? _GEN_884 : dirty_29_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1141 = io_cpu_M_mem_write ? _GEN_885 : dirty_29_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1142 = io_cpu_M_mem_write ? _GEN_886 : dirty_30_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1143 = io_cpu_M_mem_write ? _GEN_887 : dirty_30_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1144 = io_cpu_M_mem_write ? _GEN_888 : dirty_31_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1145 = io_cpu_M_mem_write ? _GEN_889 : dirty_31_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1146 = io_cpu_M_mem_write ? _GEN_890 : dirty_32_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1147 = io_cpu_M_mem_write ? _GEN_891 : dirty_32_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1148 = io_cpu_M_mem_write ? _GEN_892 : dirty_33_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1149 = io_cpu_M_mem_write ? _GEN_893 : dirty_33_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1150 = io_cpu_M_mem_write ? _GEN_894 : dirty_34_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1151 = io_cpu_M_mem_write ? _GEN_895 : dirty_34_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1152 = io_cpu_M_mem_write ? _GEN_896 : dirty_35_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1153 = io_cpu_M_mem_write ? _GEN_897 : dirty_35_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1154 = io_cpu_M_mem_write ? _GEN_898 : dirty_36_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1155 = io_cpu_M_mem_write ? _GEN_899 : dirty_36_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1156 = io_cpu_M_mem_write ? _GEN_900 : dirty_37_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1157 = io_cpu_M_mem_write ? _GEN_901 : dirty_37_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1158 = io_cpu_M_mem_write ? _GEN_902 : dirty_38_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1159 = io_cpu_M_mem_write ? _GEN_903 : dirty_38_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1160 = io_cpu_M_mem_write ? _GEN_904 : dirty_39_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1161 = io_cpu_M_mem_write ? _GEN_905 : dirty_39_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1162 = io_cpu_M_mem_write ? _GEN_906 : dirty_40_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1163 = io_cpu_M_mem_write ? _GEN_907 : dirty_40_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1164 = io_cpu_M_mem_write ? _GEN_908 : dirty_41_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1165 = io_cpu_M_mem_write ? _GEN_909 : dirty_41_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1166 = io_cpu_M_mem_write ? _GEN_910 : dirty_42_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1167 = io_cpu_M_mem_write ? _GEN_911 : dirty_42_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1168 = io_cpu_M_mem_write ? _GEN_912 : dirty_43_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1169 = io_cpu_M_mem_write ? _GEN_913 : dirty_43_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1170 = io_cpu_M_mem_write ? _GEN_914 : dirty_44_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1171 = io_cpu_M_mem_write ? _GEN_915 : dirty_44_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1172 = io_cpu_M_mem_write ? _GEN_916 : dirty_45_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1173 = io_cpu_M_mem_write ? _GEN_917 : dirty_45_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1174 = io_cpu_M_mem_write ? _GEN_918 : dirty_46_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1175 = io_cpu_M_mem_write ? _GEN_919 : dirty_46_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1176 = io_cpu_M_mem_write ? _GEN_920 : dirty_47_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1177 = io_cpu_M_mem_write ? _GEN_921 : dirty_47_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1178 = io_cpu_M_mem_write ? _GEN_922 : dirty_48_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1179 = io_cpu_M_mem_write ? _GEN_923 : dirty_48_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1180 = io_cpu_M_mem_write ? _GEN_924 : dirty_49_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1181 = io_cpu_M_mem_write ? _GEN_925 : dirty_49_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1182 = io_cpu_M_mem_write ? _GEN_926 : dirty_50_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1183 = io_cpu_M_mem_write ? _GEN_927 : dirty_50_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1184 = io_cpu_M_mem_write ? _GEN_928 : dirty_51_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1185 = io_cpu_M_mem_write ? _GEN_929 : dirty_51_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1186 = io_cpu_M_mem_write ? _GEN_930 : dirty_52_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1187 = io_cpu_M_mem_write ? _GEN_931 : dirty_52_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1188 = io_cpu_M_mem_write ? _GEN_932 : dirty_53_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1189 = io_cpu_M_mem_write ? _GEN_933 : dirty_53_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1190 = io_cpu_M_mem_write ? _GEN_934 : dirty_54_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1191 = io_cpu_M_mem_write ? _GEN_935 : dirty_54_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1192 = io_cpu_M_mem_write ? _GEN_936 : dirty_55_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1193 = io_cpu_M_mem_write ? _GEN_937 : dirty_55_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1194 = io_cpu_M_mem_write ? _GEN_938 : dirty_56_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1195 = io_cpu_M_mem_write ? _GEN_939 : dirty_56_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1196 = io_cpu_M_mem_write ? _GEN_940 : dirty_57_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1197 = io_cpu_M_mem_write ? _GEN_941 : dirty_57_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1198 = io_cpu_M_mem_write ? _GEN_942 : dirty_58_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1199 = io_cpu_M_mem_write ? _GEN_943 : dirty_58_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1200 = io_cpu_M_mem_write ? _GEN_944 : dirty_59_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1201 = io_cpu_M_mem_write ? _GEN_945 : dirty_59_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1202 = io_cpu_M_mem_write ? _GEN_946 : dirty_60_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1203 = io_cpu_M_mem_write ? _GEN_947 : dirty_60_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1204 = io_cpu_M_mem_write ? _GEN_948 : dirty_61_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1205 = io_cpu_M_mem_write ? _GEN_949 : dirty_61_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1206 = io_cpu_M_mem_write ? _GEN_950 : dirty_62_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1207 = io_cpu_M_mem_write ? _GEN_951 : dirty_62_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1208 = io_cpu_M_mem_write ? _GEN_952 : dirty_63_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1209 = io_cpu_M_mem_write ? _GEN_953 : dirty_63_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1210 = io_cpu_M_mem_write ? _GEN_954 : dirty_64_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1211 = io_cpu_M_mem_write ? _GEN_955 : dirty_64_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1212 = io_cpu_M_mem_write ? _GEN_956 : dirty_65_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1213 = io_cpu_M_mem_write ? _GEN_957 : dirty_65_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1214 = io_cpu_M_mem_write ? _GEN_958 : dirty_66_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1215 = io_cpu_M_mem_write ? _GEN_959 : dirty_66_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1216 = io_cpu_M_mem_write ? _GEN_960 : dirty_67_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1217 = io_cpu_M_mem_write ? _GEN_961 : dirty_67_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1218 = io_cpu_M_mem_write ? _GEN_962 : dirty_68_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1219 = io_cpu_M_mem_write ? _GEN_963 : dirty_68_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1220 = io_cpu_M_mem_write ? _GEN_964 : dirty_69_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1221 = io_cpu_M_mem_write ? _GEN_965 : dirty_69_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1222 = io_cpu_M_mem_write ? _GEN_966 : dirty_70_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1223 = io_cpu_M_mem_write ? _GEN_967 : dirty_70_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1224 = io_cpu_M_mem_write ? _GEN_968 : dirty_71_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1225 = io_cpu_M_mem_write ? _GEN_969 : dirty_71_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1226 = io_cpu_M_mem_write ? _GEN_970 : dirty_72_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1227 = io_cpu_M_mem_write ? _GEN_971 : dirty_72_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1228 = io_cpu_M_mem_write ? _GEN_972 : dirty_73_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1229 = io_cpu_M_mem_write ? _GEN_973 : dirty_73_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1230 = io_cpu_M_mem_write ? _GEN_974 : dirty_74_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1231 = io_cpu_M_mem_write ? _GEN_975 : dirty_74_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1232 = io_cpu_M_mem_write ? _GEN_976 : dirty_75_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1233 = io_cpu_M_mem_write ? _GEN_977 : dirty_75_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1234 = io_cpu_M_mem_write ? _GEN_978 : dirty_76_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1235 = io_cpu_M_mem_write ? _GEN_979 : dirty_76_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1236 = io_cpu_M_mem_write ? _GEN_980 : dirty_77_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1237 = io_cpu_M_mem_write ? _GEN_981 : dirty_77_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1238 = io_cpu_M_mem_write ? _GEN_982 : dirty_78_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1239 = io_cpu_M_mem_write ? _GEN_983 : dirty_78_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1240 = io_cpu_M_mem_write ? _GEN_984 : dirty_79_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1241 = io_cpu_M_mem_write ? _GEN_985 : dirty_79_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1242 = io_cpu_M_mem_write ? _GEN_986 : dirty_80_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1243 = io_cpu_M_mem_write ? _GEN_987 : dirty_80_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1244 = io_cpu_M_mem_write ? _GEN_988 : dirty_81_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1245 = io_cpu_M_mem_write ? _GEN_989 : dirty_81_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1246 = io_cpu_M_mem_write ? _GEN_990 : dirty_82_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1247 = io_cpu_M_mem_write ? _GEN_991 : dirty_82_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1248 = io_cpu_M_mem_write ? _GEN_992 : dirty_83_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1249 = io_cpu_M_mem_write ? _GEN_993 : dirty_83_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1250 = io_cpu_M_mem_write ? _GEN_994 : dirty_84_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1251 = io_cpu_M_mem_write ? _GEN_995 : dirty_84_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1252 = io_cpu_M_mem_write ? _GEN_996 : dirty_85_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1253 = io_cpu_M_mem_write ? _GEN_997 : dirty_85_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1254 = io_cpu_M_mem_write ? _GEN_998 : dirty_86_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1255 = io_cpu_M_mem_write ? _GEN_999 : dirty_86_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1256 = io_cpu_M_mem_write ? _GEN_1000 : dirty_87_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1257 = io_cpu_M_mem_write ? _GEN_1001 : dirty_87_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1258 = io_cpu_M_mem_write ? _GEN_1002 : dirty_88_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1259 = io_cpu_M_mem_write ? _GEN_1003 : dirty_88_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1260 = io_cpu_M_mem_write ? _GEN_1004 : dirty_89_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1261 = io_cpu_M_mem_write ? _GEN_1005 : dirty_89_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1262 = io_cpu_M_mem_write ? _GEN_1006 : dirty_90_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1263 = io_cpu_M_mem_write ? _GEN_1007 : dirty_90_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1264 = io_cpu_M_mem_write ? _GEN_1008 : dirty_91_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1265 = io_cpu_M_mem_write ? _GEN_1009 : dirty_91_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1266 = io_cpu_M_mem_write ? _GEN_1010 : dirty_92_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1267 = io_cpu_M_mem_write ? _GEN_1011 : dirty_92_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1268 = io_cpu_M_mem_write ? _GEN_1012 : dirty_93_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1269 = io_cpu_M_mem_write ? _GEN_1013 : dirty_93_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1270 = io_cpu_M_mem_write ? _GEN_1014 : dirty_94_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1271 = io_cpu_M_mem_write ? _GEN_1015 : dirty_94_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1272 = io_cpu_M_mem_write ? _GEN_1016 : dirty_95_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1273 = io_cpu_M_mem_write ? _GEN_1017 : dirty_95_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1274 = io_cpu_M_mem_write ? _GEN_1018 : dirty_96_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1275 = io_cpu_M_mem_write ? _GEN_1019 : dirty_96_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1276 = io_cpu_M_mem_write ? _GEN_1020 : dirty_97_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1277 = io_cpu_M_mem_write ? _GEN_1021 : dirty_97_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1278 = io_cpu_M_mem_write ? _GEN_1022 : dirty_98_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1279 = io_cpu_M_mem_write ? _GEN_1023 : dirty_98_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1280 = io_cpu_M_mem_write ? _GEN_1024 : dirty_99_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1281 = io_cpu_M_mem_write ? _GEN_1025 : dirty_99_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1282 = io_cpu_M_mem_write ? _GEN_1026 : dirty_100_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1283 = io_cpu_M_mem_write ? _GEN_1027 : dirty_100_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1284 = io_cpu_M_mem_write ? _GEN_1028 : dirty_101_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1285 = io_cpu_M_mem_write ? _GEN_1029 : dirty_101_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1286 = io_cpu_M_mem_write ? _GEN_1030 : dirty_102_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1287 = io_cpu_M_mem_write ? _GEN_1031 : dirty_102_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1288 = io_cpu_M_mem_write ? _GEN_1032 : dirty_103_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1289 = io_cpu_M_mem_write ? _GEN_1033 : dirty_103_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1290 = io_cpu_M_mem_write ? _GEN_1034 : dirty_104_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1291 = io_cpu_M_mem_write ? _GEN_1035 : dirty_104_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1292 = io_cpu_M_mem_write ? _GEN_1036 : dirty_105_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1293 = io_cpu_M_mem_write ? _GEN_1037 : dirty_105_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1294 = io_cpu_M_mem_write ? _GEN_1038 : dirty_106_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1295 = io_cpu_M_mem_write ? _GEN_1039 : dirty_106_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1296 = io_cpu_M_mem_write ? _GEN_1040 : dirty_107_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1297 = io_cpu_M_mem_write ? _GEN_1041 : dirty_107_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1298 = io_cpu_M_mem_write ? _GEN_1042 : dirty_108_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1299 = io_cpu_M_mem_write ? _GEN_1043 : dirty_108_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1300 = io_cpu_M_mem_write ? _GEN_1044 : dirty_109_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1301 = io_cpu_M_mem_write ? _GEN_1045 : dirty_109_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1302 = io_cpu_M_mem_write ? _GEN_1046 : dirty_110_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1303 = io_cpu_M_mem_write ? _GEN_1047 : dirty_110_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1304 = io_cpu_M_mem_write ? _GEN_1048 : dirty_111_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1305 = io_cpu_M_mem_write ? _GEN_1049 : dirty_111_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1306 = io_cpu_M_mem_write ? _GEN_1050 : dirty_112_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1307 = io_cpu_M_mem_write ? _GEN_1051 : dirty_112_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1308 = io_cpu_M_mem_write ? _GEN_1052 : dirty_113_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1309 = io_cpu_M_mem_write ? _GEN_1053 : dirty_113_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1310 = io_cpu_M_mem_write ? _GEN_1054 : dirty_114_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1311 = io_cpu_M_mem_write ? _GEN_1055 : dirty_114_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1312 = io_cpu_M_mem_write ? _GEN_1056 : dirty_115_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1313 = io_cpu_M_mem_write ? _GEN_1057 : dirty_115_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1314 = io_cpu_M_mem_write ? _GEN_1058 : dirty_116_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1315 = io_cpu_M_mem_write ? _GEN_1059 : dirty_116_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1316 = io_cpu_M_mem_write ? _GEN_1060 : dirty_117_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1317 = io_cpu_M_mem_write ? _GEN_1061 : dirty_117_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1318 = io_cpu_M_mem_write ? _GEN_1062 : dirty_118_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1319 = io_cpu_M_mem_write ? _GEN_1063 : dirty_118_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1320 = io_cpu_M_mem_write ? _GEN_1064 : dirty_119_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1321 = io_cpu_M_mem_write ? _GEN_1065 : dirty_119_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1322 = io_cpu_M_mem_write ? _GEN_1066 : dirty_120_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1323 = io_cpu_M_mem_write ? _GEN_1067 : dirty_120_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1324 = io_cpu_M_mem_write ? _GEN_1068 : dirty_121_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1325 = io_cpu_M_mem_write ? _GEN_1069 : dirty_121_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1326 = io_cpu_M_mem_write ? _GEN_1070 : dirty_122_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1327 = io_cpu_M_mem_write ? _GEN_1071 : dirty_122_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1328 = io_cpu_M_mem_write ? _GEN_1072 : dirty_123_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1329 = io_cpu_M_mem_write ? _GEN_1073 : dirty_123_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1330 = io_cpu_M_mem_write ? _GEN_1074 : dirty_124_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1331 = io_cpu_M_mem_write ? _GEN_1075 : dirty_124_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1332 = io_cpu_M_mem_write ? _GEN_1076 : dirty_125_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1333 = io_cpu_M_mem_write ? _GEN_1077 : dirty_125_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1334 = io_cpu_M_mem_write ? _GEN_1078 : dirty_126_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1335 = io_cpu_M_mem_write ? _GEN_1079 : dirty_126_1; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1336 = io_cpu_M_mem_write ? _GEN_1080 : dirty_127_0; // @[DCache.scala 312:33 69:22]
  wire  _GEN_1337 = io_cpu_M_mem_write ? _GEN_1081 : dirty_127_1; // @[DCache.scala 312:33 69:22]
  wire [31:0] _GEN_1338 = io_cpu_stallM ? _GEN_1 : saved_rdata; // @[DCache.scala 141:28 315:28 316:29]
  wire [2:0] _GEN_1339 = io_cpu_stallM ? 3'h5 : state; // @[DCache.scala 315:28 317:29 65:96]
  wire  _GEN_1340 = _T_8 ? _GEN_698 : lru_0; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1341 = _T_8 ? _GEN_699 : lru_1; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1342 = _T_8 ? _GEN_700 : lru_2; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1343 = _T_8 ? _GEN_701 : lru_3; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1344 = _T_8 ? _GEN_702 : lru_4; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1345 = _T_8 ? _GEN_703 : lru_5; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1346 = _T_8 ? _GEN_704 : lru_6; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1347 = _T_8 ? _GEN_705 : lru_7; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1348 = _T_8 ? _GEN_706 : lru_8; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1349 = _T_8 ? _GEN_707 : lru_9; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1350 = _T_8 ? _GEN_708 : lru_10; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1351 = _T_8 ? _GEN_709 : lru_11; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1352 = _T_8 ? _GEN_710 : lru_12; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1353 = _T_8 ? _GEN_711 : lru_13; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1354 = _T_8 ? _GEN_712 : lru_14; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1355 = _T_8 ? _GEN_713 : lru_15; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1356 = _T_8 ? _GEN_714 : lru_16; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1357 = _T_8 ? _GEN_715 : lru_17; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1358 = _T_8 ? _GEN_716 : lru_18; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1359 = _T_8 ? _GEN_717 : lru_19; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1360 = _T_8 ? _GEN_718 : lru_20; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1361 = _T_8 ? _GEN_719 : lru_21; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1362 = _T_8 ? _GEN_720 : lru_22; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1363 = _T_8 ? _GEN_721 : lru_23; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1364 = _T_8 ? _GEN_722 : lru_24; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1365 = _T_8 ? _GEN_723 : lru_25; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1366 = _T_8 ? _GEN_724 : lru_26; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1367 = _T_8 ? _GEN_725 : lru_27; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1368 = _T_8 ? _GEN_726 : lru_28; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1369 = _T_8 ? _GEN_727 : lru_29; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1370 = _T_8 ? _GEN_728 : lru_30; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1371 = _T_8 ? _GEN_729 : lru_31; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1372 = _T_8 ? _GEN_730 : lru_32; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1373 = _T_8 ? _GEN_731 : lru_33; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1374 = _T_8 ? _GEN_732 : lru_34; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1375 = _T_8 ? _GEN_733 : lru_35; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1376 = _T_8 ? _GEN_734 : lru_36; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1377 = _T_8 ? _GEN_735 : lru_37; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1378 = _T_8 ? _GEN_736 : lru_38; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1379 = _T_8 ? _GEN_737 : lru_39; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1380 = _T_8 ? _GEN_738 : lru_40; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1381 = _T_8 ? _GEN_739 : lru_41; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1382 = _T_8 ? _GEN_740 : lru_42; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1383 = _T_8 ? _GEN_741 : lru_43; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1384 = _T_8 ? _GEN_742 : lru_44; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1385 = _T_8 ? _GEN_743 : lru_45; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1386 = _T_8 ? _GEN_744 : lru_46; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1387 = _T_8 ? _GEN_745 : lru_47; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1388 = _T_8 ? _GEN_746 : lru_48; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1389 = _T_8 ? _GEN_747 : lru_49; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1390 = _T_8 ? _GEN_748 : lru_50; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1391 = _T_8 ? _GEN_749 : lru_51; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1392 = _T_8 ? _GEN_750 : lru_52; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1393 = _T_8 ? _GEN_751 : lru_53; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1394 = _T_8 ? _GEN_752 : lru_54; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1395 = _T_8 ? _GEN_753 : lru_55; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1396 = _T_8 ? _GEN_754 : lru_56; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1397 = _T_8 ? _GEN_755 : lru_57; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1398 = _T_8 ? _GEN_756 : lru_58; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1399 = _T_8 ? _GEN_757 : lru_59; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1400 = _T_8 ? _GEN_758 : lru_60; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1401 = _T_8 ? _GEN_759 : lru_61; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1402 = _T_8 ? _GEN_760 : lru_62; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1403 = _T_8 ? _GEN_761 : lru_63; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1404 = _T_8 ? _GEN_762 : lru_64; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1405 = _T_8 ? _GEN_763 : lru_65; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1406 = _T_8 ? _GEN_764 : lru_66; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1407 = _T_8 ? _GEN_765 : lru_67; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1408 = _T_8 ? _GEN_766 : lru_68; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1409 = _T_8 ? _GEN_767 : lru_69; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1410 = _T_8 ? _GEN_768 : lru_70; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1411 = _T_8 ? _GEN_769 : lru_71; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1412 = _T_8 ? _GEN_770 : lru_72; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1413 = _T_8 ? _GEN_771 : lru_73; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1414 = _T_8 ? _GEN_772 : lru_74; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1415 = _T_8 ? _GEN_773 : lru_75; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1416 = _T_8 ? _GEN_774 : lru_76; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1417 = _T_8 ? _GEN_775 : lru_77; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1418 = _T_8 ? _GEN_776 : lru_78; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1419 = _T_8 ? _GEN_777 : lru_79; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1420 = _T_8 ? _GEN_778 : lru_80; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1421 = _T_8 ? _GEN_779 : lru_81; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1422 = _T_8 ? _GEN_780 : lru_82; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1423 = _T_8 ? _GEN_781 : lru_83; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1424 = _T_8 ? _GEN_782 : lru_84; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1425 = _T_8 ? _GEN_783 : lru_85; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1426 = _T_8 ? _GEN_784 : lru_86; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1427 = _T_8 ? _GEN_785 : lru_87; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1428 = _T_8 ? _GEN_786 : lru_88; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1429 = _T_8 ? _GEN_787 : lru_89; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1430 = _T_8 ? _GEN_788 : lru_90; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1431 = _T_8 ? _GEN_789 : lru_91; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1432 = _T_8 ? _GEN_790 : lru_92; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1433 = _T_8 ? _GEN_791 : lru_93; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1434 = _T_8 ? _GEN_792 : lru_94; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1435 = _T_8 ? _GEN_793 : lru_95; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1436 = _T_8 ? _GEN_794 : lru_96; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1437 = _T_8 ? _GEN_795 : lru_97; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1438 = _T_8 ? _GEN_796 : lru_98; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1439 = _T_8 ? _GEN_797 : lru_99; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1440 = _T_8 ? _GEN_798 : lru_100; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1441 = _T_8 ? _GEN_799 : lru_101; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1442 = _T_8 ? _GEN_800 : lru_102; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1443 = _T_8 ? _GEN_801 : lru_103; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1444 = _T_8 ? _GEN_802 : lru_104; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1445 = _T_8 ? _GEN_803 : lru_105; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1446 = _T_8 ? _GEN_804 : lru_106; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1447 = _T_8 ? _GEN_805 : lru_107; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1448 = _T_8 ? _GEN_806 : lru_108; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1449 = _T_8 ? _GEN_807 : lru_109; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1450 = _T_8 ? _GEN_808 : lru_110; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1451 = _T_8 ? _GEN_809 : lru_111; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1452 = _T_8 ? _GEN_810 : lru_112; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1453 = _T_8 ? _GEN_811 : lru_113; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1454 = _T_8 ? _GEN_812 : lru_114; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1455 = _T_8 ? _GEN_813 : lru_115; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1456 = _T_8 ? _GEN_814 : lru_116; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1457 = _T_8 ? _GEN_815 : lru_117; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1458 = _T_8 ? _GEN_816 : lru_118; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1459 = _T_8 ? _GEN_817 : lru_119; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1460 = _T_8 ? _GEN_818 : lru_120; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1461 = _T_8 ? _GEN_819 : lru_121; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1462 = _T_8 ? _GEN_820 : lru_122; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1463 = _T_8 ? _GEN_821 : lru_123; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1464 = _T_8 ? _GEN_822 : lru_124; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1465 = _T_8 ? _GEN_823 : lru_125; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1466 = _T_8 ? _GEN_824 : lru_126; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1467 = _T_8 ? _GEN_825 : lru_127; // @[DCache.scala 309:34 70:22]
  wire  _GEN_1468 = _T_8 ? _GEN_1082 : dirty_0_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1469 = _T_8 ? _GEN_1083 : dirty_0_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1470 = _T_8 ? _GEN_1084 : dirty_1_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1471 = _T_8 ? _GEN_1085 : dirty_1_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1472 = _T_8 ? _GEN_1086 : dirty_2_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1473 = _T_8 ? _GEN_1087 : dirty_2_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1474 = _T_8 ? _GEN_1088 : dirty_3_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1475 = _T_8 ? _GEN_1089 : dirty_3_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1476 = _T_8 ? _GEN_1090 : dirty_4_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1477 = _T_8 ? _GEN_1091 : dirty_4_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1478 = _T_8 ? _GEN_1092 : dirty_5_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1479 = _T_8 ? _GEN_1093 : dirty_5_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1480 = _T_8 ? _GEN_1094 : dirty_6_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1481 = _T_8 ? _GEN_1095 : dirty_6_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1482 = _T_8 ? _GEN_1096 : dirty_7_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1483 = _T_8 ? _GEN_1097 : dirty_7_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1484 = _T_8 ? _GEN_1098 : dirty_8_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1485 = _T_8 ? _GEN_1099 : dirty_8_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1486 = _T_8 ? _GEN_1100 : dirty_9_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1487 = _T_8 ? _GEN_1101 : dirty_9_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1488 = _T_8 ? _GEN_1102 : dirty_10_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1489 = _T_8 ? _GEN_1103 : dirty_10_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1490 = _T_8 ? _GEN_1104 : dirty_11_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1491 = _T_8 ? _GEN_1105 : dirty_11_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1492 = _T_8 ? _GEN_1106 : dirty_12_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1493 = _T_8 ? _GEN_1107 : dirty_12_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1494 = _T_8 ? _GEN_1108 : dirty_13_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1495 = _T_8 ? _GEN_1109 : dirty_13_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1496 = _T_8 ? _GEN_1110 : dirty_14_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1497 = _T_8 ? _GEN_1111 : dirty_14_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1498 = _T_8 ? _GEN_1112 : dirty_15_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1499 = _T_8 ? _GEN_1113 : dirty_15_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1500 = _T_8 ? _GEN_1114 : dirty_16_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1501 = _T_8 ? _GEN_1115 : dirty_16_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1502 = _T_8 ? _GEN_1116 : dirty_17_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1503 = _T_8 ? _GEN_1117 : dirty_17_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1504 = _T_8 ? _GEN_1118 : dirty_18_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1505 = _T_8 ? _GEN_1119 : dirty_18_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1506 = _T_8 ? _GEN_1120 : dirty_19_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1507 = _T_8 ? _GEN_1121 : dirty_19_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1508 = _T_8 ? _GEN_1122 : dirty_20_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1509 = _T_8 ? _GEN_1123 : dirty_20_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1510 = _T_8 ? _GEN_1124 : dirty_21_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1511 = _T_8 ? _GEN_1125 : dirty_21_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1512 = _T_8 ? _GEN_1126 : dirty_22_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1513 = _T_8 ? _GEN_1127 : dirty_22_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1514 = _T_8 ? _GEN_1128 : dirty_23_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1515 = _T_8 ? _GEN_1129 : dirty_23_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1516 = _T_8 ? _GEN_1130 : dirty_24_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1517 = _T_8 ? _GEN_1131 : dirty_24_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1518 = _T_8 ? _GEN_1132 : dirty_25_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1519 = _T_8 ? _GEN_1133 : dirty_25_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1520 = _T_8 ? _GEN_1134 : dirty_26_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1521 = _T_8 ? _GEN_1135 : dirty_26_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1522 = _T_8 ? _GEN_1136 : dirty_27_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1523 = _T_8 ? _GEN_1137 : dirty_27_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1524 = _T_8 ? _GEN_1138 : dirty_28_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1525 = _T_8 ? _GEN_1139 : dirty_28_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1526 = _T_8 ? _GEN_1140 : dirty_29_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1527 = _T_8 ? _GEN_1141 : dirty_29_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1528 = _T_8 ? _GEN_1142 : dirty_30_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1529 = _T_8 ? _GEN_1143 : dirty_30_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1530 = _T_8 ? _GEN_1144 : dirty_31_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1531 = _T_8 ? _GEN_1145 : dirty_31_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1532 = _T_8 ? _GEN_1146 : dirty_32_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1533 = _T_8 ? _GEN_1147 : dirty_32_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1534 = _T_8 ? _GEN_1148 : dirty_33_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1535 = _T_8 ? _GEN_1149 : dirty_33_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1536 = _T_8 ? _GEN_1150 : dirty_34_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1537 = _T_8 ? _GEN_1151 : dirty_34_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1538 = _T_8 ? _GEN_1152 : dirty_35_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1539 = _T_8 ? _GEN_1153 : dirty_35_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1540 = _T_8 ? _GEN_1154 : dirty_36_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1541 = _T_8 ? _GEN_1155 : dirty_36_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1542 = _T_8 ? _GEN_1156 : dirty_37_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1543 = _T_8 ? _GEN_1157 : dirty_37_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1544 = _T_8 ? _GEN_1158 : dirty_38_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1545 = _T_8 ? _GEN_1159 : dirty_38_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1546 = _T_8 ? _GEN_1160 : dirty_39_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1547 = _T_8 ? _GEN_1161 : dirty_39_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1548 = _T_8 ? _GEN_1162 : dirty_40_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1549 = _T_8 ? _GEN_1163 : dirty_40_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1550 = _T_8 ? _GEN_1164 : dirty_41_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1551 = _T_8 ? _GEN_1165 : dirty_41_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1552 = _T_8 ? _GEN_1166 : dirty_42_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1553 = _T_8 ? _GEN_1167 : dirty_42_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1554 = _T_8 ? _GEN_1168 : dirty_43_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1555 = _T_8 ? _GEN_1169 : dirty_43_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1556 = _T_8 ? _GEN_1170 : dirty_44_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1557 = _T_8 ? _GEN_1171 : dirty_44_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1558 = _T_8 ? _GEN_1172 : dirty_45_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1559 = _T_8 ? _GEN_1173 : dirty_45_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1560 = _T_8 ? _GEN_1174 : dirty_46_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1561 = _T_8 ? _GEN_1175 : dirty_46_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1562 = _T_8 ? _GEN_1176 : dirty_47_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1563 = _T_8 ? _GEN_1177 : dirty_47_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1564 = _T_8 ? _GEN_1178 : dirty_48_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1565 = _T_8 ? _GEN_1179 : dirty_48_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1566 = _T_8 ? _GEN_1180 : dirty_49_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1567 = _T_8 ? _GEN_1181 : dirty_49_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1568 = _T_8 ? _GEN_1182 : dirty_50_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1569 = _T_8 ? _GEN_1183 : dirty_50_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1570 = _T_8 ? _GEN_1184 : dirty_51_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1571 = _T_8 ? _GEN_1185 : dirty_51_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1572 = _T_8 ? _GEN_1186 : dirty_52_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1573 = _T_8 ? _GEN_1187 : dirty_52_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1574 = _T_8 ? _GEN_1188 : dirty_53_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1575 = _T_8 ? _GEN_1189 : dirty_53_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1576 = _T_8 ? _GEN_1190 : dirty_54_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1577 = _T_8 ? _GEN_1191 : dirty_54_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1578 = _T_8 ? _GEN_1192 : dirty_55_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1579 = _T_8 ? _GEN_1193 : dirty_55_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1580 = _T_8 ? _GEN_1194 : dirty_56_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1581 = _T_8 ? _GEN_1195 : dirty_56_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1582 = _T_8 ? _GEN_1196 : dirty_57_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1583 = _T_8 ? _GEN_1197 : dirty_57_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1584 = _T_8 ? _GEN_1198 : dirty_58_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1585 = _T_8 ? _GEN_1199 : dirty_58_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1586 = _T_8 ? _GEN_1200 : dirty_59_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1587 = _T_8 ? _GEN_1201 : dirty_59_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1588 = _T_8 ? _GEN_1202 : dirty_60_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1589 = _T_8 ? _GEN_1203 : dirty_60_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1590 = _T_8 ? _GEN_1204 : dirty_61_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1591 = _T_8 ? _GEN_1205 : dirty_61_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1592 = _T_8 ? _GEN_1206 : dirty_62_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1593 = _T_8 ? _GEN_1207 : dirty_62_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1594 = _T_8 ? _GEN_1208 : dirty_63_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1595 = _T_8 ? _GEN_1209 : dirty_63_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1596 = _T_8 ? _GEN_1210 : dirty_64_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1597 = _T_8 ? _GEN_1211 : dirty_64_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1598 = _T_8 ? _GEN_1212 : dirty_65_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1599 = _T_8 ? _GEN_1213 : dirty_65_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1600 = _T_8 ? _GEN_1214 : dirty_66_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1601 = _T_8 ? _GEN_1215 : dirty_66_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1602 = _T_8 ? _GEN_1216 : dirty_67_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1603 = _T_8 ? _GEN_1217 : dirty_67_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1604 = _T_8 ? _GEN_1218 : dirty_68_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1605 = _T_8 ? _GEN_1219 : dirty_68_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1606 = _T_8 ? _GEN_1220 : dirty_69_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1607 = _T_8 ? _GEN_1221 : dirty_69_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1608 = _T_8 ? _GEN_1222 : dirty_70_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1609 = _T_8 ? _GEN_1223 : dirty_70_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1610 = _T_8 ? _GEN_1224 : dirty_71_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1611 = _T_8 ? _GEN_1225 : dirty_71_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1612 = _T_8 ? _GEN_1226 : dirty_72_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1613 = _T_8 ? _GEN_1227 : dirty_72_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1614 = _T_8 ? _GEN_1228 : dirty_73_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1615 = _T_8 ? _GEN_1229 : dirty_73_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1616 = _T_8 ? _GEN_1230 : dirty_74_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1617 = _T_8 ? _GEN_1231 : dirty_74_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1618 = _T_8 ? _GEN_1232 : dirty_75_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1619 = _T_8 ? _GEN_1233 : dirty_75_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1620 = _T_8 ? _GEN_1234 : dirty_76_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1621 = _T_8 ? _GEN_1235 : dirty_76_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1622 = _T_8 ? _GEN_1236 : dirty_77_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1623 = _T_8 ? _GEN_1237 : dirty_77_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1624 = _T_8 ? _GEN_1238 : dirty_78_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1625 = _T_8 ? _GEN_1239 : dirty_78_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1626 = _T_8 ? _GEN_1240 : dirty_79_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1627 = _T_8 ? _GEN_1241 : dirty_79_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1628 = _T_8 ? _GEN_1242 : dirty_80_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1629 = _T_8 ? _GEN_1243 : dirty_80_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1630 = _T_8 ? _GEN_1244 : dirty_81_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1631 = _T_8 ? _GEN_1245 : dirty_81_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1632 = _T_8 ? _GEN_1246 : dirty_82_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1633 = _T_8 ? _GEN_1247 : dirty_82_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1634 = _T_8 ? _GEN_1248 : dirty_83_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1635 = _T_8 ? _GEN_1249 : dirty_83_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1636 = _T_8 ? _GEN_1250 : dirty_84_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1637 = _T_8 ? _GEN_1251 : dirty_84_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1638 = _T_8 ? _GEN_1252 : dirty_85_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1639 = _T_8 ? _GEN_1253 : dirty_85_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1640 = _T_8 ? _GEN_1254 : dirty_86_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1641 = _T_8 ? _GEN_1255 : dirty_86_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1642 = _T_8 ? _GEN_1256 : dirty_87_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1643 = _T_8 ? _GEN_1257 : dirty_87_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1644 = _T_8 ? _GEN_1258 : dirty_88_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1645 = _T_8 ? _GEN_1259 : dirty_88_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1646 = _T_8 ? _GEN_1260 : dirty_89_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1647 = _T_8 ? _GEN_1261 : dirty_89_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1648 = _T_8 ? _GEN_1262 : dirty_90_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1649 = _T_8 ? _GEN_1263 : dirty_90_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1650 = _T_8 ? _GEN_1264 : dirty_91_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1651 = _T_8 ? _GEN_1265 : dirty_91_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1652 = _T_8 ? _GEN_1266 : dirty_92_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1653 = _T_8 ? _GEN_1267 : dirty_92_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1654 = _T_8 ? _GEN_1268 : dirty_93_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1655 = _T_8 ? _GEN_1269 : dirty_93_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1656 = _T_8 ? _GEN_1270 : dirty_94_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1657 = _T_8 ? _GEN_1271 : dirty_94_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1658 = _T_8 ? _GEN_1272 : dirty_95_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1659 = _T_8 ? _GEN_1273 : dirty_95_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1660 = _T_8 ? _GEN_1274 : dirty_96_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1661 = _T_8 ? _GEN_1275 : dirty_96_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1662 = _T_8 ? _GEN_1276 : dirty_97_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1663 = _T_8 ? _GEN_1277 : dirty_97_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1664 = _T_8 ? _GEN_1278 : dirty_98_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1665 = _T_8 ? _GEN_1279 : dirty_98_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1666 = _T_8 ? _GEN_1280 : dirty_99_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1667 = _T_8 ? _GEN_1281 : dirty_99_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1668 = _T_8 ? _GEN_1282 : dirty_100_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1669 = _T_8 ? _GEN_1283 : dirty_100_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1670 = _T_8 ? _GEN_1284 : dirty_101_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1671 = _T_8 ? _GEN_1285 : dirty_101_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1672 = _T_8 ? _GEN_1286 : dirty_102_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1673 = _T_8 ? _GEN_1287 : dirty_102_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1674 = _T_8 ? _GEN_1288 : dirty_103_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1675 = _T_8 ? _GEN_1289 : dirty_103_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1676 = _T_8 ? _GEN_1290 : dirty_104_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1677 = _T_8 ? _GEN_1291 : dirty_104_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1678 = _T_8 ? _GEN_1292 : dirty_105_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1679 = _T_8 ? _GEN_1293 : dirty_105_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1680 = _T_8 ? _GEN_1294 : dirty_106_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1681 = _T_8 ? _GEN_1295 : dirty_106_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1682 = _T_8 ? _GEN_1296 : dirty_107_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1683 = _T_8 ? _GEN_1297 : dirty_107_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1684 = _T_8 ? _GEN_1298 : dirty_108_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1685 = _T_8 ? _GEN_1299 : dirty_108_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1686 = _T_8 ? _GEN_1300 : dirty_109_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1687 = _T_8 ? _GEN_1301 : dirty_109_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1688 = _T_8 ? _GEN_1302 : dirty_110_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1689 = _T_8 ? _GEN_1303 : dirty_110_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1690 = _T_8 ? _GEN_1304 : dirty_111_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1691 = _T_8 ? _GEN_1305 : dirty_111_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1692 = _T_8 ? _GEN_1306 : dirty_112_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1693 = _T_8 ? _GEN_1307 : dirty_112_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1694 = _T_8 ? _GEN_1308 : dirty_113_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1695 = _T_8 ? _GEN_1309 : dirty_113_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1696 = _T_8 ? _GEN_1310 : dirty_114_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1697 = _T_8 ? _GEN_1311 : dirty_114_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1698 = _T_8 ? _GEN_1312 : dirty_115_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1699 = _T_8 ? _GEN_1313 : dirty_115_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1700 = _T_8 ? _GEN_1314 : dirty_116_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1701 = _T_8 ? _GEN_1315 : dirty_116_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1702 = _T_8 ? _GEN_1316 : dirty_117_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1703 = _T_8 ? _GEN_1317 : dirty_117_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1704 = _T_8 ? _GEN_1318 : dirty_118_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1705 = _T_8 ? _GEN_1319 : dirty_118_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1706 = _T_8 ? _GEN_1320 : dirty_119_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1707 = _T_8 ? _GEN_1321 : dirty_119_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1708 = _T_8 ? _GEN_1322 : dirty_120_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1709 = _T_8 ? _GEN_1323 : dirty_120_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1710 = _T_8 ? _GEN_1324 : dirty_121_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1711 = _T_8 ? _GEN_1325 : dirty_121_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1712 = _T_8 ? _GEN_1326 : dirty_122_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1713 = _T_8 ? _GEN_1327 : dirty_122_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1714 = _T_8 ? _GEN_1328 : dirty_123_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1715 = _T_8 ? _GEN_1329 : dirty_123_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1716 = _T_8 ? _GEN_1330 : dirty_124_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1717 = _T_8 ? _GEN_1331 : dirty_124_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1718 = _T_8 ? _GEN_1332 : dirty_125_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1719 = _T_8 ? _GEN_1333 : dirty_125_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1720 = _T_8 ? _GEN_1334 : dirty_126_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1721 = _T_8 ? _GEN_1335 : dirty_126_1; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1722 = _T_8 ? _GEN_1336 : dirty_127_0; // @[DCache.scala 309:34 69:22]
  wire  _GEN_1723 = _T_8 ? _GEN_1337 : dirty_127_1; // @[DCache.scala 309:34 69:22]
  wire [31:0] _GEN_1724 = _T_8 ? _GEN_1338 : saved_rdata; // @[DCache.scala 141:28 309:34]
  wire [2:0] _GEN_1725 = _T_8 ? _GEN_1339 : state; // @[DCache.scala 309:34 65:96]
  wire [2:0] _GEN_1726 = _cached_stall_T_1 ? 3'h4 : _GEN_1725; // @[DCache.scala 298:28 299:37]
  wire [3:0] _GEN_1727 = _cached_stall_T_1 ? 4'h0 : axi_wcnt; // @[DCache.scala 298:28 300:37 89:40]
  wire [9:0] _GEN_1728 = _cached_stall_T_1 ? _bram_replace_addr_T : bram_replace_addr; // @[DCache.scala 298:28 301:37 90:40]
  wire [9:0] _GEN_1729 = _cached_stall_T_1 ? _bram_replace_addr_T : bram_read_ready_addr; // @[DCache.scala 298:28 302:37 91:40]
  wire [9:0] _GEN_1730 = _cached_stall_T_1 ? _bram_replace_addr_T : bram_replace_write_addr; // @[DCache.scala 298:28 303:37 92:40]
  wire  _GEN_1732 = _cached_stall_T_1 | bram_use_replace_addr; // @[DCache.scala 298:28 305:37 95:40]
  wire  _GEN_1734 = _cached_stall_T_1 ? _GEN_697 : replace_writeback; // @[DCache.scala 298:28 307:37 101:40]
  wire  _GEN_1735 = _cached_stall_T_1 ? lru_0 : _GEN_1340; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1736 = _cached_stall_T_1 ? lru_1 : _GEN_1341; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1737 = _cached_stall_T_1 ? lru_2 : _GEN_1342; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1738 = _cached_stall_T_1 ? lru_3 : _GEN_1343; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1739 = _cached_stall_T_1 ? lru_4 : _GEN_1344; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1740 = _cached_stall_T_1 ? lru_5 : _GEN_1345; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1741 = _cached_stall_T_1 ? lru_6 : _GEN_1346; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1742 = _cached_stall_T_1 ? lru_7 : _GEN_1347; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1743 = _cached_stall_T_1 ? lru_8 : _GEN_1348; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1744 = _cached_stall_T_1 ? lru_9 : _GEN_1349; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1745 = _cached_stall_T_1 ? lru_10 : _GEN_1350; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1746 = _cached_stall_T_1 ? lru_11 : _GEN_1351; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1747 = _cached_stall_T_1 ? lru_12 : _GEN_1352; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1748 = _cached_stall_T_1 ? lru_13 : _GEN_1353; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1749 = _cached_stall_T_1 ? lru_14 : _GEN_1354; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1750 = _cached_stall_T_1 ? lru_15 : _GEN_1355; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1751 = _cached_stall_T_1 ? lru_16 : _GEN_1356; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1752 = _cached_stall_T_1 ? lru_17 : _GEN_1357; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1753 = _cached_stall_T_1 ? lru_18 : _GEN_1358; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1754 = _cached_stall_T_1 ? lru_19 : _GEN_1359; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1755 = _cached_stall_T_1 ? lru_20 : _GEN_1360; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1756 = _cached_stall_T_1 ? lru_21 : _GEN_1361; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1757 = _cached_stall_T_1 ? lru_22 : _GEN_1362; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1758 = _cached_stall_T_1 ? lru_23 : _GEN_1363; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1759 = _cached_stall_T_1 ? lru_24 : _GEN_1364; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1760 = _cached_stall_T_1 ? lru_25 : _GEN_1365; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1761 = _cached_stall_T_1 ? lru_26 : _GEN_1366; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1762 = _cached_stall_T_1 ? lru_27 : _GEN_1367; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1763 = _cached_stall_T_1 ? lru_28 : _GEN_1368; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1764 = _cached_stall_T_1 ? lru_29 : _GEN_1369; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1765 = _cached_stall_T_1 ? lru_30 : _GEN_1370; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1766 = _cached_stall_T_1 ? lru_31 : _GEN_1371; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1767 = _cached_stall_T_1 ? lru_32 : _GEN_1372; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1768 = _cached_stall_T_1 ? lru_33 : _GEN_1373; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1769 = _cached_stall_T_1 ? lru_34 : _GEN_1374; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1770 = _cached_stall_T_1 ? lru_35 : _GEN_1375; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1771 = _cached_stall_T_1 ? lru_36 : _GEN_1376; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1772 = _cached_stall_T_1 ? lru_37 : _GEN_1377; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1773 = _cached_stall_T_1 ? lru_38 : _GEN_1378; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1774 = _cached_stall_T_1 ? lru_39 : _GEN_1379; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1775 = _cached_stall_T_1 ? lru_40 : _GEN_1380; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1776 = _cached_stall_T_1 ? lru_41 : _GEN_1381; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1777 = _cached_stall_T_1 ? lru_42 : _GEN_1382; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1778 = _cached_stall_T_1 ? lru_43 : _GEN_1383; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1779 = _cached_stall_T_1 ? lru_44 : _GEN_1384; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1780 = _cached_stall_T_1 ? lru_45 : _GEN_1385; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1781 = _cached_stall_T_1 ? lru_46 : _GEN_1386; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1782 = _cached_stall_T_1 ? lru_47 : _GEN_1387; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1783 = _cached_stall_T_1 ? lru_48 : _GEN_1388; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1784 = _cached_stall_T_1 ? lru_49 : _GEN_1389; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1785 = _cached_stall_T_1 ? lru_50 : _GEN_1390; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1786 = _cached_stall_T_1 ? lru_51 : _GEN_1391; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1787 = _cached_stall_T_1 ? lru_52 : _GEN_1392; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1788 = _cached_stall_T_1 ? lru_53 : _GEN_1393; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1789 = _cached_stall_T_1 ? lru_54 : _GEN_1394; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1790 = _cached_stall_T_1 ? lru_55 : _GEN_1395; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1791 = _cached_stall_T_1 ? lru_56 : _GEN_1396; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1792 = _cached_stall_T_1 ? lru_57 : _GEN_1397; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1793 = _cached_stall_T_1 ? lru_58 : _GEN_1398; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1794 = _cached_stall_T_1 ? lru_59 : _GEN_1399; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1795 = _cached_stall_T_1 ? lru_60 : _GEN_1400; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1796 = _cached_stall_T_1 ? lru_61 : _GEN_1401; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1797 = _cached_stall_T_1 ? lru_62 : _GEN_1402; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1798 = _cached_stall_T_1 ? lru_63 : _GEN_1403; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1799 = _cached_stall_T_1 ? lru_64 : _GEN_1404; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1800 = _cached_stall_T_1 ? lru_65 : _GEN_1405; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1801 = _cached_stall_T_1 ? lru_66 : _GEN_1406; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1802 = _cached_stall_T_1 ? lru_67 : _GEN_1407; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1803 = _cached_stall_T_1 ? lru_68 : _GEN_1408; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1804 = _cached_stall_T_1 ? lru_69 : _GEN_1409; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1805 = _cached_stall_T_1 ? lru_70 : _GEN_1410; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1806 = _cached_stall_T_1 ? lru_71 : _GEN_1411; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1807 = _cached_stall_T_1 ? lru_72 : _GEN_1412; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1808 = _cached_stall_T_1 ? lru_73 : _GEN_1413; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1809 = _cached_stall_T_1 ? lru_74 : _GEN_1414; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1810 = _cached_stall_T_1 ? lru_75 : _GEN_1415; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1811 = _cached_stall_T_1 ? lru_76 : _GEN_1416; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1812 = _cached_stall_T_1 ? lru_77 : _GEN_1417; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1813 = _cached_stall_T_1 ? lru_78 : _GEN_1418; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1814 = _cached_stall_T_1 ? lru_79 : _GEN_1419; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1815 = _cached_stall_T_1 ? lru_80 : _GEN_1420; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1816 = _cached_stall_T_1 ? lru_81 : _GEN_1421; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1817 = _cached_stall_T_1 ? lru_82 : _GEN_1422; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1818 = _cached_stall_T_1 ? lru_83 : _GEN_1423; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1819 = _cached_stall_T_1 ? lru_84 : _GEN_1424; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1820 = _cached_stall_T_1 ? lru_85 : _GEN_1425; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1821 = _cached_stall_T_1 ? lru_86 : _GEN_1426; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1822 = _cached_stall_T_1 ? lru_87 : _GEN_1427; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1823 = _cached_stall_T_1 ? lru_88 : _GEN_1428; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1824 = _cached_stall_T_1 ? lru_89 : _GEN_1429; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1825 = _cached_stall_T_1 ? lru_90 : _GEN_1430; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1826 = _cached_stall_T_1 ? lru_91 : _GEN_1431; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1827 = _cached_stall_T_1 ? lru_92 : _GEN_1432; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1828 = _cached_stall_T_1 ? lru_93 : _GEN_1433; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1829 = _cached_stall_T_1 ? lru_94 : _GEN_1434; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1830 = _cached_stall_T_1 ? lru_95 : _GEN_1435; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1831 = _cached_stall_T_1 ? lru_96 : _GEN_1436; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1832 = _cached_stall_T_1 ? lru_97 : _GEN_1437; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1833 = _cached_stall_T_1 ? lru_98 : _GEN_1438; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1834 = _cached_stall_T_1 ? lru_99 : _GEN_1439; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1835 = _cached_stall_T_1 ? lru_100 : _GEN_1440; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1836 = _cached_stall_T_1 ? lru_101 : _GEN_1441; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1837 = _cached_stall_T_1 ? lru_102 : _GEN_1442; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1838 = _cached_stall_T_1 ? lru_103 : _GEN_1443; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1839 = _cached_stall_T_1 ? lru_104 : _GEN_1444; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1840 = _cached_stall_T_1 ? lru_105 : _GEN_1445; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1841 = _cached_stall_T_1 ? lru_106 : _GEN_1446; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1842 = _cached_stall_T_1 ? lru_107 : _GEN_1447; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1843 = _cached_stall_T_1 ? lru_108 : _GEN_1448; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1844 = _cached_stall_T_1 ? lru_109 : _GEN_1449; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1845 = _cached_stall_T_1 ? lru_110 : _GEN_1450; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1846 = _cached_stall_T_1 ? lru_111 : _GEN_1451; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1847 = _cached_stall_T_1 ? lru_112 : _GEN_1452; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1848 = _cached_stall_T_1 ? lru_113 : _GEN_1453; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1849 = _cached_stall_T_1 ? lru_114 : _GEN_1454; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1850 = _cached_stall_T_1 ? lru_115 : _GEN_1455; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1851 = _cached_stall_T_1 ? lru_116 : _GEN_1456; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1852 = _cached_stall_T_1 ? lru_117 : _GEN_1457; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1853 = _cached_stall_T_1 ? lru_118 : _GEN_1458; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1854 = _cached_stall_T_1 ? lru_119 : _GEN_1459; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1855 = _cached_stall_T_1 ? lru_120 : _GEN_1460; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1856 = _cached_stall_T_1 ? lru_121 : _GEN_1461; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1857 = _cached_stall_T_1 ? lru_122 : _GEN_1462; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1858 = _cached_stall_T_1 ? lru_123 : _GEN_1463; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1859 = _cached_stall_T_1 ? lru_124 : _GEN_1464; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1860 = _cached_stall_T_1 ? lru_125 : _GEN_1465; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1861 = _cached_stall_T_1 ? lru_126 : _GEN_1466; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1862 = _cached_stall_T_1 ? lru_127 : _GEN_1467; // @[DCache.scala 298:28 70:22]
  wire  _GEN_1863 = _cached_stall_T_1 ? dirty_0_0 : _GEN_1468; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1864 = _cached_stall_T_1 ? dirty_0_1 : _GEN_1469; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1865 = _cached_stall_T_1 ? dirty_1_0 : _GEN_1470; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1866 = _cached_stall_T_1 ? dirty_1_1 : _GEN_1471; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1867 = _cached_stall_T_1 ? dirty_2_0 : _GEN_1472; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1868 = _cached_stall_T_1 ? dirty_2_1 : _GEN_1473; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1869 = _cached_stall_T_1 ? dirty_3_0 : _GEN_1474; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1870 = _cached_stall_T_1 ? dirty_3_1 : _GEN_1475; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1871 = _cached_stall_T_1 ? dirty_4_0 : _GEN_1476; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1872 = _cached_stall_T_1 ? dirty_4_1 : _GEN_1477; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1873 = _cached_stall_T_1 ? dirty_5_0 : _GEN_1478; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1874 = _cached_stall_T_1 ? dirty_5_1 : _GEN_1479; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1875 = _cached_stall_T_1 ? dirty_6_0 : _GEN_1480; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1876 = _cached_stall_T_1 ? dirty_6_1 : _GEN_1481; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1877 = _cached_stall_T_1 ? dirty_7_0 : _GEN_1482; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1878 = _cached_stall_T_1 ? dirty_7_1 : _GEN_1483; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1879 = _cached_stall_T_1 ? dirty_8_0 : _GEN_1484; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1880 = _cached_stall_T_1 ? dirty_8_1 : _GEN_1485; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1881 = _cached_stall_T_1 ? dirty_9_0 : _GEN_1486; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1882 = _cached_stall_T_1 ? dirty_9_1 : _GEN_1487; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1883 = _cached_stall_T_1 ? dirty_10_0 : _GEN_1488; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1884 = _cached_stall_T_1 ? dirty_10_1 : _GEN_1489; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1885 = _cached_stall_T_1 ? dirty_11_0 : _GEN_1490; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1886 = _cached_stall_T_1 ? dirty_11_1 : _GEN_1491; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1887 = _cached_stall_T_1 ? dirty_12_0 : _GEN_1492; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1888 = _cached_stall_T_1 ? dirty_12_1 : _GEN_1493; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1889 = _cached_stall_T_1 ? dirty_13_0 : _GEN_1494; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1890 = _cached_stall_T_1 ? dirty_13_1 : _GEN_1495; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1891 = _cached_stall_T_1 ? dirty_14_0 : _GEN_1496; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1892 = _cached_stall_T_1 ? dirty_14_1 : _GEN_1497; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1893 = _cached_stall_T_1 ? dirty_15_0 : _GEN_1498; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1894 = _cached_stall_T_1 ? dirty_15_1 : _GEN_1499; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1895 = _cached_stall_T_1 ? dirty_16_0 : _GEN_1500; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1896 = _cached_stall_T_1 ? dirty_16_1 : _GEN_1501; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1897 = _cached_stall_T_1 ? dirty_17_0 : _GEN_1502; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1898 = _cached_stall_T_1 ? dirty_17_1 : _GEN_1503; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1899 = _cached_stall_T_1 ? dirty_18_0 : _GEN_1504; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1900 = _cached_stall_T_1 ? dirty_18_1 : _GEN_1505; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1901 = _cached_stall_T_1 ? dirty_19_0 : _GEN_1506; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1902 = _cached_stall_T_1 ? dirty_19_1 : _GEN_1507; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1903 = _cached_stall_T_1 ? dirty_20_0 : _GEN_1508; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1904 = _cached_stall_T_1 ? dirty_20_1 : _GEN_1509; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1905 = _cached_stall_T_1 ? dirty_21_0 : _GEN_1510; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1906 = _cached_stall_T_1 ? dirty_21_1 : _GEN_1511; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1907 = _cached_stall_T_1 ? dirty_22_0 : _GEN_1512; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1908 = _cached_stall_T_1 ? dirty_22_1 : _GEN_1513; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1909 = _cached_stall_T_1 ? dirty_23_0 : _GEN_1514; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1910 = _cached_stall_T_1 ? dirty_23_1 : _GEN_1515; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1911 = _cached_stall_T_1 ? dirty_24_0 : _GEN_1516; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1912 = _cached_stall_T_1 ? dirty_24_1 : _GEN_1517; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1913 = _cached_stall_T_1 ? dirty_25_0 : _GEN_1518; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1914 = _cached_stall_T_1 ? dirty_25_1 : _GEN_1519; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1915 = _cached_stall_T_1 ? dirty_26_0 : _GEN_1520; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1916 = _cached_stall_T_1 ? dirty_26_1 : _GEN_1521; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1917 = _cached_stall_T_1 ? dirty_27_0 : _GEN_1522; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1918 = _cached_stall_T_1 ? dirty_27_1 : _GEN_1523; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1919 = _cached_stall_T_1 ? dirty_28_0 : _GEN_1524; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1920 = _cached_stall_T_1 ? dirty_28_1 : _GEN_1525; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1921 = _cached_stall_T_1 ? dirty_29_0 : _GEN_1526; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1922 = _cached_stall_T_1 ? dirty_29_1 : _GEN_1527; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1923 = _cached_stall_T_1 ? dirty_30_0 : _GEN_1528; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1924 = _cached_stall_T_1 ? dirty_30_1 : _GEN_1529; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1925 = _cached_stall_T_1 ? dirty_31_0 : _GEN_1530; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1926 = _cached_stall_T_1 ? dirty_31_1 : _GEN_1531; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1927 = _cached_stall_T_1 ? dirty_32_0 : _GEN_1532; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1928 = _cached_stall_T_1 ? dirty_32_1 : _GEN_1533; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1929 = _cached_stall_T_1 ? dirty_33_0 : _GEN_1534; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1930 = _cached_stall_T_1 ? dirty_33_1 : _GEN_1535; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1931 = _cached_stall_T_1 ? dirty_34_0 : _GEN_1536; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1932 = _cached_stall_T_1 ? dirty_34_1 : _GEN_1537; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1933 = _cached_stall_T_1 ? dirty_35_0 : _GEN_1538; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1934 = _cached_stall_T_1 ? dirty_35_1 : _GEN_1539; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1935 = _cached_stall_T_1 ? dirty_36_0 : _GEN_1540; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1936 = _cached_stall_T_1 ? dirty_36_1 : _GEN_1541; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1937 = _cached_stall_T_1 ? dirty_37_0 : _GEN_1542; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1938 = _cached_stall_T_1 ? dirty_37_1 : _GEN_1543; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1939 = _cached_stall_T_1 ? dirty_38_0 : _GEN_1544; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1940 = _cached_stall_T_1 ? dirty_38_1 : _GEN_1545; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1941 = _cached_stall_T_1 ? dirty_39_0 : _GEN_1546; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1942 = _cached_stall_T_1 ? dirty_39_1 : _GEN_1547; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1943 = _cached_stall_T_1 ? dirty_40_0 : _GEN_1548; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1944 = _cached_stall_T_1 ? dirty_40_1 : _GEN_1549; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1945 = _cached_stall_T_1 ? dirty_41_0 : _GEN_1550; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1946 = _cached_stall_T_1 ? dirty_41_1 : _GEN_1551; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1947 = _cached_stall_T_1 ? dirty_42_0 : _GEN_1552; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1948 = _cached_stall_T_1 ? dirty_42_1 : _GEN_1553; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1949 = _cached_stall_T_1 ? dirty_43_0 : _GEN_1554; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1950 = _cached_stall_T_1 ? dirty_43_1 : _GEN_1555; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1951 = _cached_stall_T_1 ? dirty_44_0 : _GEN_1556; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1952 = _cached_stall_T_1 ? dirty_44_1 : _GEN_1557; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1953 = _cached_stall_T_1 ? dirty_45_0 : _GEN_1558; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1954 = _cached_stall_T_1 ? dirty_45_1 : _GEN_1559; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1955 = _cached_stall_T_1 ? dirty_46_0 : _GEN_1560; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1956 = _cached_stall_T_1 ? dirty_46_1 : _GEN_1561; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1957 = _cached_stall_T_1 ? dirty_47_0 : _GEN_1562; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1958 = _cached_stall_T_1 ? dirty_47_1 : _GEN_1563; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1959 = _cached_stall_T_1 ? dirty_48_0 : _GEN_1564; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1960 = _cached_stall_T_1 ? dirty_48_1 : _GEN_1565; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1961 = _cached_stall_T_1 ? dirty_49_0 : _GEN_1566; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1962 = _cached_stall_T_1 ? dirty_49_1 : _GEN_1567; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1963 = _cached_stall_T_1 ? dirty_50_0 : _GEN_1568; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1964 = _cached_stall_T_1 ? dirty_50_1 : _GEN_1569; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1965 = _cached_stall_T_1 ? dirty_51_0 : _GEN_1570; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1966 = _cached_stall_T_1 ? dirty_51_1 : _GEN_1571; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1967 = _cached_stall_T_1 ? dirty_52_0 : _GEN_1572; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1968 = _cached_stall_T_1 ? dirty_52_1 : _GEN_1573; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1969 = _cached_stall_T_1 ? dirty_53_0 : _GEN_1574; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1970 = _cached_stall_T_1 ? dirty_53_1 : _GEN_1575; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1971 = _cached_stall_T_1 ? dirty_54_0 : _GEN_1576; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1972 = _cached_stall_T_1 ? dirty_54_1 : _GEN_1577; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1973 = _cached_stall_T_1 ? dirty_55_0 : _GEN_1578; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1974 = _cached_stall_T_1 ? dirty_55_1 : _GEN_1579; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1975 = _cached_stall_T_1 ? dirty_56_0 : _GEN_1580; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1976 = _cached_stall_T_1 ? dirty_56_1 : _GEN_1581; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1977 = _cached_stall_T_1 ? dirty_57_0 : _GEN_1582; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1978 = _cached_stall_T_1 ? dirty_57_1 : _GEN_1583; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1979 = _cached_stall_T_1 ? dirty_58_0 : _GEN_1584; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1980 = _cached_stall_T_1 ? dirty_58_1 : _GEN_1585; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1981 = _cached_stall_T_1 ? dirty_59_0 : _GEN_1586; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1982 = _cached_stall_T_1 ? dirty_59_1 : _GEN_1587; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1983 = _cached_stall_T_1 ? dirty_60_0 : _GEN_1588; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1984 = _cached_stall_T_1 ? dirty_60_1 : _GEN_1589; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1985 = _cached_stall_T_1 ? dirty_61_0 : _GEN_1590; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1986 = _cached_stall_T_1 ? dirty_61_1 : _GEN_1591; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1987 = _cached_stall_T_1 ? dirty_62_0 : _GEN_1592; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1988 = _cached_stall_T_1 ? dirty_62_1 : _GEN_1593; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1989 = _cached_stall_T_1 ? dirty_63_0 : _GEN_1594; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1990 = _cached_stall_T_1 ? dirty_63_1 : _GEN_1595; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1991 = _cached_stall_T_1 ? dirty_64_0 : _GEN_1596; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1992 = _cached_stall_T_1 ? dirty_64_1 : _GEN_1597; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1993 = _cached_stall_T_1 ? dirty_65_0 : _GEN_1598; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1994 = _cached_stall_T_1 ? dirty_65_1 : _GEN_1599; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1995 = _cached_stall_T_1 ? dirty_66_0 : _GEN_1600; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1996 = _cached_stall_T_1 ? dirty_66_1 : _GEN_1601; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1997 = _cached_stall_T_1 ? dirty_67_0 : _GEN_1602; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1998 = _cached_stall_T_1 ? dirty_67_1 : _GEN_1603; // @[DCache.scala 298:28 69:22]
  wire  _GEN_1999 = _cached_stall_T_1 ? dirty_68_0 : _GEN_1604; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2000 = _cached_stall_T_1 ? dirty_68_1 : _GEN_1605; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2001 = _cached_stall_T_1 ? dirty_69_0 : _GEN_1606; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2002 = _cached_stall_T_1 ? dirty_69_1 : _GEN_1607; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2003 = _cached_stall_T_1 ? dirty_70_0 : _GEN_1608; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2004 = _cached_stall_T_1 ? dirty_70_1 : _GEN_1609; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2005 = _cached_stall_T_1 ? dirty_71_0 : _GEN_1610; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2006 = _cached_stall_T_1 ? dirty_71_1 : _GEN_1611; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2007 = _cached_stall_T_1 ? dirty_72_0 : _GEN_1612; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2008 = _cached_stall_T_1 ? dirty_72_1 : _GEN_1613; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2009 = _cached_stall_T_1 ? dirty_73_0 : _GEN_1614; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2010 = _cached_stall_T_1 ? dirty_73_1 : _GEN_1615; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2011 = _cached_stall_T_1 ? dirty_74_0 : _GEN_1616; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2012 = _cached_stall_T_1 ? dirty_74_1 : _GEN_1617; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2013 = _cached_stall_T_1 ? dirty_75_0 : _GEN_1618; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2014 = _cached_stall_T_1 ? dirty_75_1 : _GEN_1619; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2015 = _cached_stall_T_1 ? dirty_76_0 : _GEN_1620; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2016 = _cached_stall_T_1 ? dirty_76_1 : _GEN_1621; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2017 = _cached_stall_T_1 ? dirty_77_0 : _GEN_1622; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2018 = _cached_stall_T_1 ? dirty_77_1 : _GEN_1623; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2019 = _cached_stall_T_1 ? dirty_78_0 : _GEN_1624; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2020 = _cached_stall_T_1 ? dirty_78_1 : _GEN_1625; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2021 = _cached_stall_T_1 ? dirty_79_0 : _GEN_1626; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2022 = _cached_stall_T_1 ? dirty_79_1 : _GEN_1627; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2023 = _cached_stall_T_1 ? dirty_80_0 : _GEN_1628; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2024 = _cached_stall_T_1 ? dirty_80_1 : _GEN_1629; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2025 = _cached_stall_T_1 ? dirty_81_0 : _GEN_1630; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2026 = _cached_stall_T_1 ? dirty_81_1 : _GEN_1631; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2027 = _cached_stall_T_1 ? dirty_82_0 : _GEN_1632; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2028 = _cached_stall_T_1 ? dirty_82_1 : _GEN_1633; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2029 = _cached_stall_T_1 ? dirty_83_0 : _GEN_1634; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2030 = _cached_stall_T_1 ? dirty_83_1 : _GEN_1635; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2031 = _cached_stall_T_1 ? dirty_84_0 : _GEN_1636; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2032 = _cached_stall_T_1 ? dirty_84_1 : _GEN_1637; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2033 = _cached_stall_T_1 ? dirty_85_0 : _GEN_1638; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2034 = _cached_stall_T_1 ? dirty_85_1 : _GEN_1639; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2035 = _cached_stall_T_1 ? dirty_86_0 : _GEN_1640; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2036 = _cached_stall_T_1 ? dirty_86_1 : _GEN_1641; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2037 = _cached_stall_T_1 ? dirty_87_0 : _GEN_1642; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2038 = _cached_stall_T_1 ? dirty_87_1 : _GEN_1643; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2039 = _cached_stall_T_1 ? dirty_88_0 : _GEN_1644; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2040 = _cached_stall_T_1 ? dirty_88_1 : _GEN_1645; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2041 = _cached_stall_T_1 ? dirty_89_0 : _GEN_1646; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2042 = _cached_stall_T_1 ? dirty_89_1 : _GEN_1647; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2043 = _cached_stall_T_1 ? dirty_90_0 : _GEN_1648; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2044 = _cached_stall_T_1 ? dirty_90_1 : _GEN_1649; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2045 = _cached_stall_T_1 ? dirty_91_0 : _GEN_1650; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2046 = _cached_stall_T_1 ? dirty_91_1 : _GEN_1651; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2047 = _cached_stall_T_1 ? dirty_92_0 : _GEN_1652; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2048 = _cached_stall_T_1 ? dirty_92_1 : _GEN_1653; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2049 = _cached_stall_T_1 ? dirty_93_0 : _GEN_1654; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2050 = _cached_stall_T_1 ? dirty_93_1 : _GEN_1655; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2051 = _cached_stall_T_1 ? dirty_94_0 : _GEN_1656; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2052 = _cached_stall_T_1 ? dirty_94_1 : _GEN_1657; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2053 = _cached_stall_T_1 ? dirty_95_0 : _GEN_1658; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2054 = _cached_stall_T_1 ? dirty_95_1 : _GEN_1659; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2055 = _cached_stall_T_1 ? dirty_96_0 : _GEN_1660; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2056 = _cached_stall_T_1 ? dirty_96_1 : _GEN_1661; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2057 = _cached_stall_T_1 ? dirty_97_0 : _GEN_1662; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2058 = _cached_stall_T_1 ? dirty_97_1 : _GEN_1663; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2059 = _cached_stall_T_1 ? dirty_98_0 : _GEN_1664; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2060 = _cached_stall_T_1 ? dirty_98_1 : _GEN_1665; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2061 = _cached_stall_T_1 ? dirty_99_0 : _GEN_1666; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2062 = _cached_stall_T_1 ? dirty_99_1 : _GEN_1667; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2063 = _cached_stall_T_1 ? dirty_100_0 : _GEN_1668; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2064 = _cached_stall_T_1 ? dirty_100_1 : _GEN_1669; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2065 = _cached_stall_T_1 ? dirty_101_0 : _GEN_1670; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2066 = _cached_stall_T_1 ? dirty_101_1 : _GEN_1671; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2067 = _cached_stall_T_1 ? dirty_102_0 : _GEN_1672; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2068 = _cached_stall_T_1 ? dirty_102_1 : _GEN_1673; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2069 = _cached_stall_T_1 ? dirty_103_0 : _GEN_1674; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2070 = _cached_stall_T_1 ? dirty_103_1 : _GEN_1675; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2071 = _cached_stall_T_1 ? dirty_104_0 : _GEN_1676; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2072 = _cached_stall_T_1 ? dirty_104_1 : _GEN_1677; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2073 = _cached_stall_T_1 ? dirty_105_0 : _GEN_1678; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2074 = _cached_stall_T_1 ? dirty_105_1 : _GEN_1679; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2075 = _cached_stall_T_1 ? dirty_106_0 : _GEN_1680; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2076 = _cached_stall_T_1 ? dirty_106_1 : _GEN_1681; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2077 = _cached_stall_T_1 ? dirty_107_0 : _GEN_1682; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2078 = _cached_stall_T_1 ? dirty_107_1 : _GEN_1683; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2079 = _cached_stall_T_1 ? dirty_108_0 : _GEN_1684; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2080 = _cached_stall_T_1 ? dirty_108_1 : _GEN_1685; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2081 = _cached_stall_T_1 ? dirty_109_0 : _GEN_1686; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2082 = _cached_stall_T_1 ? dirty_109_1 : _GEN_1687; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2083 = _cached_stall_T_1 ? dirty_110_0 : _GEN_1688; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2084 = _cached_stall_T_1 ? dirty_110_1 : _GEN_1689; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2085 = _cached_stall_T_1 ? dirty_111_0 : _GEN_1690; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2086 = _cached_stall_T_1 ? dirty_111_1 : _GEN_1691; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2087 = _cached_stall_T_1 ? dirty_112_0 : _GEN_1692; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2088 = _cached_stall_T_1 ? dirty_112_1 : _GEN_1693; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2089 = _cached_stall_T_1 ? dirty_113_0 : _GEN_1694; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2090 = _cached_stall_T_1 ? dirty_113_1 : _GEN_1695; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2091 = _cached_stall_T_1 ? dirty_114_0 : _GEN_1696; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2092 = _cached_stall_T_1 ? dirty_114_1 : _GEN_1697; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2093 = _cached_stall_T_1 ? dirty_115_0 : _GEN_1698; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2094 = _cached_stall_T_1 ? dirty_115_1 : _GEN_1699; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2095 = _cached_stall_T_1 ? dirty_116_0 : _GEN_1700; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2096 = _cached_stall_T_1 ? dirty_116_1 : _GEN_1701; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2097 = _cached_stall_T_1 ? dirty_117_0 : _GEN_1702; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2098 = _cached_stall_T_1 ? dirty_117_1 : _GEN_1703; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2099 = _cached_stall_T_1 ? dirty_118_0 : _GEN_1704; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2100 = _cached_stall_T_1 ? dirty_118_1 : _GEN_1705; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2101 = _cached_stall_T_1 ? dirty_119_0 : _GEN_1706; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2102 = _cached_stall_T_1 ? dirty_119_1 : _GEN_1707; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2103 = _cached_stall_T_1 ? dirty_120_0 : _GEN_1708; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2104 = _cached_stall_T_1 ? dirty_120_1 : _GEN_1709; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2105 = _cached_stall_T_1 ? dirty_121_0 : _GEN_1710; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2106 = _cached_stall_T_1 ? dirty_121_1 : _GEN_1711; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2107 = _cached_stall_T_1 ? dirty_122_0 : _GEN_1712; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2108 = _cached_stall_T_1 ? dirty_122_1 : _GEN_1713; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2109 = _cached_stall_T_1 ? dirty_123_0 : _GEN_1714; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2110 = _cached_stall_T_1 ? dirty_123_1 : _GEN_1715; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2111 = _cached_stall_T_1 ? dirty_124_0 : _GEN_1716; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2112 = _cached_stall_T_1 ? dirty_124_1 : _GEN_1717; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2113 = _cached_stall_T_1 ? dirty_125_0 : _GEN_1718; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2114 = _cached_stall_T_1 ? dirty_125_1 : _GEN_1719; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2115 = _cached_stall_T_1 ? dirty_126_0 : _GEN_1720; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2116 = _cached_stall_T_1 ? dirty_126_1 : _GEN_1721; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2117 = _cached_stall_T_1 ? dirty_127_0 : _GEN_1722; // @[DCache.scala 298:28 69:22]
  wire  _GEN_2118 = _cached_stall_T_1 ? dirty_127_1 : _GEN_1723; // @[DCache.scala 298:28 69:22]
  wire [31:0] _GEN_2119 = _cached_stall_T_1 ? saved_rdata : _GEN_1724; // @[DCache.scala 141:28 298:28]
  wire  _GEN_2120 = M_mem_uncached & _GEN_302; // @[DCache.scala 271:36 83:29]
  wire [31:0] _GEN_2121 = M_mem_uncached ? _GEN_303 : 32'h0; // @[DCache.scala 271:36 84:29]
  wire [1:0] _GEN_2122 = M_mem_uncached ? _GEN_304 : 2'h0; // @[DCache.scala 271:36 84:29]
  wire [3:0] _GEN_2123 = M_mem_uncached ? _GEN_305 : 4'h0; // @[DCache.scala 271:36 84:29]
  wire [31:0] _GEN_2124 = M_mem_uncached ? _GEN_306 : 32'h0; // @[DCache.scala 271:36 84:29]
  wire  _GEN_2125 = M_mem_uncached ? _GEN_307 : current_mmio_write_saved; // @[DCache.scala 271:36 216:41]
  wire [31:0] _GEN_2126 = M_mem_uncached ? _GEN_308 : ar_addr; // @[DCache.scala 199:24 271:36]
  wire [7:0] _GEN_2127 = M_mem_uncached ? _GEN_309 : ar_len; // @[DCache.scala 199:24 271:36]
  wire [2:0] _GEN_2128 = M_mem_uncached ? _GEN_310 : ar_size; // @[DCache.scala 199:24 271:36]
  wire  _GEN_2129 = M_mem_uncached ? _GEN_311 : arvalid; // @[DCache.scala 200:24 271:36]
  wire [2:0] _GEN_2130 = M_mem_uncached ? _GEN_312 : _GEN_1726; // @[DCache.scala 271:36]
  wire  _GEN_2131 = M_mem_uncached ? _GEN_313 : rready; // @[DCache.scala 203:23 271:36]
  wire [3:0] _GEN_2132 = M_mem_uncached ? axi_wcnt : _GEN_1727; // @[DCache.scala 271:36 89:40]
  wire [9:0] _GEN_2133 = M_mem_uncached ? bram_replace_addr : _GEN_1728; // @[DCache.scala 271:36 90:40]
  wire [9:0] _GEN_2134 = M_mem_uncached ? bram_read_ready_addr : _GEN_1729; // @[DCache.scala 271:36 91:40]
  wire [9:0] _GEN_2135 = M_mem_uncached ? bram_replace_write_addr : _GEN_1730; // @[DCache.scala 271:36 92:40]
  wire  _GEN_2137 = M_mem_uncached ? bram_use_replace_addr : _GEN_1732; // @[DCache.scala 271:36 95:40]
  wire  _GEN_2139 = M_mem_uncached ? replace_writeback : _GEN_1734; // @[DCache.scala 271:36 101:40]
  wire  _GEN_2140 = M_mem_uncached ? lru_0 : _GEN_1735; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2141 = M_mem_uncached ? lru_1 : _GEN_1736; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2142 = M_mem_uncached ? lru_2 : _GEN_1737; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2143 = M_mem_uncached ? lru_3 : _GEN_1738; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2144 = M_mem_uncached ? lru_4 : _GEN_1739; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2145 = M_mem_uncached ? lru_5 : _GEN_1740; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2146 = M_mem_uncached ? lru_6 : _GEN_1741; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2147 = M_mem_uncached ? lru_7 : _GEN_1742; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2148 = M_mem_uncached ? lru_8 : _GEN_1743; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2149 = M_mem_uncached ? lru_9 : _GEN_1744; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2150 = M_mem_uncached ? lru_10 : _GEN_1745; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2151 = M_mem_uncached ? lru_11 : _GEN_1746; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2152 = M_mem_uncached ? lru_12 : _GEN_1747; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2153 = M_mem_uncached ? lru_13 : _GEN_1748; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2154 = M_mem_uncached ? lru_14 : _GEN_1749; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2155 = M_mem_uncached ? lru_15 : _GEN_1750; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2156 = M_mem_uncached ? lru_16 : _GEN_1751; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2157 = M_mem_uncached ? lru_17 : _GEN_1752; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2158 = M_mem_uncached ? lru_18 : _GEN_1753; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2159 = M_mem_uncached ? lru_19 : _GEN_1754; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2160 = M_mem_uncached ? lru_20 : _GEN_1755; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2161 = M_mem_uncached ? lru_21 : _GEN_1756; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2162 = M_mem_uncached ? lru_22 : _GEN_1757; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2163 = M_mem_uncached ? lru_23 : _GEN_1758; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2164 = M_mem_uncached ? lru_24 : _GEN_1759; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2165 = M_mem_uncached ? lru_25 : _GEN_1760; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2166 = M_mem_uncached ? lru_26 : _GEN_1761; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2167 = M_mem_uncached ? lru_27 : _GEN_1762; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2168 = M_mem_uncached ? lru_28 : _GEN_1763; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2169 = M_mem_uncached ? lru_29 : _GEN_1764; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2170 = M_mem_uncached ? lru_30 : _GEN_1765; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2171 = M_mem_uncached ? lru_31 : _GEN_1766; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2172 = M_mem_uncached ? lru_32 : _GEN_1767; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2173 = M_mem_uncached ? lru_33 : _GEN_1768; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2174 = M_mem_uncached ? lru_34 : _GEN_1769; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2175 = M_mem_uncached ? lru_35 : _GEN_1770; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2176 = M_mem_uncached ? lru_36 : _GEN_1771; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2177 = M_mem_uncached ? lru_37 : _GEN_1772; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2178 = M_mem_uncached ? lru_38 : _GEN_1773; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2179 = M_mem_uncached ? lru_39 : _GEN_1774; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2180 = M_mem_uncached ? lru_40 : _GEN_1775; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2181 = M_mem_uncached ? lru_41 : _GEN_1776; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2182 = M_mem_uncached ? lru_42 : _GEN_1777; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2183 = M_mem_uncached ? lru_43 : _GEN_1778; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2184 = M_mem_uncached ? lru_44 : _GEN_1779; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2185 = M_mem_uncached ? lru_45 : _GEN_1780; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2186 = M_mem_uncached ? lru_46 : _GEN_1781; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2187 = M_mem_uncached ? lru_47 : _GEN_1782; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2188 = M_mem_uncached ? lru_48 : _GEN_1783; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2189 = M_mem_uncached ? lru_49 : _GEN_1784; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2190 = M_mem_uncached ? lru_50 : _GEN_1785; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2191 = M_mem_uncached ? lru_51 : _GEN_1786; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2192 = M_mem_uncached ? lru_52 : _GEN_1787; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2193 = M_mem_uncached ? lru_53 : _GEN_1788; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2194 = M_mem_uncached ? lru_54 : _GEN_1789; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2195 = M_mem_uncached ? lru_55 : _GEN_1790; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2196 = M_mem_uncached ? lru_56 : _GEN_1791; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2197 = M_mem_uncached ? lru_57 : _GEN_1792; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2198 = M_mem_uncached ? lru_58 : _GEN_1793; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2199 = M_mem_uncached ? lru_59 : _GEN_1794; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2200 = M_mem_uncached ? lru_60 : _GEN_1795; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2201 = M_mem_uncached ? lru_61 : _GEN_1796; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2202 = M_mem_uncached ? lru_62 : _GEN_1797; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2203 = M_mem_uncached ? lru_63 : _GEN_1798; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2204 = M_mem_uncached ? lru_64 : _GEN_1799; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2205 = M_mem_uncached ? lru_65 : _GEN_1800; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2206 = M_mem_uncached ? lru_66 : _GEN_1801; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2207 = M_mem_uncached ? lru_67 : _GEN_1802; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2208 = M_mem_uncached ? lru_68 : _GEN_1803; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2209 = M_mem_uncached ? lru_69 : _GEN_1804; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2210 = M_mem_uncached ? lru_70 : _GEN_1805; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2211 = M_mem_uncached ? lru_71 : _GEN_1806; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2212 = M_mem_uncached ? lru_72 : _GEN_1807; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2213 = M_mem_uncached ? lru_73 : _GEN_1808; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2214 = M_mem_uncached ? lru_74 : _GEN_1809; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2215 = M_mem_uncached ? lru_75 : _GEN_1810; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2216 = M_mem_uncached ? lru_76 : _GEN_1811; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2217 = M_mem_uncached ? lru_77 : _GEN_1812; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2218 = M_mem_uncached ? lru_78 : _GEN_1813; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2219 = M_mem_uncached ? lru_79 : _GEN_1814; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2220 = M_mem_uncached ? lru_80 : _GEN_1815; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2221 = M_mem_uncached ? lru_81 : _GEN_1816; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2222 = M_mem_uncached ? lru_82 : _GEN_1817; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2223 = M_mem_uncached ? lru_83 : _GEN_1818; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2224 = M_mem_uncached ? lru_84 : _GEN_1819; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2225 = M_mem_uncached ? lru_85 : _GEN_1820; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2226 = M_mem_uncached ? lru_86 : _GEN_1821; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2227 = M_mem_uncached ? lru_87 : _GEN_1822; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2228 = M_mem_uncached ? lru_88 : _GEN_1823; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2229 = M_mem_uncached ? lru_89 : _GEN_1824; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2230 = M_mem_uncached ? lru_90 : _GEN_1825; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2231 = M_mem_uncached ? lru_91 : _GEN_1826; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2232 = M_mem_uncached ? lru_92 : _GEN_1827; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2233 = M_mem_uncached ? lru_93 : _GEN_1828; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2234 = M_mem_uncached ? lru_94 : _GEN_1829; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2235 = M_mem_uncached ? lru_95 : _GEN_1830; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2236 = M_mem_uncached ? lru_96 : _GEN_1831; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2237 = M_mem_uncached ? lru_97 : _GEN_1832; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2238 = M_mem_uncached ? lru_98 : _GEN_1833; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2239 = M_mem_uncached ? lru_99 : _GEN_1834; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2240 = M_mem_uncached ? lru_100 : _GEN_1835; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2241 = M_mem_uncached ? lru_101 : _GEN_1836; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2242 = M_mem_uncached ? lru_102 : _GEN_1837; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2243 = M_mem_uncached ? lru_103 : _GEN_1838; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2244 = M_mem_uncached ? lru_104 : _GEN_1839; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2245 = M_mem_uncached ? lru_105 : _GEN_1840; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2246 = M_mem_uncached ? lru_106 : _GEN_1841; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2247 = M_mem_uncached ? lru_107 : _GEN_1842; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2248 = M_mem_uncached ? lru_108 : _GEN_1843; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2249 = M_mem_uncached ? lru_109 : _GEN_1844; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2250 = M_mem_uncached ? lru_110 : _GEN_1845; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2251 = M_mem_uncached ? lru_111 : _GEN_1846; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2252 = M_mem_uncached ? lru_112 : _GEN_1847; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2253 = M_mem_uncached ? lru_113 : _GEN_1848; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2254 = M_mem_uncached ? lru_114 : _GEN_1849; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2255 = M_mem_uncached ? lru_115 : _GEN_1850; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2256 = M_mem_uncached ? lru_116 : _GEN_1851; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2257 = M_mem_uncached ? lru_117 : _GEN_1852; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2258 = M_mem_uncached ? lru_118 : _GEN_1853; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2259 = M_mem_uncached ? lru_119 : _GEN_1854; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2260 = M_mem_uncached ? lru_120 : _GEN_1855; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2261 = M_mem_uncached ? lru_121 : _GEN_1856; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2262 = M_mem_uncached ? lru_122 : _GEN_1857; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2263 = M_mem_uncached ? lru_123 : _GEN_1858; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2264 = M_mem_uncached ? lru_124 : _GEN_1859; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2265 = M_mem_uncached ? lru_125 : _GEN_1860; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2266 = M_mem_uncached ? lru_126 : _GEN_1861; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2267 = M_mem_uncached ? lru_127 : _GEN_1862; // @[DCache.scala 271:36 70:22]
  wire  _GEN_2268 = M_mem_uncached ? dirty_0_0 : _GEN_1863; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2269 = M_mem_uncached ? dirty_0_1 : _GEN_1864; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2270 = M_mem_uncached ? dirty_1_0 : _GEN_1865; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2271 = M_mem_uncached ? dirty_1_1 : _GEN_1866; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2272 = M_mem_uncached ? dirty_2_0 : _GEN_1867; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2273 = M_mem_uncached ? dirty_2_1 : _GEN_1868; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2274 = M_mem_uncached ? dirty_3_0 : _GEN_1869; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2275 = M_mem_uncached ? dirty_3_1 : _GEN_1870; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2276 = M_mem_uncached ? dirty_4_0 : _GEN_1871; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2277 = M_mem_uncached ? dirty_4_1 : _GEN_1872; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2278 = M_mem_uncached ? dirty_5_0 : _GEN_1873; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2279 = M_mem_uncached ? dirty_5_1 : _GEN_1874; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2280 = M_mem_uncached ? dirty_6_0 : _GEN_1875; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2281 = M_mem_uncached ? dirty_6_1 : _GEN_1876; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2282 = M_mem_uncached ? dirty_7_0 : _GEN_1877; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2283 = M_mem_uncached ? dirty_7_1 : _GEN_1878; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2284 = M_mem_uncached ? dirty_8_0 : _GEN_1879; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2285 = M_mem_uncached ? dirty_8_1 : _GEN_1880; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2286 = M_mem_uncached ? dirty_9_0 : _GEN_1881; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2287 = M_mem_uncached ? dirty_9_1 : _GEN_1882; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2288 = M_mem_uncached ? dirty_10_0 : _GEN_1883; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2289 = M_mem_uncached ? dirty_10_1 : _GEN_1884; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2290 = M_mem_uncached ? dirty_11_0 : _GEN_1885; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2291 = M_mem_uncached ? dirty_11_1 : _GEN_1886; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2292 = M_mem_uncached ? dirty_12_0 : _GEN_1887; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2293 = M_mem_uncached ? dirty_12_1 : _GEN_1888; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2294 = M_mem_uncached ? dirty_13_0 : _GEN_1889; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2295 = M_mem_uncached ? dirty_13_1 : _GEN_1890; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2296 = M_mem_uncached ? dirty_14_0 : _GEN_1891; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2297 = M_mem_uncached ? dirty_14_1 : _GEN_1892; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2298 = M_mem_uncached ? dirty_15_0 : _GEN_1893; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2299 = M_mem_uncached ? dirty_15_1 : _GEN_1894; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2300 = M_mem_uncached ? dirty_16_0 : _GEN_1895; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2301 = M_mem_uncached ? dirty_16_1 : _GEN_1896; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2302 = M_mem_uncached ? dirty_17_0 : _GEN_1897; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2303 = M_mem_uncached ? dirty_17_1 : _GEN_1898; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2304 = M_mem_uncached ? dirty_18_0 : _GEN_1899; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2305 = M_mem_uncached ? dirty_18_1 : _GEN_1900; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2306 = M_mem_uncached ? dirty_19_0 : _GEN_1901; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2307 = M_mem_uncached ? dirty_19_1 : _GEN_1902; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2308 = M_mem_uncached ? dirty_20_0 : _GEN_1903; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2309 = M_mem_uncached ? dirty_20_1 : _GEN_1904; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2310 = M_mem_uncached ? dirty_21_0 : _GEN_1905; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2311 = M_mem_uncached ? dirty_21_1 : _GEN_1906; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2312 = M_mem_uncached ? dirty_22_0 : _GEN_1907; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2313 = M_mem_uncached ? dirty_22_1 : _GEN_1908; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2314 = M_mem_uncached ? dirty_23_0 : _GEN_1909; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2315 = M_mem_uncached ? dirty_23_1 : _GEN_1910; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2316 = M_mem_uncached ? dirty_24_0 : _GEN_1911; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2317 = M_mem_uncached ? dirty_24_1 : _GEN_1912; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2318 = M_mem_uncached ? dirty_25_0 : _GEN_1913; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2319 = M_mem_uncached ? dirty_25_1 : _GEN_1914; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2320 = M_mem_uncached ? dirty_26_0 : _GEN_1915; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2321 = M_mem_uncached ? dirty_26_1 : _GEN_1916; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2322 = M_mem_uncached ? dirty_27_0 : _GEN_1917; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2323 = M_mem_uncached ? dirty_27_1 : _GEN_1918; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2324 = M_mem_uncached ? dirty_28_0 : _GEN_1919; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2325 = M_mem_uncached ? dirty_28_1 : _GEN_1920; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2326 = M_mem_uncached ? dirty_29_0 : _GEN_1921; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2327 = M_mem_uncached ? dirty_29_1 : _GEN_1922; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2328 = M_mem_uncached ? dirty_30_0 : _GEN_1923; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2329 = M_mem_uncached ? dirty_30_1 : _GEN_1924; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2330 = M_mem_uncached ? dirty_31_0 : _GEN_1925; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2331 = M_mem_uncached ? dirty_31_1 : _GEN_1926; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2332 = M_mem_uncached ? dirty_32_0 : _GEN_1927; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2333 = M_mem_uncached ? dirty_32_1 : _GEN_1928; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2334 = M_mem_uncached ? dirty_33_0 : _GEN_1929; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2335 = M_mem_uncached ? dirty_33_1 : _GEN_1930; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2336 = M_mem_uncached ? dirty_34_0 : _GEN_1931; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2337 = M_mem_uncached ? dirty_34_1 : _GEN_1932; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2338 = M_mem_uncached ? dirty_35_0 : _GEN_1933; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2339 = M_mem_uncached ? dirty_35_1 : _GEN_1934; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2340 = M_mem_uncached ? dirty_36_0 : _GEN_1935; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2341 = M_mem_uncached ? dirty_36_1 : _GEN_1936; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2342 = M_mem_uncached ? dirty_37_0 : _GEN_1937; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2343 = M_mem_uncached ? dirty_37_1 : _GEN_1938; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2344 = M_mem_uncached ? dirty_38_0 : _GEN_1939; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2345 = M_mem_uncached ? dirty_38_1 : _GEN_1940; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2346 = M_mem_uncached ? dirty_39_0 : _GEN_1941; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2347 = M_mem_uncached ? dirty_39_1 : _GEN_1942; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2348 = M_mem_uncached ? dirty_40_0 : _GEN_1943; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2349 = M_mem_uncached ? dirty_40_1 : _GEN_1944; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2350 = M_mem_uncached ? dirty_41_0 : _GEN_1945; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2351 = M_mem_uncached ? dirty_41_1 : _GEN_1946; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2352 = M_mem_uncached ? dirty_42_0 : _GEN_1947; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2353 = M_mem_uncached ? dirty_42_1 : _GEN_1948; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2354 = M_mem_uncached ? dirty_43_0 : _GEN_1949; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2355 = M_mem_uncached ? dirty_43_1 : _GEN_1950; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2356 = M_mem_uncached ? dirty_44_0 : _GEN_1951; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2357 = M_mem_uncached ? dirty_44_1 : _GEN_1952; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2358 = M_mem_uncached ? dirty_45_0 : _GEN_1953; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2359 = M_mem_uncached ? dirty_45_1 : _GEN_1954; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2360 = M_mem_uncached ? dirty_46_0 : _GEN_1955; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2361 = M_mem_uncached ? dirty_46_1 : _GEN_1956; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2362 = M_mem_uncached ? dirty_47_0 : _GEN_1957; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2363 = M_mem_uncached ? dirty_47_1 : _GEN_1958; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2364 = M_mem_uncached ? dirty_48_0 : _GEN_1959; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2365 = M_mem_uncached ? dirty_48_1 : _GEN_1960; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2366 = M_mem_uncached ? dirty_49_0 : _GEN_1961; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2367 = M_mem_uncached ? dirty_49_1 : _GEN_1962; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2368 = M_mem_uncached ? dirty_50_0 : _GEN_1963; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2369 = M_mem_uncached ? dirty_50_1 : _GEN_1964; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2370 = M_mem_uncached ? dirty_51_0 : _GEN_1965; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2371 = M_mem_uncached ? dirty_51_1 : _GEN_1966; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2372 = M_mem_uncached ? dirty_52_0 : _GEN_1967; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2373 = M_mem_uncached ? dirty_52_1 : _GEN_1968; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2374 = M_mem_uncached ? dirty_53_0 : _GEN_1969; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2375 = M_mem_uncached ? dirty_53_1 : _GEN_1970; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2376 = M_mem_uncached ? dirty_54_0 : _GEN_1971; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2377 = M_mem_uncached ? dirty_54_1 : _GEN_1972; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2378 = M_mem_uncached ? dirty_55_0 : _GEN_1973; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2379 = M_mem_uncached ? dirty_55_1 : _GEN_1974; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2380 = M_mem_uncached ? dirty_56_0 : _GEN_1975; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2381 = M_mem_uncached ? dirty_56_1 : _GEN_1976; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2382 = M_mem_uncached ? dirty_57_0 : _GEN_1977; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2383 = M_mem_uncached ? dirty_57_1 : _GEN_1978; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2384 = M_mem_uncached ? dirty_58_0 : _GEN_1979; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2385 = M_mem_uncached ? dirty_58_1 : _GEN_1980; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2386 = M_mem_uncached ? dirty_59_0 : _GEN_1981; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2387 = M_mem_uncached ? dirty_59_1 : _GEN_1982; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2388 = M_mem_uncached ? dirty_60_0 : _GEN_1983; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2389 = M_mem_uncached ? dirty_60_1 : _GEN_1984; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2390 = M_mem_uncached ? dirty_61_0 : _GEN_1985; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2391 = M_mem_uncached ? dirty_61_1 : _GEN_1986; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2392 = M_mem_uncached ? dirty_62_0 : _GEN_1987; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2393 = M_mem_uncached ? dirty_62_1 : _GEN_1988; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2394 = M_mem_uncached ? dirty_63_0 : _GEN_1989; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2395 = M_mem_uncached ? dirty_63_1 : _GEN_1990; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2396 = M_mem_uncached ? dirty_64_0 : _GEN_1991; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2397 = M_mem_uncached ? dirty_64_1 : _GEN_1992; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2398 = M_mem_uncached ? dirty_65_0 : _GEN_1993; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2399 = M_mem_uncached ? dirty_65_1 : _GEN_1994; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2400 = M_mem_uncached ? dirty_66_0 : _GEN_1995; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2401 = M_mem_uncached ? dirty_66_1 : _GEN_1996; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2402 = M_mem_uncached ? dirty_67_0 : _GEN_1997; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2403 = M_mem_uncached ? dirty_67_1 : _GEN_1998; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2404 = M_mem_uncached ? dirty_68_0 : _GEN_1999; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2405 = M_mem_uncached ? dirty_68_1 : _GEN_2000; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2406 = M_mem_uncached ? dirty_69_0 : _GEN_2001; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2407 = M_mem_uncached ? dirty_69_1 : _GEN_2002; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2408 = M_mem_uncached ? dirty_70_0 : _GEN_2003; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2409 = M_mem_uncached ? dirty_70_1 : _GEN_2004; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2410 = M_mem_uncached ? dirty_71_0 : _GEN_2005; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2411 = M_mem_uncached ? dirty_71_1 : _GEN_2006; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2412 = M_mem_uncached ? dirty_72_0 : _GEN_2007; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2413 = M_mem_uncached ? dirty_72_1 : _GEN_2008; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2414 = M_mem_uncached ? dirty_73_0 : _GEN_2009; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2415 = M_mem_uncached ? dirty_73_1 : _GEN_2010; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2416 = M_mem_uncached ? dirty_74_0 : _GEN_2011; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2417 = M_mem_uncached ? dirty_74_1 : _GEN_2012; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2418 = M_mem_uncached ? dirty_75_0 : _GEN_2013; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2419 = M_mem_uncached ? dirty_75_1 : _GEN_2014; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2420 = M_mem_uncached ? dirty_76_0 : _GEN_2015; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2421 = M_mem_uncached ? dirty_76_1 : _GEN_2016; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2422 = M_mem_uncached ? dirty_77_0 : _GEN_2017; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2423 = M_mem_uncached ? dirty_77_1 : _GEN_2018; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2424 = M_mem_uncached ? dirty_78_0 : _GEN_2019; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2425 = M_mem_uncached ? dirty_78_1 : _GEN_2020; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2426 = M_mem_uncached ? dirty_79_0 : _GEN_2021; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2427 = M_mem_uncached ? dirty_79_1 : _GEN_2022; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2428 = M_mem_uncached ? dirty_80_0 : _GEN_2023; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2429 = M_mem_uncached ? dirty_80_1 : _GEN_2024; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2430 = M_mem_uncached ? dirty_81_0 : _GEN_2025; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2431 = M_mem_uncached ? dirty_81_1 : _GEN_2026; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2432 = M_mem_uncached ? dirty_82_0 : _GEN_2027; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2433 = M_mem_uncached ? dirty_82_1 : _GEN_2028; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2434 = M_mem_uncached ? dirty_83_0 : _GEN_2029; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2435 = M_mem_uncached ? dirty_83_1 : _GEN_2030; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2436 = M_mem_uncached ? dirty_84_0 : _GEN_2031; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2437 = M_mem_uncached ? dirty_84_1 : _GEN_2032; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2438 = M_mem_uncached ? dirty_85_0 : _GEN_2033; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2439 = M_mem_uncached ? dirty_85_1 : _GEN_2034; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2440 = M_mem_uncached ? dirty_86_0 : _GEN_2035; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2441 = M_mem_uncached ? dirty_86_1 : _GEN_2036; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2442 = M_mem_uncached ? dirty_87_0 : _GEN_2037; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2443 = M_mem_uncached ? dirty_87_1 : _GEN_2038; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2444 = M_mem_uncached ? dirty_88_0 : _GEN_2039; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2445 = M_mem_uncached ? dirty_88_1 : _GEN_2040; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2446 = M_mem_uncached ? dirty_89_0 : _GEN_2041; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2447 = M_mem_uncached ? dirty_89_1 : _GEN_2042; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2448 = M_mem_uncached ? dirty_90_0 : _GEN_2043; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2449 = M_mem_uncached ? dirty_90_1 : _GEN_2044; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2450 = M_mem_uncached ? dirty_91_0 : _GEN_2045; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2451 = M_mem_uncached ? dirty_91_1 : _GEN_2046; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2452 = M_mem_uncached ? dirty_92_0 : _GEN_2047; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2453 = M_mem_uncached ? dirty_92_1 : _GEN_2048; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2454 = M_mem_uncached ? dirty_93_0 : _GEN_2049; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2455 = M_mem_uncached ? dirty_93_1 : _GEN_2050; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2456 = M_mem_uncached ? dirty_94_0 : _GEN_2051; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2457 = M_mem_uncached ? dirty_94_1 : _GEN_2052; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2458 = M_mem_uncached ? dirty_95_0 : _GEN_2053; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2459 = M_mem_uncached ? dirty_95_1 : _GEN_2054; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2460 = M_mem_uncached ? dirty_96_0 : _GEN_2055; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2461 = M_mem_uncached ? dirty_96_1 : _GEN_2056; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2462 = M_mem_uncached ? dirty_97_0 : _GEN_2057; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2463 = M_mem_uncached ? dirty_97_1 : _GEN_2058; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2464 = M_mem_uncached ? dirty_98_0 : _GEN_2059; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2465 = M_mem_uncached ? dirty_98_1 : _GEN_2060; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2466 = M_mem_uncached ? dirty_99_0 : _GEN_2061; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2467 = M_mem_uncached ? dirty_99_1 : _GEN_2062; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2468 = M_mem_uncached ? dirty_100_0 : _GEN_2063; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2469 = M_mem_uncached ? dirty_100_1 : _GEN_2064; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2470 = M_mem_uncached ? dirty_101_0 : _GEN_2065; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2471 = M_mem_uncached ? dirty_101_1 : _GEN_2066; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2472 = M_mem_uncached ? dirty_102_0 : _GEN_2067; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2473 = M_mem_uncached ? dirty_102_1 : _GEN_2068; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2474 = M_mem_uncached ? dirty_103_0 : _GEN_2069; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2475 = M_mem_uncached ? dirty_103_1 : _GEN_2070; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2476 = M_mem_uncached ? dirty_104_0 : _GEN_2071; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2477 = M_mem_uncached ? dirty_104_1 : _GEN_2072; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2478 = M_mem_uncached ? dirty_105_0 : _GEN_2073; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2479 = M_mem_uncached ? dirty_105_1 : _GEN_2074; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2480 = M_mem_uncached ? dirty_106_0 : _GEN_2075; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2481 = M_mem_uncached ? dirty_106_1 : _GEN_2076; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2482 = M_mem_uncached ? dirty_107_0 : _GEN_2077; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2483 = M_mem_uncached ? dirty_107_1 : _GEN_2078; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2484 = M_mem_uncached ? dirty_108_0 : _GEN_2079; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2485 = M_mem_uncached ? dirty_108_1 : _GEN_2080; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2486 = M_mem_uncached ? dirty_109_0 : _GEN_2081; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2487 = M_mem_uncached ? dirty_109_1 : _GEN_2082; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2488 = M_mem_uncached ? dirty_110_0 : _GEN_2083; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2489 = M_mem_uncached ? dirty_110_1 : _GEN_2084; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2490 = M_mem_uncached ? dirty_111_0 : _GEN_2085; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2491 = M_mem_uncached ? dirty_111_1 : _GEN_2086; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2492 = M_mem_uncached ? dirty_112_0 : _GEN_2087; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2493 = M_mem_uncached ? dirty_112_1 : _GEN_2088; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2494 = M_mem_uncached ? dirty_113_0 : _GEN_2089; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2495 = M_mem_uncached ? dirty_113_1 : _GEN_2090; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2496 = M_mem_uncached ? dirty_114_0 : _GEN_2091; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2497 = M_mem_uncached ? dirty_114_1 : _GEN_2092; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2498 = M_mem_uncached ? dirty_115_0 : _GEN_2093; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2499 = M_mem_uncached ? dirty_115_1 : _GEN_2094; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2500 = M_mem_uncached ? dirty_116_0 : _GEN_2095; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2501 = M_mem_uncached ? dirty_116_1 : _GEN_2096; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2502 = M_mem_uncached ? dirty_117_0 : _GEN_2097; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2503 = M_mem_uncached ? dirty_117_1 : _GEN_2098; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2504 = M_mem_uncached ? dirty_118_0 : _GEN_2099; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2505 = M_mem_uncached ? dirty_118_1 : _GEN_2100; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2506 = M_mem_uncached ? dirty_119_0 : _GEN_2101; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2507 = M_mem_uncached ? dirty_119_1 : _GEN_2102; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2508 = M_mem_uncached ? dirty_120_0 : _GEN_2103; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2509 = M_mem_uncached ? dirty_120_1 : _GEN_2104; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2510 = M_mem_uncached ? dirty_121_0 : _GEN_2105; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2511 = M_mem_uncached ? dirty_121_1 : _GEN_2106; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2512 = M_mem_uncached ? dirty_122_0 : _GEN_2107; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2513 = M_mem_uncached ? dirty_122_1 : _GEN_2108; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2514 = M_mem_uncached ? dirty_123_0 : _GEN_2109; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2515 = M_mem_uncached ? dirty_123_1 : _GEN_2110; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2516 = M_mem_uncached ? dirty_124_0 : _GEN_2111; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2517 = M_mem_uncached ? dirty_124_1 : _GEN_2112; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2518 = M_mem_uncached ? dirty_125_0 : _GEN_2113; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2519 = M_mem_uncached ? dirty_125_1 : _GEN_2114; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2520 = M_mem_uncached ? dirty_126_0 : _GEN_2115; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2521 = M_mem_uncached ? dirty_126_1 : _GEN_2116; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2522 = M_mem_uncached ? dirty_127_0 : _GEN_2117; // @[DCache.scala 271:36 69:22]
  wire  _GEN_2523 = M_mem_uncached ? dirty_127_1 : _GEN_2118; // @[DCache.scala 271:36 69:22]
  wire [31:0] _GEN_2524 = M_mem_uncached ? saved_rdata : _GEN_2119; // @[DCache.scala 141:28 271:36]
  wire [19:0] _GEN_2527 = tlb_stall ? _GEN_288 : {{1'd0}, tlb2_vpn}; // @[DCache.scala 245:21 263:31]
  wire  _GEN_2528 = tlb_stall ? 1'h0 : _GEN_2120; // @[DCache.scala 263:31 83:29]
  wire [31:0] _GEN_2529 = tlb_stall ? 32'h0 : _GEN_2121; // @[DCache.scala 263:31 84:29]
  wire [1:0] _GEN_2530 = tlb_stall ? 2'h0 : _GEN_2122; // @[DCache.scala 263:31 84:29]
  wire [3:0] _GEN_2531 = tlb_stall ? 4'h0 : _GEN_2123; // @[DCache.scala 263:31 84:29]
  wire [31:0] _GEN_2532 = tlb_stall ? 32'h0 : _GEN_2124; // @[DCache.scala 263:31 84:29]
  wire  _GEN_2933 = 6'h1 == fence_line_addr ? dirty_1_0 : dirty_0_0; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2934 = 6'h2 == fence_line_addr ? dirty_2_0 : _GEN_2933; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2935 = 6'h3 == fence_line_addr ? dirty_3_0 : _GEN_2934; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2936 = 6'h4 == fence_line_addr ? dirty_4_0 : _GEN_2935; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2937 = 6'h5 == fence_line_addr ? dirty_5_0 : _GEN_2936; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2938 = 6'h6 == fence_line_addr ? dirty_6_0 : _GEN_2937; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2939 = 6'h7 == fence_line_addr ? dirty_7_0 : _GEN_2938; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2940 = 6'h8 == fence_line_addr ? dirty_8_0 : _GEN_2939; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2941 = 6'h9 == fence_line_addr ? dirty_9_0 : _GEN_2940; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2942 = 6'ha == fence_line_addr ? dirty_10_0 : _GEN_2941; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2943 = 6'hb == fence_line_addr ? dirty_11_0 : _GEN_2942; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2944 = 6'hc == fence_line_addr ? dirty_12_0 : _GEN_2943; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2945 = 6'hd == fence_line_addr ? dirty_13_0 : _GEN_2944; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2946 = 6'he == fence_line_addr ? dirty_14_0 : _GEN_2945; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2947 = 6'hf == fence_line_addr ? dirty_15_0 : _GEN_2946; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2948 = 6'h10 == fence_line_addr ? dirty_16_0 : _GEN_2947; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2949 = 6'h11 == fence_line_addr ? dirty_17_0 : _GEN_2948; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2950 = 6'h12 == fence_line_addr ? dirty_18_0 : _GEN_2949; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2951 = 6'h13 == fence_line_addr ? dirty_19_0 : _GEN_2950; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2952 = 6'h14 == fence_line_addr ? dirty_20_0 : _GEN_2951; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2953 = 6'h15 == fence_line_addr ? dirty_21_0 : _GEN_2952; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2954 = 6'h16 == fence_line_addr ? dirty_22_0 : _GEN_2953; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2955 = 6'h17 == fence_line_addr ? dirty_23_0 : _GEN_2954; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2956 = 6'h18 == fence_line_addr ? dirty_24_0 : _GEN_2955; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2957 = 6'h19 == fence_line_addr ? dirty_25_0 : _GEN_2956; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2958 = 6'h1a == fence_line_addr ? dirty_26_0 : _GEN_2957; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2959 = 6'h1b == fence_line_addr ? dirty_27_0 : _GEN_2958; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2960 = 6'h1c == fence_line_addr ? dirty_28_0 : _GEN_2959; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2961 = 6'h1d == fence_line_addr ? dirty_29_0 : _GEN_2960; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2962 = 6'h1e == fence_line_addr ? dirty_30_0 : _GEN_2961; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2963 = 6'h1f == fence_line_addr ? dirty_31_0 : _GEN_2962; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2964 = 6'h20 == fence_line_addr ? dirty_32_0 : _GEN_2963; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2965 = 6'h21 == fence_line_addr ? dirty_33_0 : _GEN_2964; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2966 = 6'h22 == fence_line_addr ? dirty_34_0 : _GEN_2965; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2967 = 6'h23 == fence_line_addr ? dirty_35_0 : _GEN_2966; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2968 = 6'h24 == fence_line_addr ? dirty_36_0 : _GEN_2967; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2969 = 6'h25 == fence_line_addr ? dirty_37_0 : _GEN_2968; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2970 = 6'h26 == fence_line_addr ? dirty_38_0 : _GEN_2969; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2971 = 6'h27 == fence_line_addr ? dirty_39_0 : _GEN_2970; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2972 = 6'h28 == fence_line_addr ? dirty_40_0 : _GEN_2971; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2973 = 6'h29 == fence_line_addr ? dirty_41_0 : _GEN_2972; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2974 = 6'h2a == fence_line_addr ? dirty_42_0 : _GEN_2973; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2975 = 6'h2b == fence_line_addr ? dirty_43_0 : _GEN_2974; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2976 = 6'h2c == fence_line_addr ? dirty_44_0 : _GEN_2975; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2977 = 6'h2d == fence_line_addr ? dirty_45_0 : _GEN_2976; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2978 = 6'h2e == fence_line_addr ? dirty_46_0 : _GEN_2977; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2979 = 6'h2f == fence_line_addr ? dirty_47_0 : _GEN_2978; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2980 = 6'h30 == fence_line_addr ? dirty_48_0 : _GEN_2979; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2981 = 6'h31 == fence_line_addr ? dirty_49_0 : _GEN_2980; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2982 = 6'h32 == fence_line_addr ? dirty_50_0 : _GEN_2981; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2983 = 6'h33 == fence_line_addr ? dirty_51_0 : _GEN_2982; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2984 = 6'h34 == fence_line_addr ? dirty_52_0 : _GEN_2983; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2985 = 6'h35 == fence_line_addr ? dirty_53_0 : _GEN_2984; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2986 = 6'h36 == fence_line_addr ? dirty_54_0 : _GEN_2985; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2987 = 6'h37 == fence_line_addr ? dirty_55_0 : _GEN_2986; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2988 = 6'h38 == fence_line_addr ? dirty_56_0 : _GEN_2987; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2989 = 6'h39 == fence_line_addr ? dirty_57_0 : _GEN_2988; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2990 = 6'h3a == fence_line_addr ? dirty_58_0 : _GEN_2989; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2991 = 6'h3b == fence_line_addr ? dirty_59_0 : _GEN_2990; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2992 = 6'h3c == fence_line_addr ? dirty_60_0 : _GEN_2991; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2993 = 6'h3d == fence_line_addr ? dirty_61_0 : _GEN_2992; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2994 = 6'h3e == fence_line_addr ? dirty_62_0 : _GEN_2993; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2995 = 6'h3f == fence_line_addr ? dirty_63_0 : _GEN_2994; // @[DCache.scala 323:{45,45}]
  wire [6:0] _GEN_13029 = {{1'd0}, fence_line_addr}; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2996 = 7'h40 == _GEN_13029 ? dirty_64_0 : _GEN_2995; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2997 = 7'h41 == _GEN_13029 ? dirty_65_0 : _GEN_2996; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2998 = 7'h42 == _GEN_13029 ? dirty_66_0 : _GEN_2997; // @[DCache.scala 323:{45,45}]
  wire  _GEN_2999 = 7'h43 == _GEN_13029 ? dirty_67_0 : _GEN_2998; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3000 = 7'h44 == _GEN_13029 ? dirty_68_0 : _GEN_2999; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3001 = 7'h45 == _GEN_13029 ? dirty_69_0 : _GEN_3000; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3002 = 7'h46 == _GEN_13029 ? dirty_70_0 : _GEN_3001; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3003 = 7'h47 == _GEN_13029 ? dirty_71_0 : _GEN_3002; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3004 = 7'h48 == _GEN_13029 ? dirty_72_0 : _GEN_3003; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3005 = 7'h49 == _GEN_13029 ? dirty_73_0 : _GEN_3004; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3006 = 7'h4a == _GEN_13029 ? dirty_74_0 : _GEN_3005; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3007 = 7'h4b == _GEN_13029 ? dirty_75_0 : _GEN_3006; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3008 = 7'h4c == _GEN_13029 ? dirty_76_0 : _GEN_3007; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3009 = 7'h4d == _GEN_13029 ? dirty_77_0 : _GEN_3008; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3010 = 7'h4e == _GEN_13029 ? dirty_78_0 : _GEN_3009; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3011 = 7'h4f == _GEN_13029 ? dirty_79_0 : _GEN_3010; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3012 = 7'h50 == _GEN_13029 ? dirty_80_0 : _GEN_3011; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3013 = 7'h51 == _GEN_13029 ? dirty_81_0 : _GEN_3012; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3014 = 7'h52 == _GEN_13029 ? dirty_82_0 : _GEN_3013; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3015 = 7'h53 == _GEN_13029 ? dirty_83_0 : _GEN_3014; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3016 = 7'h54 == _GEN_13029 ? dirty_84_0 : _GEN_3015; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3017 = 7'h55 == _GEN_13029 ? dirty_85_0 : _GEN_3016; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3018 = 7'h56 == _GEN_13029 ? dirty_86_0 : _GEN_3017; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3019 = 7'h57 == _GEN_13029 ? dirty_87_0 : _GEN_3018; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3020 = 7'h58 == _GEN_13029 ? dirty_88_0 : _GEN_3019; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3021 = 7'h59 == _GEN_13029 ? dirty_89_0 : _GEN_3020; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3022 = 7'h5a == _GEN_13029 ? dirty_90_0 : _GEN_3021; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3023 = 7'h5b == _GEN_13029 ? dirty_91_0 : _GEN_3022; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3024 = 7'h5c == _GEN_13029 ? dirty_92_0 : _GEN_3023; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3025 = 7'h5d == _GEN_13029 ? dirty_93_0 : _GEN_3024; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3026 = 7'h5e == _GEN_13029 ? dirty_94_0 : _GEN_3025; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3027 = 7'h5f == _GEN_13029 ? dirty_95_0 : _GEN_3026; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3028 = 7'h60 == _GEN_13029 ? dirty_96_0 : _GEN_3027; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3029 = 7'h61 == _GEN_13029 ? dirty_97_0 : _GEN_3028; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3030 = 7'h62 == _GEN_13029 ? dirty_98_0 : _GEN_3029; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3031 = 7'h63 == _GEN_13029 ? dirty_99_0 : _GEN_3030; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3032 = 7'h64 == _GEN_13029 ? dirty_100_0 : _GEN_3031; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3033 = 7'h65 == _GEN_13029 ? dirty_101_0 : _GEN_3032; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3034 = 7'h66 == _GEN_13029 ? dirty_102_0 : _GEN_3033; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3035 = 7'h67 == _GEN_13029 ? dirty_103_0 : _GEN_3034; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3036 = 7'h68 == _GEN_13029 ? dirty_104_0 : _GEN_3035; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3037 = 7'h69 == _GEN_13029 ? dirty_105_0 : _GEN_3036; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3038 = 7'h6a == _GEN_13029 ? dirty_106_0 : _GEN_3037; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3039 = 7'h6b == _GEN_13029 ? dirty_107_0 : _GEN_3038; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3040 = 7'h6c == _GEN_13029 ? dirty_108_0 : _GEN_3039; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3041 = 7'h6d == _GEN_13029 ? dirty_109_0 : _GEN_3040; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3042 = 7'h6e == _GEN_13029 ? dirty_110_0 : _GEN_3041; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3043 = 7'h6f == _GEN_13029 ? dirty_111_0 : _GEN_3042; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3044 = 7'h70 == _GEN_13029 ? dirty_112_0 : _GEN_3043; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3045 = 7'h71 == _GEN_13029 ? dirty_113_0 : _GEN_3044; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3046 = 7'h72 == _GEN_13029 ? dirty_114_0 : _GEN_3045; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3047 = 7'h73 == _GEN_13029 ? dirty_115_0 : _GEN_3046; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3048 = 7'h74 == _GEN_13029 ? dirty_116_0 : _GEN_3047; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3049 = 7'h75 == _GEN_13029 ? dirty_117_0 : _GEN_3048; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3050 = 7'h76 == _GEN_13029 ? dirty_118_0 : _GEN_3049; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3051 = 7'h77 == _GEN_13029 ? dirty_119_0 : _GEN_3050; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3052 = 7'h78 == _GEN_13029 ? dirty_120_0 : _GEN_3051; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3053 = 7'h79 == _GEN_13029 ? dirty_121_0 : _GEN_3052; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3054 = 7'h7a == _GEN_13029 ? dirty_122_0 : _GEN_3053; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3055 = 7'h7b == _GEN_13029 ? dirty_123_0 : _GEN_3054; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3056 = 7'h7c == _GEN_13029 ? dirty_124_0 : _GEN_3055; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3057 = 7'h7d == _GEN_13029 ? dirty_125_0 : _GEN_3056; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3058 = 7'h7e == _GEN_13029 ? dirty_126_0 : _GEN_3057; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3059 = 7'h7f == _GEN_13029 ? dirty_127_0 : _GEN_3058; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3061 = 6'h1 == fence_line_addr ? dirty_1_1 : dirty_0_1; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3062 = 6'h2 == fence_line_addr ? dirty_2_1 : _GEN_3061; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3063 = 6'h3 == fence_line_addr ? dirty_3_1 : _GEN_3062; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3064 = 6'h4 == fence_line_addr ? dirty_4_1 : _GEN_3063; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3065 = 6'h5 == fence_line_addr ? dirty_5_1 : _GEN_3064; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3066 = 6'h6 == fence_line_addr ? dirty_6_1 : _GEN_3065; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3067 = 6'h7 == fence_line_addr ? dirty_7_1 : _GEN_3066; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3068 = 6'h8 == fence_line_addr ? dirty_8_1 : _GEN_3067; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3069 = 6'h9 == fence_line_addr ? dirty_9_1 : _GEN_3068; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3070 = 6'ha == fence_line_addr ? dirty_10_1 : _GEN_3069; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3071 = 6'hb == fence_line_addr ? dirty_11_1 : _GEN_3070; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3072 = 6'hc == fence_line_addr ? dirty_12_1 : _GEN_3071; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3073 = 6'hd == fence_line_addr ? dirty_13_1 : _GEN_3072; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3074 = 6'he == fence_line_addr ? dirty_14_1 : _GEN_3073; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3075 = 6'hf == fence_line_addr ? dirty_15_1 : _GEN_3074; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3076 = 6'h10 == fence_line_addr ? dirty_16_1 : _GEN_3075; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3077 = 6'h11 == fence_line_addr ? dirty_17_1 : _GEN_3076; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3078 = 6'h12 == fence_line_addr ? dirty_18_1 : _GEN_3077; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3079 = 6'h13 == fence_line_addr ? dirty_19_1 : _GEN_3078; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3080 = 6'h14 == fence_line_addr ? dirty_20_1 : _GEN_3079; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3081 = 6'h15 == fence_line_addr ? dirty_21_1 : _GEN_3080; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3082 = 6'h16 == fence_line_addr ? dirty_22_1 : _GEN_3081; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3083 = 6'h17 == fence_line_addr ? dirty_23_1 : _GEN_3082; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3084 = 6'h18 == fence_line_addr ? dirty_24_1 : _GEN_3083; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3085 = 6'h19 == fence_line_addr ? dirty_25_1 : _GEN_3084; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3086 = 6'h1a == fence_line_addr ? dirty_26_1 : _GEN_3085; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3087 = 6'h1b == fence_line_addr ? dirty_27_1 : _GEN_3086; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3088 = 6'h1c == fence_line_addr ? dirty_28_1 : _GEN_3087; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3089 = 6'h1d == fence_line_addr ? dirty_29_1 : _GEN_3088; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3090 = 6'h1e == fence_line_addr ? dirty_30_1 : _GEN_3089; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3091 = 6'h1f == fence_line_addr ? dirty_31_1 : _GEN_3090; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3092 = 6'h20 == fence_line_addr ? dirty_32_1 : _GEN_3091; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3093 = 6'h21 == fence_line_addr ? dirty_33_1 : _GEN_3092; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3094 = 6'h22 == fence_line_addr ? dirty_34_1 : _GEN_3093; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3095 = 6'h23 == fence_line_addr ? dirty_35_1 : _GEN_3094; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3096 = 6'h24 == fence_line_addr ? dirty_36_1 : _GEN_3095; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3097 = 6'h25 == fence_line_addr ? dirty_37_1 : _GEN_3096; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3098 = 6'h26 == fence_line_addr ? dirty_38_1 : _GEN_3097; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3099 = 6'h27 == fence_line_addr ? dirty_39_1 : _GEN_3098; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3100 = 6'h28 == fence_line_addr ? dirty_40_1 : _GEN_3099; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3101 = 6'h29 == fence_line_addr ? dirty_41_1 : _GEN_3100; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3102 = 6'h2a == fence_line_addr ? dirty_42_1 : _GEN_3101; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3103 = 6'h2b == fence_line_addr ? dirty_43_1 : _GEN_3102; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3104 = 6'h2c == fence_line_addr ? dirty_44_1 : _GEN_3103; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3105 = 6'h2d == fence_line_addr ? dirty_45_1 : _GEN_3104; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3106 = 6'h2e == fence_line_addr ? dirty_46_1 : _GEN_3105; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3107 = 6'h2f == fence_line_addr ? dirty_47_1 : _GEN_3106; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3108 = 6'h30 == fence_line_addr ? dirty_48_1 : _GEN_3107; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3109 = 6'h31 == fence_line_addr ? dirty_49_1 : _GEN_3108; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3110 = 6'h32 == fence_line_addr ? dirty_50_1 : _GEN_3109; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3111 = 6'h33 == fence_line_addr ? dirty_51_1 : _GEN_3110; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3112 = 6'h34 == fence_line_addr ? dirty_52_1 : _GEN_3111; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3113 = 6'h35 == fence_line_addr ? dirty_53_1 : _GEN_3112; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3114 = 6'h36 == fence_line_addr ? dirty_54_1 : _GEN_3113; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3115 = 6'h37 == fence_line_addr ? dirty_55_1 : _GEN_3114; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3116 = 6'h38 == fence_line_addr ? dirty_56_1 : _GEN_3115; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3117 = 6'h39 == fence_line_addr ? dirty_57_1 : _GEN_3116; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3118 = 6'h3a == fence_line_addr ? dirty_58_1 : _GEN_3117; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3119 = 6'h3b == fence_line_addr ? dirty_59_1 : _GEN_3118; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3120 = 6'h3c == fence_line_addr ? dirty_60_1 : _GEN_3119; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3121 = 6'h3d == fence_line_addr ? dirty_61_1 : _GEN_3120; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3122 = 6'h3e == fence_line_addr ? dirty_62_1 : _GEN_3121; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3123 = 6'h3f == fence_line_addr ? dirty_63_1 : _GEN_3122; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3124 = 7'h40 == _GEN_13029 ? dirty_64_1 : _GEN_3123; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3125 = 7'h41 == _GEN_13029 ? dirty_65_1 : _GEN_3124; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3126 = 7'h42 == _GEN_13029 ? dirty_66_1 : _GEN_3125; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3127 = 7'h43 == _GEN_13029 ? dirty_67_1 : _GEN_3126; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3128 = 7'h44 == _GEN_13029 ? dirty_68_1 : _GEN_3127; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3129 = 7'h45 == _GEN_13029 ? dirty_69_1 : _GEN_3128; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3130 = 7'h46 == _GEN_13029 ? dirty_70_1 : _GEN_3129; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3131 = 7'h47 == _GEN_13029 ? dirty_71_1 : _GEN_3130; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3132 = 7'h48 == _GEN_13029 ? dirty_72_1 : _GEN_3131; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3133 = 7'h49 == _GEN_13029 ? dirty_73_1 : _GEN_3132; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3134 = 7'h4a == _GEN_13029 ? dirty_74_1 : _GEN_3133; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3135 = 7'h4b == _GEN_13029 ? dirty_75_1 : _GEN_3134; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3136 = 7'h4c == _GEN_13029 ? dirty_76_1 : _GEN_3135; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3137 = 7'h4d == _GEN_13029 ? dirty_77_1 : _GEN_3136; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3138 = 7'h4e == _GEN_13029 ? dirty_78_1 : _GEN_3137; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3139 = 7'h4f == _GEN_13029 ? dirty_79_1 : _GEN_3138; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3140 = 7'h50 == _GEN_13029 ? dirty_80_1 : _GEN_3139; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3141 = 7'h51 == _GEN_13029 ? dirty_81_1 : _GEN_3140; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3142 = 7'h52 == _GEN_13029 ? dirty_82_1 : _GEN_3141; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3143 = 7'h53 == _GEN_13029 ? dirty_83_1 : _GEN_3142; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3144 = 7'h54 == _GEN_13029 ? dirty_84_1 : _GEN_3143; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3145 = 7'h55 == _GEN_13029 ? dirty_85_1 : _GEN_3144; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3146 = 7'h56 == _GEN_13029 ? dirty_86_1 : _GEN_3145; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3147 = 7'h57 == _GEN_13029 ? dirty_87_1 : _GEN_3146; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3148 = 7'h58 == _GEN_13029 ? dirty_88_1 : _GEN_3147; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3149 = 7'h59 == _GEN_13029 ? dirty_89_1 : _GEN_3148; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3150 = 7'h5a == _GEN_13029 ? dirty_90_1 : _GEN_3149; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3151 = 7'h5b == _GEN_13029 ? dirty_91_1 : _GEN_3150; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3152 = 7'h5c == _GEN_13029 ? dirty_92_1 : _GEN_3151; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3153 = 7'h5d == _GEN_13029 ? dirty_93_1 : _GEN_3152; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3154 = 7'h5e == _GEN_13029 ? dirty_94_1 : _GEN_3153; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3155 = 7'h5f == _GEN_13029 ? dirty_95_1 : _GEN_3154; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3156 = 7'h60 == _GEN_13029 ? dirty_96_1 : _GEN_3155; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3157 = 7'h61 == _GEN_13029 ? dirty_97_1 : _GEN_3156; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3158 = 7'h62 == _GEN_13029 ? dirty_98_1 : _GEN_3157; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3159 = 7'h63 == _GEN_13029 ? dirty_99_1 : _GEN_3158; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3160 = 7'h64 == _GEN_13029 ? dirty_100_1 : _GEN_3159; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3161 = 7'h65 == _GEN_13029 ? dirty_101_1 : _GEN_3160; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3162 = 7'h66 == _GEN_13029 ? dirty_102_1 : _GEN_3161; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3163 = 7'h67 == _GEN_13029 ? dirty_103_1 : _GEN_3162; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3164 = 7'h68 == _GEN_13029 ? dirty_104_1 : _GEN_3163; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3165 = 7'h69 == _GEN_13029 ? dirty_105_1 : _GEN_3164; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3166 = 7'h6a == _GEN_13029 ? dirty_106_1 : _GEN_3165; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3167 = 7'h6b == _GEN_13029 ? dirty_107_1 : _GEN_3166; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3168 = 7'h6c == _GEN_13029 ? dirty_108_1 : _GEN_3167; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3169 = 7'h6d == _GEN_13029 ? dirty_109_1 : _GEN_3168; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3170 = 7'h6e == _GEN_13029 ? dirty_110_1 : _GEN_3169; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3171 = 7'h6f == _GEN_13029 ? dirty_111_1 : _GEN_3170; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3172 = 7'h70 == _GEN_13029 ? dirty_112_1 : _GEN_3171; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3173 = 7'h71 == _GEN_13029 ? dirty_113_1 : _GEN_3172; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3174 = 7'h72 == _GEN_13029 ? dirty_114_1 : _GEN_3173; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3175 = 7'h73 == _GEN_13029 ? dirty_115_1 : _GEN_3174; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3176 = 7'h74 == _GEN_13029 ? dirty_116_1 : _GEN_3175; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3177 = 7'h75 == _GEN_13029 ? dirty_117_1 : _GEN_3176; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3178 = 7'h76 == _GEN_13029 ? dirty_118_1 : _GEN_3177; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3179 = 7'h77 == _GEN_13029 ? dirty_119_1 : _GEN_3178; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3180 = 7'h78 == _GEN_13029 ? dirty_120_1 : _GEN_3179; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3181 = 7'h79 == _GEN_13029 ? dirty_121_1 : _GEN_3180; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3182 = 7'h7a == _GEN_13029 ? dirty_122_1 : _GEN_3181; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3183 = 7'h7b == _GEN_13029 ? dirty_123_1 : _GEN_3182; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3184 = 7'h7c == _GEN_13029 ? dirty_124_1 : _GEN_3183; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3185 = 7'h7d == _GEN_13029 ? dirty_125_1 : _GEN_3184; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3186 = 7'h7e == _GEN_13029 ? dirty_126_1 : _GEN_3185; // @[DCache.scala 323:{45,45}]
  wire  _GEN_3187 = 7'h7f == _GEN_13029 ? dirty_127_1 : _GEN_3186; // @[DCache.scala 323:{45,45}]
  wire [9:0] _bram_replace_addr_T_2 = {fence_line_addr,4'h0}; // @[Cat.scala 33:92]
  wire [2:0] _GEN_3188 = _T_12 ? 3'h3 : state; // @[DCache.scala 324:71 325:35 65:96]
  wire [3:0] _GEN_3189 = _T_12 ? 4'h0 : axi_wcnt; // @[DCache.scala 324:71 326:35 89:40]
  wire [9:0] _GEN_3190 = _T_12 ? _bram_replace_addr_T_2 : bram_replace_addr; // @[DCache.scala 324:71 327:35 90:40]
  wire [9:0] _GEN_3191 = _T_12 ? _bram_replace_addr_T_2 : bram_read_ready_addr; // @[DCache.scala 324:71 328:35 91:40]
  wire  _GEN_3193 = _T_12 | bram_use_replace_addr; // @[DCache.scala 324:71 330:35 95:40]
  wire  _GEN_3196 = 6'h1 == fence_line_addr ? valid_1_0 : valid_0_0; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3197 = 6'h2 == fence_line_addr ? valid_2_0 : _GEN_3196; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3198 = 6'h3 == fence_line_addr ? valid_3_0 : _GEN_3197; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3199 = 6'h4 == fence_line_addr ? valid_4_0 : _GEN_3198; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3200 = 6'h5 == fence_line_addr ? valid_5_0 : _GEN_3199; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3201 = 6'h6 == fence_line_addr ? valid_6_0 : _GEN_3200; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3202 = 6'h7 == fence_line_addr ? valid_7_0 : _GEN_3201; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3203 = 6'h8 == fence_line_addr ? valid_8_0 : _GEN_3202; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3204 = 6'h9 == fence_line_addr ? valid_9_0 : _GEN_3203; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3205 = 6'ha == fence_line_addr ? valid_10_0 : _GEN_3204; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3206 = 6'hb == fence_line_addr ? valid_11_0 : _GEN_3205; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3207 = 6'hc == fence_line_addr ? valid_12_0 : _GEN_3206; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3208 = 6'hd == fence_line_addr ? valid_13_0 : _GEN_3207; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3209 = 6'he == fence_line_addr ? valid_14_0 : _GEN_3208; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3210 = 6'hf == fence_line_addr ? valid_15_0 : _GEN_3209; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3211 = 6'h10 == fence_line_addr ? valid_16_0 : _GEN_3210; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3212 = 6'h11 == fence_line_addr ? valid_17_0 : _GEN_3211; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3213 = 6'h12 == fence_line_addr ? valid_18_0 : _GEN_3212; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3214 = 6'h13 == fence_line_addr ? valid_19_0 : _GEN_3213; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3215 = 6'h14 == fence_line_addr ? valid_20_0 : _GEN_3214; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3216 = 6'h15 == fence_line_addr ? valid_21_0 : _GEN_3215; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3217 = 6'h16 == fence_line_addr ? valid_22_0 : _GEN_3216; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3218 = 6'h17 == fence_line_addr ? valid_23_0 : _GEN_3217; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3219 = 6'h18 == fence_line_addr ? valid_24_0 : _GEN_3218; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3220 = 6'h19 == fence_line_addr ? valid_25_0 : _GEN_3219; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3221 = 6'h1a == fence_line_addr ? valid_26_0 : _GEN_3220; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3222 = 6'h1b == fence_line_addr ? valid_27_0 : _GEN_3221; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3223 = 6'h1c == fence_line_addr ? valid_28_0 : _GEN_3222; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3224 = 6'h1d == fence_line_addr ? valid_29_0 : _GEN_3223; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3225 = 6'h1e == fence_line_addr ? valid_30_0 : _GEN_3224; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3226 = 6'h1f == fence_line_addr ? valid_31_0 : _GEN_3225; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3227 = 6'h20 == fence_line_addr ? valid_32_0 : _GEN_3226; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3228 = 6'h21 == fence_line_addr ? valid_33_0 : _GEN_3227; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3229 = 6'h22 == fence_line_addr ? valid_34_0 : _GEN_3228; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3230 = 6'h23 == fence_line_addr ? valid_35_0 : _GEN_3229; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3231 = 6'h24 == fence_line_addr ? valid_36_0 : _GEN_3230; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3232 = 6'h25 == fence_line_addr ? valid_37_0 : _GEN_3231; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3233 = 6'h26 == fence_line_addr ? valid_38_0 : _GEN_3232; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3234 = 6'h27 == fence_line_addr ? valid_39_0 : _GEN_3233; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3235 = 6'h28 == fence_line_addr ? valid_40_0 : _GEN_3234; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3236 = 6'h29 == fence_line_addr ? valid_41_0 : _GEN_3235; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3237 = 6'h2a == fence_line_addr ? valid_42_0 : _GEN_3236; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3238 = 6'h2b == fence_line_addr ? valid_43_0 : _GEN_3237; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3239 = 6'h2c == fence_line_addr ? valid_44_0 : _GEN_3238; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3240 = 6'h2d == fence_line_addr ? valid_45_0 : _GEN_3239; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3241 = 6'h2e == fence_line_addr ? valid_46_0 : _GEN_3240; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3242 = 6'h2f == fence_line_addr ? valid_47_0 : _GEN_3241; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3243 = 6'h30 == fence_line_addr ? valid_48_0 : _GEN_3242; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3244 = 6'h31 == fence_line_addr ? valid_49_0 : _GEN_3243; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3245 = 6'h32 == fence_line_addr ? valid_50_0 : _GEN_3244; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3246 = 6'h33 == fence_line_addr ? valid_51_0 : _GEN_3245; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3247 = 6'h34 == fence_line_addr ? valid_52_0 : _GEN_3246; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3248 = 6'h35 == fence_line_addr ? valid_53_0 : _GEN_3247; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3249 = 6'h36 == fence_line_addr ? valid_54_0 : _GEN_3248; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3250 = 6'h37 == fence_line_addr ? valid_55_0 : _GEN_3249; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3251 = 6'h38 == fence_line_addr ? valid_56_0 : _GEN_3250; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3252 = 6'h39 == fence_line_addr ? valid_57_0 : _GEN_3251; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3253 = 6'h3a == fence_line_addr ? valid_58_0 : _GEN_3252; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3254 = 6'h3b == fence_line_addr ? valid_59_0 : _GEN_3253; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3255 = 6'h3c == fence_line_addr ? valid_60_0 : _GEN_3254; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3256 = 6'h3d == fence_line_addr ? valid_61_0 : _GEN_3255; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3257 = 6'h3e == fence_line_addr ? valid_62_0 : _GEN_3256; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3258 = 6'h3f == fence_line_addr ? valid_63_0 : _GEN_3257; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3259 = 7'h40 == _GEN_13029 ? valid_64_0 : _GEN_3258; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3260 = 7'h41 == _GEN_13029 ? valid_65_0 : _GEN_3259; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3261 = 7'h42 == _GEN_13029 ? valid_66_0 : _GEN_3260; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3262 = 7'h43 == _GEN_13029 ? valid_67_0 : _GEN_3261; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3263 = 7'h44 == _GEN_13029 ? valid_68_0 : _GEN_3262; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3264 = 7'h45 == _GEN_13029 ? valid_69_0 : _GEN_3263; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3265 = 7'h46 == _GEN_13029 ? valid_70_0 : _GEN_3264; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3266 = 7'h47 == _GEN_13029 ? valid_71_0 : _GEN_3265; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3267 = 7'h48 == _GEN_13029 ? valid_72_0 : _GEN_3266; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3268 = 7'h49 == _GEN_13029 ? valid_73_0 : _GEN_3267; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3269 = 7'h4a == _GEN_13029 ? valid_74_0 : _GEN_3268; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3270 = 7'h4b == _GEN_13029 ? valid_75_0 : _GEN_3269; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3271 = 7'h4c == _GEN_13029 ? valid_76_0 : _GEN_3270; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3272 = 7'h4d == _GEN_13029 ? valid_77_0 : _GEN_3271; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3273 = 7'h4e == _GEN_13029 ? valid_78_0 : _GEN_3272; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3274 = 7'h4f == _GEN_13029 ? valid_79_0 : _GEN_3273; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3275 = 7'h50 == _GEN_13029 ? valid_80_0 : _GEN_3274; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3276 = 7'h51 == _GEN_13029 ? valid_81_0 : _GEN_3275; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3277 = 7'h52 == _GEN_13029 ? valid_82_0 : _GEN_3276; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3278 = 7'h53 == _GEN_13029 ? valid_83_0 : _GEN_3277; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3279 = 7'h54 == _GEN_13029 ? valid_84_0 : _GEN_3278; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3280 = 7'h55 == _GEN_13029 ? valid_85_0 : _GEN_3279; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3281 = 7'h56 == _GEN_13029 ? valid_86_0 : _GEN_3280; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3282 = 7'h57 == _GEN_13029 ? valid_87_0 : _GEN_3281; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3283 = 7'h58 == _GEN_13029 ? valid_88_0 : _GEN_3282; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3284 = 7'h59 == _GEN_13029 ? valid_89_0 : _GEN_3283; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3285 = 7'h5a == _GEN_13029 ? valid_90_0 : _GEN_3284; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3286 = 7'h5b == _GEN_13029 ? valid_91_0 : _GEN_3285; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3287 = 7'h5c == _GEN_13029 ? valid_92_0 : _GEN_3286; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3288 = 7'h5d == _GEN_13029 ? valid_93_0 : _GEN_3287; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3289 = 7'h5e == _GEN_13029 ? valid_94_0 : _GEN_3288; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3290 = 7'h5f == _GEN_13029 ? valid_95_0 : _GEN_3289; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3291 = 7'h60 == _GEN_13029 ? valid_96_0 : _GEN_3290; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3292 = 7'h61 == _GEN_13029 ? valid_97_0 : _GEN_3291; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3293 = 7'h62 == _GEN_13029 ? valid_98_0 : _GEN_3292; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3294 = 7'h63 == _GEN_13029 ? valid_99_0 : _GEN_3293; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3295 = 7'h64 == _GEN_13029 ? valid_100_0 : _GEN_3294; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3296 = 7'h65 == _GEN_13029 ? valid_101_0 : _GEN_3295; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3297 = 7'h66 == _GEN_13029 ? valid_102_0 : _GEN_3296; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3298 = 7'h67 == _GEN_13029 ? valid_103_0 : _GEN_3297; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3299 = 7'h68 == _GEN_13029 ? valid_104_0 : _GEN_3298; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3300 = 7'h69 == _GEN_13029 ? valid_105_0 : _GEN_3299; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3301 = 7'h6a == _GEN_13029 ? valid_106_0 : _GEN_3300; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3302 = 7'h6b == _GEN_13029 ? valid_107_0 : _GEN_3301; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3303 = 7'h6c == _GEN_13029 ? valid_108_0 : _GEN_3302; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3304 = 7'h6d == _GEN_13029 ? valid_109_0 : _GEN_3303; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3305 = 7'h6e == _GEN_13029 ? valid_110_0 : _GEN_3304; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3306 = 7'h6f == _GEN_13029 ? valid_111_0 : _GEN_3305; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3307 = 7'h70 == _GEN_13029 ? valid_112_0 : _GEN_3306; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3308 = 7'h71 == _GEN_13029 ? valid_113_0 : _GEN_3307; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3309 = 7'h72 == _GEN_13029 ? valid_114_0 : _GEN_3308; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3310 = 7'h73 == _GEN_13029 ? valid_115_0 : _GEN_3309; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3311 = 7'h74 == _GEN_13029 ? valid_116_0 : _GEN_3310; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3312 = 7'h75 == _GEN_13029 ? valid_117_0 : _GEN_3311; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3313 = 7'h76 == _GEN_13029 ? valid_118_0 : _GEN_3312; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3314 = 7'h77 == _GEN_13029 ? valid_119_0 : _GEN_3313; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3315 = 7'h78 == _GEN_13029 ? valid_120_0 : _GEN_3314; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3316 = 7'h79 == _GEN_13029 ? valid_121_0 : _GEN_3315; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3317 = 7'h7a == _GEN_13029 ? valid_122_0 : _GEN_3316; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3318 = 7'h7b == _GEN_13029 ? valid_123_0 : _GEN_3317; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3319 = 7'h7c == _GEN_13029 ? valid_124_0 : _GEN_3318; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3320 = 7'h7d == _GEN_13029 ? valid_125_0 : _GEN_3319; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3321 = 7'h7e == _GEN_13029 ? valid_126_0 : _GEN_3320; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3322 = 7'h7f == _GEN_13029 ? valid_127_0 : _GEN_3321; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3324 = 6'h1 == fence_line_addr ? valid_1_1 : valid_0_1; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3325 = 6'h2 == fence_line_addr ? valid_2_1 : _GEN_3324; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3326 = 6'h3 == fence_line_addr ? valid_3_1 : _GEN_3325; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3327 = 6'h4 == fence_line_addr ? valid_4_1 : _GEN_3326; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3328 = 6'h5 == fence_line_addr ? valid_5_1 : _GEN_3327; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3329 = 6'h6 == fence_line_addr ? valid_6_1 : _GEN_3328; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3330 = 6'h7 == fence_line_addr ? valid_7_1 : _GEN_3329; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3331 = 6'h8 == fence_line_addr ? valid_8_1 : _GEN_3330; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3332 = 6'h9 == fence_line_addr ? valid_9_1 : _GEN_3331; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3333 = 6'ha == fence_line_addr ? valid_10_1 : _GEN_3332; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3334 = 6'hb == fence_line_addr ? valid_11_1 : _GEN_3333; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3335 = 6'hc == fence_line_addr ? valid_12_1 : _GEN_3334; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3336 = 6'hd == fence_line_addr ? valid_13_1 : _GEN_3335; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3337 = 6'he == fence_line_addr ? valid_14_1 : _GEN_3336; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3338 = 6'hf == fence_line_addr ? valid_15_1 : _GEN_3337; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3339 = 6'h10 == fence_line_addr ? valid_16_1 : _GEN_3338; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3340 = 6'h11 == fence_line_addr ? valid_17_1 : _GEN_3339; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3341 = 6'h12 == fence_line_addr ? valid_18_1 : _GEN_3340; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3342 = 6'h13 == fence_line_addr ? valid_19_1 : _GEN_3341; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3343 = 6'h14 == fence_line_addr ? valid_20_1 : _GEN_3342; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3344 = 6'h15 == fence_line_addr ? valid_21_1 : _GEN_3343; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3345 = 6'h16 == fence_line_addr ? valid_22_1 : _GEN_3344; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3346 = 6'h17 == fence_line_addr ? valid_23_1 : _GEN_3345; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3347 = 6'h18 == fence_line_addr ? valid_24_1 : _GEN_3346; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3348 = 6'h19 == fence_line_addr ? valid_25_1 : _GEN_3347; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3349 = 6'h1a == fence_line_addr ? valid_26_1 : _GEN_3348; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3350 = 6'h1b == fence_line_addr ? valid_27_1 : _GEN_3349; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3351 = 6'h1c == fence_line_addr ? valid_28_1 : _GEN_3350; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3352 = 6'h1d == fence_line_addr ? valid_29_1 : _GEN_3351; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3353 = 6'h1e == fence_line_addr ? valid_30_1 : _GEN_3352; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3354 = 6'h1f == fence_line_addr ? valid_31_1 : _GEN_3353; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3355 = 6'h20 == fence_line_addr ? valid_32_1 : _GEN_3354; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3356 = 6'h21 == fence_line_addr ? valid_33_1 : _GEN_3355; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3357 = 6'h22 == fence_line_addr ? valid_34_1 : _GEN_3356; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3358 = 6'h23 == fence_line_addr ? valid_35_1 : _GEN_3357; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3359 = 6'h24 == fence_line_addr ? valid_36_1 : _GEN_3358; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3360 = 6'h25 == fence_line_addr ? valid_37_1 : _GEN_3359; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3361 = 6'h26 == fence_line_addr ? valid_38_1 : _GEN_3360; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3362 = 6'h27 == fence_line_addr ? valid_39_1 : _GEN_3361; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3363 = 6'h28 == fence_line_addr ? valid_40_1 : _GEN_3362; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3364 = 6'h29 == fence_line_addr ? valid_41_1 : _GEN_3363; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3365 = 6'h2a == fence_line_addr ? valid_42_1 : _GEN_3364; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3366 = 6'h2b == fence_line_addr ? valid_43_1 : _GEN_3365; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3367 = 6'h2c == fence_line_addr ? valid_44_1 : _GEN_3366; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3368 = 6'h2d == fence_line_addr ? valid_45_1 : _GEN_3367; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3369 = 6'h2e == fence_line_addr ? valid_46_1 : _GEN_3368; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3370 = 6'h2f == fence_line_addr ? valid_47_1 : _GEN_3369; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3371 = 6'h30 == fence_line_addr ? valid_48_1 : _GEN_3370; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3372 = 6'h31 == fence_line_addr ? valid_49_1 : _GEN_3371; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3373 = 6'h32 == fence_line_addr ? valid_50_1 : _GEN_3372; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3374 = 6'h33 == fence_line_addr ? valid_51_1 : _GEN_3373; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3375 = 6'h34 == fence_line_addr ? valid_52_1 : _GEN_3374; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3376 = 6'h35 == fence_line_addr ? valid_53_1 : _GEN_3375; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3377 = 6'h36 == fence_line_addr ? valid_54_1 : _GEN_3376; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3378 = 6'h37 == fence_line_addr ? valid_55_1 : _GEN_3377; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3379 = 6'h38 == fence_line_addr ? valid_56_1 : _GEN_3378; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3380 = 6'h39 == fence_line_addr ? valid_57_1 : _GEN_3379; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3381 = 6'h3a == fence_line_addr ? valid_58_1 : _GEN_3380; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3382 = 6'h3b == fence_line_addr ? valid_59_1 : _GEN_3381; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3383 = 6'h3c == fence_line_addr ? valid_60_1 : _GEN_3382; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3384 = 6'h3d == fence_line_addr ? valid_61_1 : _GEN_3383; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3385 = 6'h3e == fence_line_addr ? valid_62_1 : _GEN_3384; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3386 = 6'h3f == fence_line_addr ? valid_63_1 : _GEN_3385; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3387 = 7'h40 == _GEN_13029 ? valid_64_1 : _GEN_3386; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3388 = 7'h41 == _GEN_13029 ? valid_65_1 : _GEN_3387; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3389 = 7'h42 == _GEN_13029 ? valid_66_1 : _GEN_3388; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3390 = 7'h43 == _GEN_13029 ? valid_67_1 : _GEN_3389; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3391 = 7'h44 == _GEN_13029 ? valid_68_1 : _GEN_3390; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3392 = 7'h45 == _GEN_13029 ? valid_69_1 : _GEN_3391; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3393 = 7'h46 == _GEN_13029 ? valid_70_1 : _GEN_3392; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3394 = 7'h47 == _GEN_13029 ? valid_71_1 : _GEN_3393; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3395 = 7'h48 == _GEN_13029 ? valid_72_1 : _GEN_3394; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3396 = 7'h49 == _GEN_13029 ? valid_73_1 : _GEN_3395; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3397 = 7'h4a == _GEN_13029 ? valid_74_1 : _GEN_3396; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3398 = 7'h4b == _GEN_13029 ? valid_75_1 : _GEN_3397; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3399 = 7'h4c == _GEN_13029 ? valid_76_1 : _GEN_3398; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3400 = 7'h4d == _GEN_13029 ? valid_77_1 : _GEN_3399; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3401 = 7'h4e == _GEN_13029 ? valid_78_1 : _GEN_3400; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3402 = 7'h4f == _GEN_13029 ? valid_79_1 : _GEN_3401; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3403 = 7'h50 == _GEN_13029 ? valid_80_1 : _GEN_3402; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3404 = 7'h51 == _GEN_13029 ? valid_81_1 : _GEN_3403; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3405 = 7'h52 == _GEN_13029 ? valid_82_1 : _GEN_3404; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3406 = 7'h53 == _GEN_13029 ? valid_83_1 : _GEN_3405; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3407 = 7'h54 == _GEN_13029 ? valid_84_1 : _GEN_3406; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3408 = 7'h55 == _GEN_13029 ? valid_85_1 : _GEN_3407; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3409 = 7'h56 == _GEN_13029 ? valid_86_1 : _GEN_3408; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3410 = 7'h57 == _GEN_13029 ? valid_87_1 : _GEN_3409; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3411 = 7'h58 == _GEN_13029 ? valid_88_1 : _GEN_3410; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3412 = 7'h59 == _GEN_13029 ? valid_89_1 : _GEN_3411; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3413 = 7'h5a == _GEN_13029 ? valid_90_1 : _GEN_3412; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3414 = 7'h5b == _GEN_13029 ? valid_91_1 : _GEN_3413; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3415 = 7'h5c == _GEN_13029 ? valid_92_1 : _GEN_3414; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3416 = 7'h5d == _GEN_13029 ? valid_93_1 : _GEN_3415; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3417 = 7'h5e == _GEN_13029 ? valid_94_1 : _GEN_3416; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3418 = 7'h5f == _GEN_13029 ? valid_95_1 : _GEN_3417; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3419 = 7'h60 == _GEN_13029 ? valid_96_1 : _GEN_3418; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3420 = 7'h61 == _GEN_13029 ? valid_97_1 : _GEN_3419; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3421 = 7'h62 == _GEN_13029 ? valid_98_1 : _GEN_3420; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3422 = 7'h63 == _GEN_13029 ? valid_99_1 : _GEN_3421; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3423 = 7'h64 == _GEN_13029 ? valid_100_1 : _GEN_3422; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3424 = 7'h65 == _GEN_13029 ? valid_101_1 : _GEN_3423; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3425 = 7'h66 == _GEN_13029 ? valid_102_1 : _GEN_3424; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3426 = 7'h67 == _GEN_13029 ? valid_103_1 : _GEN_3425; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3427 = 7'h68 == _GEN_13029 ? valid_104_1 : _GEN_3426; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3428 = 7'h69 == _GEN_13029 ? valid_105_1 : _GEN_3427; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3429 = 7'h6a == _GEN_13029 ? valid_106_1 : _GEN_3428; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3430 = 7'h6b == _GEN_13029 ? valid_107_1 : _GEN_3429; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3431 = 7'h6c == _GEN_13029 ? valid_108_1 : _GEN_3430; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3432 = 7'h6d == _GEN_13029 ? valid_109_1 : _GEN_3431; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3433 = 7'h6e == _GEN_13029 ? valid_110_1 : _GEN_3432; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3434 = 7'h6f == _GEN_13029 ? valid_111_1 : _GEN_3433; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3435 = 7'h70 == _GEN_13029 ? valid_112_1 : _GEN_3434; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3436 = 7'h71 == _GEN_13029 ? valid_113_1 : _GEN_3435; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3437 = 7'h72 == _GEN_13029 ? valid_114_1 : _GEN_3436; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3438 = 7'h73 == _GEN_13029 ? valid_115_1 : _GEN_3437; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3439 = 7'h74 == _GEN_13029 ? valid_116_1 : _GEN_3438; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3440 = 7'h75 == _GEN_13029 ? valid_117_1 : _GEN_3439; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3441 = 7'h76 == _GEN_13029 ? valid_118_1 : _GEN_3440; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3442 = 7'h77 == _GEN_13029 ? valid_119_1 : _GEN_3441; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3443 = 7'h78 == _GEN_13029 ? valid_120_1 : _GEN_3442; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3444 = 7'h79 == _GEN_13029 ? valid_121_1 : _GEN_3443; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3445 = 7'h7a == _GEN_13029 ? valid_122_1 : _GEN_3444; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3446 = 7'h7b == _GEN_13029 ? valid_123_1 : _GEN_3445; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3447 = 7'h7c == _GEN_13029 ? valid_124_1 : _GEN_3446; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3448 = 7'h7d == _GEN_13029 ? valid_125_1 : _GEN_3447; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3449 = 7'h7e == _GEN_13029 ? valid_126_1 : _GEN_3448; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3450 = 7'h7f == _GEN_13029 ? valid_127_1 : _GEN_3449; // @[DCache.scala 334:{47,47}]
  wire  _GEN_3451 = 6'h0 == fence_line_addr ? 1'h0 : valid_0_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3452 = 6'h1 == fence_line_addr ? 1'h0 : valid_1_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3453 = 6'h2 == fence_line_addr ? 1'h0 : valid_2_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3454 = 6'h3 == fence_line_addr ? 1'h0 : valid_3_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3455 = 6'h4 == fence_line_addr ? 1'h0 : valid_4_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3456 = 6'h5 == fence_line_addr ? 1'h0 : valid_5_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3457 = 6'h6 == fence_line_addr ? 1'h0 : valid_6_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3458 = 6'h7 == fence_line_addr ? 1'h0 : valid_7_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3459 = 6'h8 == fence_line_addr ? 1'h0 : valid_8_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3460 = 6'h9 == fence_line_addr ? 1'h0 : valid_9_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3461 = 6'ha == fence_line_addr ? 1'h0 : valid_10_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3462 = 6'hb == fence_line_addr ? 1'h0 : valid_11_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3463 = 6'hc == fence_line_addr ? 1'h0 : valid_12_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3464 = 6'hd == fence_line_addr ? 1'h0 : valid_13_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3465 = 6'he == fence_line_addr ? 1'h0 : valid_14_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3466 = 6'hf == fence_line_addr ? 1'h0 : valid_15_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3467 = 6'h10 == fence_line_addr ? 1'h0 : valid_16_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3468 = 6'h11 == fence_line_addr ? 1'h0 : valid_17_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3469 = 6'h12 == fence_line_addr ? 1'h0 : valid_18_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3470 = 6'h13 == fence_line_addr ? 1'h0 : valid_19_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3471 = 6'h14 == fence_line_addr ? 1'h0 : valid_20_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3472 = 6'h15 == fence_line_addr ? 1'h0 : valid_21_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3473 = 6'h16 == fence_line_addr ? 1'h0 : valid_22_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3474 = 6'h17 == fence_line_addr ? 1'h0 : valid_23_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3475 = 6'h18 == fence_line_addr ? 1'h0 : valid_24_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3476 = 6'h19 == fence_line_addr ? 1'h0 : valid_25_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3477 = 6'h1a == fence_line_addr ? 1'h0 : valid_26_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3478 = 6'h1b == fence_line_addr ? 1'h0 : valid_27_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3479 = 6'h1c == fence_line_addr ? 1'h0 : valid_28_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3480 = 6'h1d == fence_line_addr ? 1'h0 : valid_29_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3481 = 6'h1e == fence_line_addr ? 1'h0 : valid_30_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3482 = 6'h1f == fence_line_addr ? 1'h0 : valid_31_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3483 = 6'h20 == fence_line_addr ? 1'h0 : valid_32_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3484 = 6'h21 == fence_line_addr ? 1'h0 : valid_33_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3485 = 6'h22 == fence_line_addr ? 1'h0 : valid_34_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3486 = 6'h23 == fence_line_addr ? 1'h0 : valid_35_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3487 = 6'h24 == fence_line_addr ? 1'h0 : valid_36_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3488 = 6'h25 == fence_line_addr ? 1'h0 : valid_37_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3489 = 6'h26 == fence_line_addr ? 1'h0 : valid_38_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3490 = 6'h27 == fence_line_addr ? 1'h0 : valid_39_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3491 = 6'h28 == fence_line_addr ? 1'h0 : valid_40_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3492 = 6'h29 == fence_line_addr ? 1'h0 : valid_41_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3493 = 6'h2a == fence_line_addr ? 1'h0 : valid_42_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3494 = 6'h2b == fence_line_addr ? 1'h0 : valid_43_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3495 = 6'h2c == fence_line_addr ? 1'h0 : valid_44_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3496 = 6'h2d == fence_line_addr ? 1'h0 : valid_45_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3497 = 6'h2e == fence_line_addr ? 1'h0 : valid_46_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3498 = 6'h2f == fence_line_addr ? 1'h0 : valid_47_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3499 = 6'h30 == fence_line_addr ? 1'h0 : valid_48_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3500 = 6'h31 == fence_line_addr ? 1'h0 : valid_49_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3501 = 6'h32 == fence_line_addr ? 1'h0 : valid_50_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3502 = 6'h33 == fence_line_addr ? 1'h0 : valid_51_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3503 = 6'h34 == fence_line_addr ? 1'h0 : valid_52_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3504 = 6'h35 == fence_line_addr ? 1'h0 : valid_53_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3505 = 6'h36 == fence_line_addr ? 1'h0 : valid_54_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3506 = 6'h37 == fence_line_addr ? 1'h0 : valid_55_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3507 = 6'h38 == fence_line_addr ? 1'h0 : valid_56_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3508 = 6'h39 == fence_line_addr ? 1'h0 : valid_57_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3509 = 6'h3a == fence_line_addr ? 1'h0 : valid_58_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3510 = 6'h3b == fence_line_addr ? 1'h0 : valid_59_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3511 = 6'h3c == fence_line_addr ? 1'h0 : valid_60_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3512 = 6'h3d == fence_line_addr ? 1'h0 : valid_61_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3513 = 6'h3e == fence_line_addr ? 1'h0 : valid_62_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3514 = 6'h3f == fence_line_addr ? 1'h0 : valid_63_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3515 = 7'h40 == _GEN_13029 ? 1'h0 : valid_64_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3516 = 7'h41 == _GEN_13029 ? 1'h0 : valid_65_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3517 = 7'h42 == _GEN_13029 ? 1'h0 : valid_66_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3518 = 7'h43 == _GEN_13029 ? 1'h0 : valid_67_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3519 = 7'h44 == _GEN_13029 ? 1'h0 : valid_68_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3520 = 7'h45 == _GEN_13029 ? 1'h0 : valid_69_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3521 = 7'h46 == _GEN_13029 ? 1'h0 : valid_70_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3522 = 7'h47 == _GEN_13029 ? 1'h0 : valid_71_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3523 = 7'h48 == _GEN_13029 ? 1'h0 : valid_72_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3524 = 7'h49 == _GEN_13029 ? 1'h0 : valid_73_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3525 = 7'h4a == _GEN_13029 ? 1'h0 : valid_74_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3526 = 7'h4b == _GEN_13029 ? 1'h0 : valid_75_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3527 = 7'h4c == _GEN_13029 ? 1'h0 : valid_76_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3528 = 7'h4d == _GEN_13029 ? 1'h0 : valid_77_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3529 = 7'h4e == _GEN_13029 ? 1'h0 : valid_78_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3530 = 7'h4f == _GEN_13029 ? 1'h0 : valid_79_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3531 = 7'h50 == _GEN_13029 ? 1'h0 : valid_80_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3532 = 7'h51 == _GEN_13029 ? 1'h0 : valid_81_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3533 = 7'h52 == _GEN_13029 ? 1'h0 : valid_82_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3534 = 7'h53 == _GEN_13029 ? 1'h0 : valid_83_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3535 = 7'h54 == _GEN_13029 ? 1'h0 : valid_84_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3536 = 7'h55 == _GEN_13029 ? 1'h0 : valid_85_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3537 = 7'h56 == _GEN_13029 ? 1'h0 : valid_86_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3538 = 7'h57 == _GEN_13029 ? 1'h0 : valid_87_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3539 = 7'h58 == _GEN_13029 ? 1'h0 : valid_88_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3540 = 7'h59 == _GEN_13029 ? 1'h0 : valid_89_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3541 = 7'h5a == _GEN_13029 ? 1'h0 : valid_90_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3542 = 7'h5b == _GEN_13029 ? 1'h0 : valid_91_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3543 = 7'h5c == _GEN_13029 ? 1'h0 : valid_92_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3544 = 7'h5d == _GEN_13029 ? 1'h0 : valid_93_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3545 = 7'h5e == _GEN_13029 ? 1'h0 : valid_94_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3546 = 7'h5f == _GEN_13029 ? 1'h0 : valid_95_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3547 = 7'h60 == _GEN_13029 ? 1'h0 : valid_96_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3548 = 7'h61 == _GEN_13029 ? 1'h0 : valid_97_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3549 = 7'h62 == _GEN_13029 ? 1'h0 : valid_98_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3550 = 7'h63 == _GEN_13029 ? 1'h0 : valid_99_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3551 = 7'h64 == _GEN_13029 ? 1'h0 : valid_100_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3552 = 7'h65 == _GEN_13029 ? 1'h0 : valid_101_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3553 = 7'h66 == _GEN_13029 ? 1'h0 : valid_102_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3554 = 7'h67 == _GEN_13029 ? 1'h0 : valid_103_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3555 = 7'h68 == _GEN_13029 ? 1'h0 : valid_104_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3556 = 7'h69 == _GEN_13029 ? 1'h0 : valid_105_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3557 = 7'h6a == _GEN_13029 ? 1'h0 : valid_106_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3558 = 7'h6b == _GEN_13029 ? 1'h0 : valid_107_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3559 = 7'h6c == _GEN_13029 ? 1'h0 : valid_108_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3560 = 7'h6d == _GEN_13029 ? 1'h0 : valid_109_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3561 = 7'h6e == _GEN_13029 ? 1'h0 : valid_110_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3562 = 7'h6f == _GEN_13029 ? 1'h0 : valid_111_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3563 = 7'h70 == _GEN_13029 ? 1'h0 : valid_112_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3564 = 7'h71 == _GEN_13029 ? 1'h0 : valid_113_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3565 = 7'h72 == _GEN_13029 ? 1'h0 : valid_114_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3566 = 7'h73 == _GEN_13029 ? 1'h0 : valid_115_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3567 = 7'h74 == _GEN_13029 ? 1'h0 : valid_116_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3568 = 7'h75 == _GEN_13029 ? 1'h0 : valid_117_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3569 = 7'h76 == _GEN_13029 ? 1'h0 : valid_118_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3570 = 7'h77 == _GEN_13029 ? 1'h0 : valid_119_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3571 = 7'h78 == _GEN_13029 ? 1'h0 : valid_120_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3572 = 7'h79 == _GEN_13029 ? 1'h0 : valid_121_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3573 = 7'h7a == _GEN_13029 ? 1'h0 : valid_122_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3574 = 7'h7b == _GEN_13029 ? 1'h0 : valid_123_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3575 = 7'h7c == _GEN_13029 ? 1'h0 : valid_124_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3576 = 7'h7d == _GEN_13029 ? 1'h0 : valid_125_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3577 = 7'h7e == _GEN_13029 ? 1'h0 : valid_126_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3578 = 7'h7f == _GEN_13029 ? 1'h0 : valid_127_0; // @[DCache.scala 335:{39,39} 68:22]
  wire  _GEN_3579 = 6'h0 == fence_line_addr ? 1'h0 : valid_0_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3580 = 6'h1 == fence_line_addr ? 1'h0 : valid_1_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3581 = 6'h2 == fence_line_addr ? 1'h0 : valid_2_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3582 = 6'h3 == fence_line_addr ? 1'h0 : valid_3_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3583 = 6'h4 == fence_line_addr ? 1'h0 : valid_4_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3584 = 6'h5 == fence_line_addr ? 1'h0 : valid_5_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3585 = 6'h6 == fence_line_addr ? 1'h0 : valid_6_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3586 = 6'h7 == fence_line_addr ? 1'h0 : valid_7_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3587 = 6'h8 == fence_line_addr ? 1'h0 : valid_8_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3588 = 6'h9 == fence_line_addr ? 1'h0 : valid_9_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3589 = 6'ha == fence_line_addr ? 1'h0 : valid_10_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3590 = 6'hb == fence_line_addr ? 1'h0 : valid_11_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3591 = 6'hc == fence_line_addr ? 1'h0 : valid_12_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3592 = 6'hd == fence_line_addr ? 1'h0 : valid_13_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3593 = 6'he == fence_line_addr ? 1'h0 : valid_14_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3594 = 6'hf == fence_line_addr ? 1'h0 : valid_15_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3595 = 6'h10 == fence_line_addr ? 1'h0 : valid_16_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3596 = 6'h11 == fence_line_addr ? 1'h0 : valid_17_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3597 = 6'h12 == fence_line_addr ? 1'h0 : valid_18_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3598 = 6'h13 == fence_line_addr ? 1'h0 : valid_19_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3599 = 6'h14 == fence_line_addr ? 1'h0 : valid_20_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3600 = 6'h15 == fence_line_addr ? 1'h0 : valid_21_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3601 = 6'h16 == fence_line_addr ? 1'h0 : valid_22_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3602 = 6'h17 == fence_line_addr ? 1'h0 : valid_23_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3603 = 6'h18 == fence_line_addr ? 1'h0 : valid_24_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3604 = 6'h19 == fence_line_addr ? 1'h0 : valid_25_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3605 = 6'h1a == fence_line_addr ? 1'h0 : valid_26_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3606 = 6'h1b == fence_line_addr ? 1'h0 : valid_27_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3607 = 6'h1c == fence_line_addr ? 1'h0 : valid_28_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3608 = 6'h1d == fence_line_addr ? 1'h0 : valid_29_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3609 = 6'h1e == fence_line_addr ? 1'h0 : valid_30_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3610 = 6'h1f == fence_line_addr ? 1'h0 : valid_31_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3611 = 6'h20 == fence_line_addr ? 1'h0 : valid_32_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3612 = 6'h21 == fence_line_addr ? 1'h0 : valid_33_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3613 = 6'h22 == fence_line_addr ? 1'h0 : valid_34_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3614 = 6'h23 == fence_line_addr ? 1'h0 : valid_35_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3615 = 6'h24 == fence_line_addr ? 1'h0 : valid_36_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3616 = 6'h25 == fence_line_addr ? 1'h0 : valid_37_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3617 = 6'h26 == fence_line_addr ? 1'h0 : valid_38_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3618 = 6'h27 == fence_line_addr ? 1'h0 : valid_39_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3619 = 6'h28 == fence_line_addr ? 1'h0 : valid_40_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3620 = 6'h29 == fence_line_addr ? 1'h0 : valid_41_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3621 = 6'h2a == fence_line_addr ? 1'h0 : valid_42_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3622 = 6'h2b == fence_line_addr ? 1'h0 : valid_43_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3623 = 6'h2c == fence_line_addr ? 1'h0 : valid_44_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3624 = 6'h2d == fence_line_addr ? 1'h0 : valid_45_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3625 = 6'h2e == fence_line_addr ? 1'h0 : valid_46_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3626 = 6'h2f == fence_line_addr ? 1'h0 : valid_47_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3627 = 6'h30 == fence_line_addr ? 1'h0 : valid_48_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3628 = 6'h31 == fence_line_addr ? 1'h0 : valid_49_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3629 = 6'h32 == fence_line_addr ? 1'h0 : valid_50_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3630 = 6'h33 == fence_line_addr ? 1'h0 : valid_51_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3631 = 6'h34 == fence_line_addr ? 1'h0 : valid_52_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3632 = 6'h35 == fence_line_addr ? 1'h0 : valid_53_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3633 = 6'h36 == fence_line_addr ? 1'h0 : valid_54_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3634 = 6'h37 == fence_line_addr ? 1'h0 : valid_55_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3635 = 6'h38 == fence_line_addr ? 1'h0 : valid_56_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3636 = 6'h39 == fence_line_addr ? 1'h0 : valid_57_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3637 = 6'h3a == fence_line_addr ? 1'h0 : valid_58_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3638 = 6'h3b == fence_line_addr ? 1'h0 : valid_59_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3639 = 6'h3c == fence_line_addr ? 1'h0 : valid_60_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3640 = 6'h3d == fence_line_addr ? 1'h0 : valid_61_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3641 = 6'h3e == fence_line_addr ? 1'h0 : valid_62_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3642 = 6'h3f == fence_line_addr ? 1'h0 : valid_63_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3643 = 7'h40 == _GEN_13029 ? 1'h0 : valid_64_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3644 = 7'h41 == _GEN_13029 ? 1'h0 : valid_65_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3645 = 7'h42 == _GEN_13029 ? 1'h0 : valid_66_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3646 = 7'h43 == _GEN_13029 ? 1'h0 : valid_67_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3647 = 7'h44 == _GEN_13029 ? 1'h0 : valid_68_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3648 = 7'h45 == _GEN_13029 ? 1'h0 : valid_69_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3649 = 7'h46 == _GEN_13029 ? 1'h0 : valid_70_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3650 = 7'h47 == _GEN_13029 ? 1'h0 : valid_71_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3651 = 7'h48 == _GEN_13029 ? 1'h0 : valid_72_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3652 = 7'h49 == _GEN_13029 ? 1'h0 : valid_73_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3653 = 7'h4a == _GEN_13029 ? 1'h0 : valid_74_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3654 = 7'h4b == _GEN_13029 ? 1'h0 : valid_75_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3655 = 7'h4c == _GEN_13029 ? 1'h0 : valid_76_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3656 = 7'h4d == _GEN_13029 ? 1'h0 : valid_77_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3657 = 7'h4e == _GEN_13029 ? 1'h0 : valid_78_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3658 = 7'h4f == _GEN_13029 ? 1'h0 : valid_79_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3659 = 7'h50 == _GEN_13029 ? 1'h0 : valid_80_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3660 = 7'h51 == _GEN_13029 ? 1'h0 : valid_81_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3661 = 7'h52 == _GEN_13029 ? 1'h0 : valid_82_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3662 = 7'h53 == _GEN_13029 ? 1'h0 : valid_83_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3663 = 7'h54 == _GEN_13029 ? 1'h0 : valid_84_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3664 = 7'h55 == _GEN_13029 ? 1'h0 : valid_85_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3665 = 7'h56 == _GEN_13029 ? 1'h0 : valid_86_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3666 = 7'h57 == _GEN_13029 ? 1'h0 : valid_87_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3667 = 7'h58 == _GEN_13029 ? 1'h0 : valid_88_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3668 = 7'h59 == _GEN_13029 ? 1'h0 : valid_89_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3669 = 7'h5a == _GEN_13029 ? 1'h0 : valid_90_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3670 = 7'h5b == _GEN_13029 ? 1'h0 : valid_91_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3671 = 7'h5c == _GEN_13029 ? 1'h0 : valid_92_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3672 = 7'h5d == _GEN_13029 ? 1'h0 : valid_93_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3673 = 7'h5e == _GEN_13029 ? 1'h0 : valid_94_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3674 = 7'h5f == _GEN_13029 ? 1'h0 : valid_95_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3675 = 7'h60 == _GEN_13029 ? 1'h0 : valid_96_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3676 = 7'h61 == _GEN_13029 ? 1'h0 : valid_97_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3677 = 7'h62 == _GEN_13029 ? 1'h0 : valid_98_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3678 = 7'h63 == _GEN_13029 ? 1'h0 : valid_99_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3679 = 7'h64 == _GEN_13029 ? 1'h0 : valid_100_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3680 = 7'h65 == _GEN_13029 ? 1'h0 : valid_101_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3681 = 7'h66 == _GEN_13029 ? 1'h0 : valid_102_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3682 = 7'h67 == _GEN_13029 ? 1'h0 : valid_103_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3683 = 7'h68 == _GEN_13029 ? 1'h0 : valid_104_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3684 = 7'h69 == _GEN_13029 ? 1'h0 : valid_105_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3685 = 7'h6a == _GEN_13029 ? 1'h0 : valid_106_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3686 = 7'h6b == _GEN_13029 ? 1'h0 : valid_107_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3687 = 7'h6c == _GEN_13029 ? 1'h0 : valid_108_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3688 = 7'h6d == _GEN_13029 ? 1'h0 : valid_109_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3689 = 7'h6e == _GEN_13029 ? 1'h0 : valid_110_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3690 = 7'h6f == _GEN_13029 ? 1'h0 : valid_111_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3691 = 7'h70 == _GEN_13029 ? 1'h0 : valid_112_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3692 = 7'h71 == _GEN_13029 ? 1'h0 : valid_113_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3693 = 7'h72 == _GEN_13029 ? 1'h0 : valid_114_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3694 = 7'h73 == _GEN_13029 ? 1'h0 : valid_115_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3695 = 7'h74 == _GEN_13029 ? 1'h0 : valid_116_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3696 = 7'h75 == _GEN_13029 ? 1'h0 : valid_117_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3697 = 7'h76 == _GEN_13029 ? 1'h0 : valid_118_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3698 = 7'h77 == _GEN_13029 ? 1'h0 : valid_119_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3699 = 7'h78 == _GEN_13029 ? 1'h0 : valid_120_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3700 = 7'h79 == _GEN_13029 ? 1'h0 : valid_121_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3701 = 7'h7a == _GEN_13029 ? 1'h0 : valid_122_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3702 = 7'h7b == _GEN_13029 ? 1'h0 : valid_123_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3703 = 7'h7c == _GEN_13029 ? 1'h0 : valid_124_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3704 = 7'h7d == _GEN_13029 ? 1'h0 : valid_125_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3705 = 7'h7e == _GEN_13029 ? 1'h0 : valid_126_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3706 = 7'h7f == _GEN_13029 ? 1'h0 : valid_127_1; // @[DCache.scala 336:{39,39} 68:22]
  wire  _GEN_3707 = _GEN_3322 | _GEN_3450 ? _GEN_3451 : valid_0_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3708 = _GEN_3322 | _GEN_3450 ? _GEN_3452 : valid_1_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3709 = _GEN_3322 | _GEN_3450 ? _GEN_3453 : valid_2_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3710 = _GEN_3322 | _GEN_3450 ? _GEN_3454 : valid_3_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3711 = _GEN_3322 | _GEN_3450 ? _GEN_3455 : valid_4_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3712 = _GEN_3322 | _GEN_3450 ? _GEN_3456 : valid_5_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3713 = _GEN_3322 | _GEN_3450 ? _GEN_3457 : valid_6_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3714 = _GEN_3322 | _GEN_3450 ? _GEN_3458 : valid_7_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3715 = _GEN_3322 | _GEN_3450 ? _GEN_3459 : valid_8_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3716 = _GEN_3322 | _GEN_3450 ? _GEN_3460 : valid_9_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3717 = _GEN_3322 | _GEN_3450 ? _GEN_3461 : valid_10_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3718 = _GEN_3322 | _GEN_3450 ? _GEN_3462 : valid_11_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3719 = _GEN_3322 | _GEN_3450 ? _GEN_3463 : valid_12_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3720 = _GEN_3322 | _GEN_3450 ? _GEN_3464 : valid_13_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3721 = _GEN_3322 | _GEN_3450 ? _GEN_3465 : valid_14_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3722 = _GEN_3322 | _GEN_3450 ? _GEN_3466 : valid_15_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3723 = _GEN_3322 | _GEN_3450 ? _GEN_3467 : valid_16_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3724 = _GEN_3322 | _GEN_3450 ? _GEN_3468 : valid_17_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3725 = _GEN_3322 | _GEN_3450 ? _GEN_3469 : valid_18_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3726 = _GEN_3322 | _GEN_3450 ? _GEN_3470 : valid_19_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3727 = _GEN_3322 | _GEN_3450 ? _GEN_3471 : valid_20_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3728 = _GEN_3322 | _GEN_3450 ? _GEN_3472 : valid_21_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3729 = _GEN_3322 | _GEN_3450 ? _GEN_3473 : valid_22_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3730 = _GEN_3322 | _GEN_3450 ? _GEN_3474 : valid_23_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3731 = _GEN_3322 | _GEN_3450 ? _GEN_3475 : valid_24_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3732 = _GEN_3322 | _GEN_3450 ? _GEN_3476 : valid_25_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3733 = _GEN_3322 | _GEN_3450 ? _GEN_3477 : valid_26_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3734 = _GEN_3322 | _GEN_3450 ? _GEN_3478 : valid_27_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3735 = _GEN_3322 | _GEN_3450 ? _GEN_3479 : valid_28_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3736 = _GEN_3322 | _GEN_3450 ? _GEN_3480 : valid_29_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3737 = _GEN_3322 | _GEN_3450 ? _GEN_3481 : valid_30_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3738 = _GEN_3322 | _GEN_3450 ? _GEN_3482 : valid_31_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3739 = _GEN_3322 | _GEN_3450 ? _GEN_3483 : valid_32_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3740 = _GEN_3322 | _GEN_3450 ? _GEN_3484 : valid_33_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3741 = _GEN_3322 | _GEN_3450 ? _GEN_3485 : valid_34_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3742 = _GEN_3322 | _GEN_3450 ? _GEN_3486 : valid_35_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3743 = _GEN_3322 | _GEN_3450 ? _GEN_3487 : valid_36_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3744 = _GEN_3322 | _GEN_3450 ? _GEN_3488 : valid_37_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3745 = _GEN_3322 | _GEN_3450 ? _GEN_3489 : valid_38_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3746 = _GEN_3322 | _GEN_3450 ? _GEN_3490 : valid_39_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3747 = _GEN_3322 | _GEN_3450 ? _GEN_3491 : valid_40_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3748 = _GEN_3322 | _GEN_3450 ? _GEN_3492 : valid_41_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3749 = _GEN_3322 | _GEN_3450 ? _GEN_3493 : valid_42_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3750 = _GEN_3322 | _GEN_3450 ? _GEN_3494 : valid_43_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3751 = _GEN_3322 | _GEN_3450 ? _GEN_3495 : valid_44_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3752 = _GEN_3322 | _GEN_3450 ? _GEN_3496 : valid_45_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3753 = _GEN_3322 | _GEN_3450 ? _GEN_3497 : valid_46_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3754 = _GEN_3322 | _GEN_3450 ? _GEN_3498 : valid_47_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3755 = _GEN_3322 | _GEN_3450 ? _GEN_3499 : valid_48_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3756 = _GEN_3322 | _GEN_3450 ? _GEN_3500 : valid_49_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3757 = _GEN_3322 | _GEN_3450 ? _GEN_3501 : valid_50_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3758 = _GEN_3322 | _GEN_3450 ? _GEN_3502 : valid_51_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3759 = _GEN_3322 | _GEN_3450 ? _GEN_3503 : valid_52_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3760 = _GEN_3322 | _GEN_3450 ? _GEN_3504 : valid_53_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3761 = _GEN_3322 | _GEN_3450 ? _GEN_3505 : valid_54_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3762 = _GEN_3322 | _GEN_3450 ? _GEN_3506 : valid_55_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3763 = _GEN_3322 | _GEN_3450 ? _GEN_3507 : valid_56_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3764 = _GEN_3322 | _GEN_3450 ? _GEN_3508 : valid_57_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3765 = _GEN_3322 | _GEN_3450 ? _GEN_3509 : valid_58_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3766 = _GEN_3322 | _GEN_3450 ? _GEN_3510 : valid_59_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3767 = _GEN_3322 | _GEN_3450 ? _GEN_3511 : valid_60_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3768 = _GEN_3322 | _GEN_3450 ? _GEN_3512 : valid_61_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3769 = _GEN_3322 | _GEN_3450 ? _GEN_3513 : valid_62_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3770 = _GEN_3322 | _GEN_3450 ? _GEN_3514 : valid_63_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3771 = _GEN_3322 | _GEN_3450 ? _GEN_3515 : valid_64_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3772 = _GEN_3322 | _GEN_3450 ? _GEN_3516 : valid_65_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3773 = _GEN_3322 | _GEN_3450 ? _GEN_3517 : valid_66_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3774 = _GEN_3322 | _GEN_3450 ? _GEN_3518 : valid_67_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3775 = _GEN_3322 | _GEN_3450 ? _GEN_3519 : valid_68_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3776 = _GEN_3322 | _GEN_3450 ? _GEN_3520 : valid_69_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3777 = _GEN_3322 | _GEN_3450 ? _GEN_3521 : valid_70_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3778 = _GEN_3322 | _GEN_3450 ? _GEN_3522 : valid_71_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3779 = _GEN_3322 | _GEN_3450 ? _GEN_3523 : valid_72_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3780 = _GEN_3322 | _GEN_3450 ? _GEN_3524 : valid_73_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3781 = _GEN_3322 | _GEN_3450 ? _GEN_3525 : valid_74_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3782 = _GEN_3322 | _GEN_3450 ? _GEN_3526 : valid_75_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3783 = _GEN_3322 | _GEN_3450 ? _GEN_3527 : valid_76_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3784 = _GEN_3322 | _GEN_3450 ? _GEN_3528 : valid_77_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3785 = _GEN_3322 | _GEN_3450 ? _GEN_3529 : valid_78_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3786 = _GEN_3322 | _GEN_3450 ? _GEN_3530 : valid_79_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3787 = _GEN_3322 | _GEN_3450 ? _GEN_3531 : valid_80_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3788 = _GEN_3322 | _GEN_3450 ? _GEN_3532 : valid_81_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3789 = _GEN_3322 | _GEN_3450 ? _GEN_3533 : valid_82_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3790 = _GEN_3322 | _GEN_3450 ? _GEN_3534 : valid_83_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3791 = _GEN_3322 | _GEN_3450 ? _GEN_3535 : valid_84_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3792 = _GEN_3322 | _GEN_3450 ? _GEN_3536 : valid_85_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3793 = _GEN_3322 | _GEN_3450 ? _GEN_3537 : valid_86_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3794 = _GEN_3322 | _GEN_3450 ? _GEN_3538 : valid_87_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3795 = _GEN_3322 | _GEN_3450 ? _GEN_3539 : valid_88_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3796 = _GEN_3322 | _GEN_3450 ? _GEN_3540 : valid_89_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3797 = _GEN_3322 | _GEN_3450 ? _GEN_3541 : valid_90_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3798 = _GEN_3322 | _GEN_3450 ? _GEN_3542 : valid_91_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3799 = _GEN_3322 | _GEN_3450 ? _GEN_3543 : valid_92_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3800 = _GEN_3322 | _GEN_3450 ? _GEN_3544 : valid_93_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3801 = _GEN_3322 | _GEN_3450 ? _GEN_3545 : valid_94_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3802 = _GEN_3322 | _GEN_3450 ? _GEN_3546 : valid_95_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3803 = _GEN_3322 | _GEN_3450 ? _GEN_3547 : valid_96_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3804 = _GEN_3322 | _GEN_3450 ? _GEN_3548 : valid_97_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3805 = _GEN_3322 | _GEN_3450 ? _GEN_3549 : valid_98_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3806 = _GEN_3322 | _GEN_3450 ? _GEN_3550 : valid_99_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3807 = _GEN_3322 | _GEN_3450 ? _GEN_3551 : valid_100_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3808 = _GEN_3322 | _GEN_3450 ? _GEN_3552 : valid_101_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3809 = _GEN_3322 | _GEN_3450 ? _GEN_3553 : valid_102_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3810 = _GEN_3322 | _GEN_3450 ? _GEN_3554 : valid_103_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3811 = _GEN_3322 | _GEN_3450 ? _GEN_3555 : valid_104_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3812 = _GEN_3322 | _GEN_3450 ? _GEN_3556 : valid_105_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3813 = _GEN_3322 | _GEN_3450 ? _GEN_3557 : valid_106_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3814 = _GEN_3322 | _GEN_3450 ? _GEN_3558 : valid_107_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3815 = _GEN_3322 | _GEN_3450 ? _GEN_3559 : valid_108_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3816 = _GEN_3322 | _GEN_3450 ? _GEN_3560 : valid_109_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3817 = _GEN_3322 | _GEN_3450 ? _GEN_3561 : valid_110_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3818 = _GEN_3322 | _GEN_3450 ? _GEN_3562 : valid_111_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3819 = _GEN_3322 | _GEN_3450 ? _GEN_3563 : valid_112_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3820 = _GEN_3322 | _GEN_3450 ? _GEN_3564 : valid_113_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3821 = _GEN_3322 | _GEN_3450 ? _GEN_3565 : valid_114_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3822 = _GEN_3322 | _GEN_3450 ? _GEN_3566 : valid_115_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3823 = _GEN_3322 | _GEN_3450 ? _GEN_3567 : valid_116_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3824 = _GEN_3322 | _GEN_3450 ? _GEN_3568 : valid_117_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3825 = _GEN_3322 | _GEN_3450 ? _GEN_3569 : valid_118_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3826 = _GEN_3322 | _GEN_3450 ? _GEN_3570 : valid_119_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3827 = _GEN_3322 | _GEN_3450 ? _GEN_3571 : valid_120_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3828 = _GEN_3322 | _GEN_3450 ? _GEN_3572 : valid_121_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3829 = _GEN_3322 | _GEN_3450 ? _GEN_3573 : valid_122_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3830 = _GEN_3322 | _GEN_3450 ? _GEN_3574 : valid_123_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3831 = _GEN_3322 | _GEN_3450 ? _GEN_3575 : valid_124_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3832 = _GEN_3322 | _GEN_3450 ? _GEN_3576 : valid_125_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3833 = _GEN_3322 | _GEN_3450 ? _GEN_3577 : valid_126_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3834 = _GEN_3322 | _GEN_3450 ? _GEN_3578 : valid_127_0; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3835 = _GEN_3322 | _GEN_3450 ? _GEN_3579 : valid_0_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3836 = _GEN_3322 | _GEN_3450 ? _GEN_3580 : valid_1_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3837 = _GEN_3322 | _GEN_3450 ? _GEN_3581 : valid_2_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3838 = _GEN_3322 | _GEN_3450 ? _GEN_3582 : valid_3_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3839 = _GEN_3322 | _GEN_3450 ? _GEN_3583 : valid_4_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3840 = _GEN_3322 | _GEN_3450 ? _GEN_3584 : valid_5_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3841 = _GEN_3322 | _GEN_3450 ? _GEN_3585 : valid_6_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3842 = _GEN_3322 | _GEN_3450 ? _GEN_3586 : valid_7_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3843 = _GEN_3322 | _GEN_3450 ? _GEN_3587 : valid_8_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3844 = _GEN_3322 | _GEN_3450 ? _GEN_3588 : valid_9_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3845 = _GEN_3322 | _GEN_3450 ? _GEN_3589 : valid_10_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3846 = _GEN_3322 | _GEN_3450 ? _GEN_3590 : valid_11_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3847 = _GEN_3322 | _GEN_3450 ? _GEN_3591 : valid_12_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3848 = _GEN_3322 | _GEN_3450 ? _GEN_3592 : valid_13_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3849 = _GEN_3322 | _GEN_3450 ? _GEN_3593 : valid_14_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3850 = _GEN_3322 | _GEN_3450 ? _GEN_3594 : valid_15_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3851 = _GEN_3322 | _GEN_3450 ? _GEN_3595 : valid_16_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3852 = _GEN_3322 | _GEN_3450 ? _GEN_3596 : valid_17_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3853 = _GEN_3322 | _GEN_3450 ? _GEN_3597 : valid_18_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3854 = _GEN_3322 | _GEN_3450 ? _GEN_3598 : valid_19_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3855 = _GEN_3322 | _GEN_3450 ? _GEN_3599 : valid_20_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3856 = _GEN_3322 | _GEN_3450 ? _GEN_3600 : valid_21_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3857 = _GEN_3322 | _GEN_3450 ? _GEN_3601 : valid_22_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3858 = _GEN_3322 | _GEN_3450 ? _GEN_3602 : valid_23_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3859 = _GEN_3322 | _GEN_3450 ? _GEN_3603 : valid_24_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3860 = _GEN_3322 | _GEN_3450 ? _GEN_3604 : valid_25_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3861 = _GEN_3322 | _GEN_3450 ? _GEN_3605 : valid_26_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3862 = _GEN_3322 | _GEN_3450 ? _GEN_3606 : valid_27_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3863 = _GEN_3322 | _GEN_3450 ? _GEN_3607 : valid_28_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3864 = _GEN_3322 | _GEN_3450 ? _GEN_3608 : valid_29_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3865 = _GEN_3322 | _GEN_3450 ? _GEN_3609 : valid_30_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3866 = _GEN_3322 | _GEN_3450 ? _GEN_3610 : valid_31_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3867 = _GEN_3322 | _GEN_3450 ? _GEN_3611 : valid_32_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3868 = _GEN_3322 | _GEN_3450 ? _GEN_3612 : valid_33_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3869 = _GEN_3322 | _GEN_3450 ? _GEN_3613 : valid_34_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3870 = _GEN_3322 | _GEN_3450 ? _GEN_3614 : valid_35_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3871 = _GEN_3322 | _GEN_3450 ? _GEN_3615 : valid_36_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3872 = _GEN_3322 | _GEN_3450 ? _GEN_3616 : valid_37_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3873 = _GEN_3322 | _GEN_3450 ? _GEN_3617 : valid_38_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3874 = _GEN_3322 | _GEN_3450 ? _GEN_3618 : valid_39_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3875 = _GEN_3322 | _GEN_3450 ? _GEN_3619 : valid_40_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3876 = _GEN_3322 | _GEN_3450 ? _GEN_3620 : valid_41_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3877 = _GEN_3322 | _GEN_3450 ? _GEN_3621 : valid_42_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3878 = _GEN_3322 | _GEN_3450 ? _GEN_3622 : valid_43_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3879 = _GEN_3322 | _GEN_3450 ? _GEN_3623 : valid_44_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3880 = _GEN_3322 | _GEN_3450 ? _GEN_3624 : valid_45_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3881 = _GEN_3322 | _GEN_3450 ? _GEN_3625 : valid_46_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3882 = _GEN_3322 | _GEN_3450 ? _GEN_3626 : valid_47_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3883 = _GEN_3322 | _GEN_3450 ? _GEN_3627 : valid_48_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3884 = _GEN_3322 | _GEN_3450 ? _GEN_3628 : valid_49_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3885 = _GEN_3322 | _GEN_3450 ? _GEN_3629 : valid_50_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3886 = _GEN_3322 | _GEN_3450 ? _GEN_3630 : valid_51_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3887 = _GEN_3322 | _GEN_3450 ? _GEN_3631 : valid_52_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3888 = _GEN_3322 | _GEN_3450 ? _GEN_3632 : valid_53_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3889 = _GEN_3322 | _GEN_3450 ? _GEN_3633 : valid_54_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3890 = _GEN_3322 | _GEN_3450 ? _GEN_3634 : valid_55_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3891 = _GEN_3322 | _GEN_3450 ? _GEN_3635 : valid_56_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3892 = _GEN_3322 | _GEN_3450 ? _GEN_3636 : valid_57_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3893 = _GEN_3322 | _GEN_3450 ? _GEN_3637 : valid_58_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3894 = _GEN_3322 | _GEN_3450 ? _GEN_3638 : valid_59_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3895 = _GEN_3322 | _GEN_3450 ? _GEN_3639 : valid_60_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3896 = _GEN_3322 | _GEN_3450 ? _GEN_3640 : valid_61_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3897 = _GEN_3322 | _GEN_3450 ? _GEN_3641 : valid_62_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3898 = _GEN_3322 | _GEN_3450 ? _GEN_3642 : valid_63_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3899 = _GEN_3322 | _GEN_3450 ? _GEN_3643 : valid_64_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3900 = _GEN_3322 | _GEN_3450 ? _GEN_3644 : valid_65_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3901 = _GEN_3322 | _GEN_3450 ? _GEN_3645 : valid_66_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3902 = _GEN_3322 | _GEN_3450 ? _GEN_3646 : valid_67_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3903 = _GEN_3322 | _GEN_3450 ? _GEN_3647 : valid_68_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3904 = _GEN_3322 | _GEN_3450 ? _GEN_3648 : valid_69_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3905 = _GEN_3322 | _GEN_3450 ? _GEN_3649 : valid_70_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3906 = _GEN_3322 | _GEN_3450 ? _GEN_3650 : valid_71_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3907 = _GEN_3322 | _GEN_3450 ? _GEN_3651 : valid_72_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3908 = _GEN_3322 | _GEN_3450 ? _GEN_3652 : valid_73_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3909 = _GEN_3322 | _GEN_3450 ? _GEN_3653 : valid_74_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3910 = _GEN_3322 | _GEN_3450 ? _GEN_3654 : valid_75_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3911 = _GEN_3322 | _GEN_3450 ? _GEN_3655 : valid_76_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3912 = _GEN_3322 | _GEN_3450 ? _GEN_3656 : valid_77_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3913 = _GEN_3322 | _GEN_3450 ? _GEN_3657 : valid_78_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3914 = _GEN_3322 | _GEN_3450 ? _GEN_3658 : valid_79_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3915 = _GEN_3322 | _GEN_3450 ? _GEN_3659 : valid_80_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3916 = _GEN_3322 | _GEN_3450 ? _GEN_3660 : valid_81_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3917 = _GEN_3322 | _GEN_3450 ? _GEN_3661 : valid_82_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3918 = _GEN_3322 | _GEN_3450 ? _GEN_3662 : valid_83_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3919 = _GEN_3322 | _GEN_3450 ? _GEN_3663 : valid_84_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3920 = _GEN_3322 | _GEN_3450 ? _GEN_3664 : valid_85_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3921 = _GEN_3322 | _GEN_3450 ? _GEN_3665 : valid_86_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3922 = _GEN_3322 | _GEN_3450 ? _GEN_3666 : valid_87_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3923 = _GEN_3322 | _GEN_3450 ? _GEN_3667 : valid_88_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3924 = _GEN_3322 | _GEN_3450 ? _GEN_3668 : valid_89_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3925 = _GEN_3322 | _GEN_3450 ? _GEN_3669 : valid_90_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3926 = _GEN_3322 | _GEN_3450 ? _GEN_3670 : valid_91_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3927 = _GEN_3322 | _GEN_3450 ? _GEN_3671 : valid_92_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3928 = _GEN_3322 | _GEN_3450 ? _GEN_3672 : valid_93_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3929 = _GEN_3322 | _GEN_3450 ? _GEN_3673 : valid_94_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3930 = _GEN_3322 | _GEN_3450 ? _GEN_3674 : valid_95_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3931 = _GEN_3322 | _GEN_3450 ? _GEN_3675 : valid_96_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3932 = _GEN_3322 | _GEN_3450 ? _GEN_3676 : valid_97_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3933 = _GEN_3322 | _GEN_3450 ? _GEN_3677 : valid_98_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3934 = _GEN_3322 | _GEN_3450 ? _GEN_3678 : valid_99_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3935 = _GEN_3322 | _GEN_3450 ? _GEN_3679 : valid_100_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3936 = _GEN_3322 | _GEN_3450 ? _GEN_3680 : valid_101_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3937 = _GEN_3322 | _GEN_3450 ? _GEN_3681 : valid_102_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3938 = _GEN_3322 | _GEN_3450 ? _GEN_3682 : valid_103_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3939 = _GEN_3322 | _GEN_3450 ? _GEN_3683 : valid_104_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3940 = _GEN_3322 | _GEN_3450 ? _GEN_3684 : valid_105_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3941 = _GEN_3322 | _GEN_3450 ? _GEN_3685 : valid_106_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3942 = _GEN_3322 | _GEN_3450 ? _GEN_3686 : valid_107_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3943 = _GEN_3322 | _GEN_3450 ? _GEN_3687 : valid_108_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3944 = _GEN_3322 | _GEN_3450 ? _GEN_3688 : valid_109_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3945 = _GEN_3322 | _GEN_3450 ? _GEN_3689 : valid_110_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3946 = _GEN_3322 | _GEN_3450 ? _GEN_3690 : valid_111_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3947 = _GEN_3322 | _GEN_3450 ? _GEN_3691 : valid_112_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3948 = _GEN_3322 | _GEN_3450 ? _GEN_3692 : valid_113_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3949 = _GEN_3322 | _GEN_3450 ? _GEN_3693 : valid_114_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3950 = _GEN_3322 | _GEN_3450 ? _GEN_3694 : valid_115_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3951 = _GEN_3322 | _GEN_3450 ? _GEN_3695 : valid_116_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3952 = _GEN_3322 | _GEN_3450 ? _GEN_3696 : valid_117_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3953 = _GEN_3322 | _GEN_3450 ? _GEN_3697 : valid_118_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3954 = _GEN_3322 | _GEN_3450 ? _GEN_3698 : valid_119_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3955 = _GEN_3322 | _GEN_3450 ? _GEN_3699 : valid_120_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3956 = _GEN_3322 | _GEN_3450 ? _GEN_3700 : valid_121_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3957 = _GEN_3322 | _GEN_3450 ? _GEN_3701 : valid_122_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3958 = _GEN_3322 | _GEN_3450 ? _GEN_3702 : valid_123_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3959 = _GEN_3322 | _GEN_3450 ? _GEN_3703 : valid_124_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3960 = _GEN_3322 | _GEN_3450 ? _GEN_3704 : valid_125_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3961 = _GEN_3322 | _GEN_3450 ? _GEN_3705 : valid_126_1; // @[DCache.scala 334:57 68:22]
  wire  _GEN_3962 = _GEN_3322 | _GEN_3450 ? _GEN_3706 : valid_127_1; // @[DCache.scala 334:57 68:22]
  wire [2:0] _GEN_3963 = _GEN_3059 | _GEN_3187 ? _GEN_3188 : 3'h5; // @[DCache.scala 323:55 338:17]
  wire [3:0] _GEN_3964 = _GEN_3059 | _GEN_3187 ? _GEN_3189 : axi_wcnt; // @[DCache.scala 323:55 89:40]
  wire [9:0] _GEN_3965 = _GEN_3059 | _GEN_3187 ? _GEN_3190 : bram_replace_addr; // @[DCache.scala 323:55 90:40]
  wire [9:0] _GEN_3966 = _GEN_3059 | _GEN_3187 ? _GEN_3191 : bram_read_ready_addr; // @[DCache.scala 323:55 91:40]
  wire  _GEN_3968 = _GEN_3059 | _GEN_3187 ? _GEN_3193 : bram_use_replace_addr; // @[DCache.scala 323:55 95:40]
  wire  _GEN_3970 = _GEN_3059 | _GEN_3187 ? valid_0_0 : _GEN_3707; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3971 = _GEN_3059 | _GEN_3187 ? valid_1_0 : _GEN_3708; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3972 = _GEN_3059 | _GEN_3187 ? valid_2_0 : _GEN_3709; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3973 = _GEN_3059 | _GEN_3187 ? valid_3_0 : _GEN_3710; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3974 = _GEN_3059 | _GEN_3187 ? valid_4_0 : _GEN_3711; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3975 = _GEN_3059 | _GEN_3187 ? valid_5_0 : _GEN_3712; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3976 = _GEN_3059 | _GEN_3187 ? valid_6_0 : _GEN_3713; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3977 = _GEN_3059 | _GEN_3187 ? valid_7_0 : _GEN_3714; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3978 = _GEN_3059 | _GEN_3187 ? valid_8_0 : _GEN_3715; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3979 = _GEN_3059 | _GEN_3187 ? valid_9_0 : _GEN_3716; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3980 = _GEN_3059 | _GEN_3187 ? valid_10_0 : _GEN_3717; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3981 = _GEN_3059 | _GEN_3187 ? valid_11_0 : _GEN_3718; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3982 = _GEN_3059 | _GEN_3187 ? valid_12_0 : _GEN_3719; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3983 = _GEN_3059 | _GEN_3187 ? valid_13_0 : _GEN_3720; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3984 = _GEN_3059 | _GEN_3187 ? valid_14_0 : _GEN_3721; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3985 = _GEN_3059 | _GEN_3187 ? valid_15_0 : _GEN_3722; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3986 = _GEN_3059 | _GEN_3187 ? valid_16_0 : _GEN_3723; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3987 = _GEN_3059 | _GEN_3187 ? valid_17_0 : _GEN_3724; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3988 = _GEN_3059 | _GEN_3187 ? valid_18_0 : _GEN_3725; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3989 = _GEN_3059 | _GEN_3187 ? valid_19_0 : _GEN_3726; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3990 = _GEN_3059 | _GEN_3187 ? valid_20_0 : _GEN_3727; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3991 = _GEN_3059 | _GEN_3187 ? valid_21_0 : _GEN_3728; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3992 = _GEN_3059 | _GEN_3187 ? valid_22_0 : _GEN_3729; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3993 = _GEN_3059 | _GEN_3187 ? valid_23_0 : _GEN_3730; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3994 = _GEN_3059 | _GEN_3187 ? valid_24_0 : _GEN_3731; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3995 = _GEN_3059 | _GEN_3187 ? valid_25_0 : _GEN_3732; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3996 = _GEN_3059 | _GEN_3187 ? valid_26_0 : _GEN_3733; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3997 = _GEN_3059 | _GEN_3187 ? valid_27_0 : _GEN_3734; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3998 = _GEN_3059 | _GEN_3187 ? valid_28_0 : _GEN_3735; // @[DCache.scala 323:55 68:22]
  wire  _GEN_3999 = _GEN_3059 | _GEN_3187 ? valid_29_0 : _GEN_3736; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4000 = _GEN_3059 | _GEN_3187 ? valid_30_0 : _GEN_3737; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4001 = _GEN_3059 | _GEN_3187 ? valid_31_0 : _GEN_3738; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4002 = _GEN_3059 | _GEN_3187 ? valid_32_0 : _GEN_3739; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4003 = _GEN_3059 | _GEN_3187 ? valid_33_0 : _GEN_3740; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4004 = _GEN_3059 | _GEN_3187 ? valid_34_0 : _GEN_3741; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4005 = _GEN_3059 | _GEN_3187 ? valid_35_0 : _GEN_3742; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4006 = _GEN_3059 | _GEN_3187 ? valid_36_0 : _GEN_3743; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4007 = _GEN_3059 | _GEN_3187 ? valid_37_0 : _GEN_3744; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4008 = _GEN_3059 | _GEN_3187 ? valid_38_0 : _GEN_3745; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4009 = _GEN_3059 | _GEN_3187 ? valid_39_0 : _GEN_3746; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4010 = _GEN_3059 | _GEN_3187 ? valid_40_0 : _GEN_3747; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4011 = _GEN_3059 | _GEN_3187 ? valid_41_0 : _GEN_3748; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4012 = _GEN_3059 | _GEN_3187 ? valid_42_0 : _GEN_3749; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4013 = _GEN_3059 | _GEN_3187 ? valid_43_0 : _GEN_3750; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4014 = _GEN_3059 | _GEN_3187 ? valid_44_0 : _GEN_3751; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4015 = _GEN_3059 | _GEN_3187 ? valid_45_0 : _GEN_3752; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4016 = _GEN_3059 | _GEN_3187 ? valid_46_0 : _GEN_3753; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4017 = _GEN_3059 | _GEN_3187 ? valid_47_0 : _GEN_3754; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4018 = _GEN_3059 | _GEN_3187 ? valid_48_0 : _GEN_3755; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4019 = _GEN_3059 | _GEN_3187 ? valid_49_0 : _GEN_3756; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4020 = _GEN_3059 | _GEN_3187 ? valid_50_0 : _GEN_3757; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4021 = _GEN_3059 | _GEN_3187 ? valid_51_0 : _GEN_3758; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4022 = _GEN_3059 | _GEN_3187 ? valid_52_0 : _GEN_3759; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4023 = _GEN_3059 | _GEN_3187 ? valid_53_0 : _GEN_3760; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4024 = _GEN_3059 | _GEN_3187 ? valid_54_0 : _GEN_3761; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4025 = _GEN_3059 | _GEN_3187 ? valid_55_0 : _GEN_3762; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4026 = _GEN_3059 | _GEN_3187 ? valid_56_0 : _GEN_3763; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4027 = _GEN_3059 | _GEN_3187 ? valid_57_0 : _GEN_3764; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4028 = _GEN_3059 | _GEN_3187 ? valid_58_0 : _GEN_3765; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4029 = _GEN_3059 | _GEN_3187 ? valid_59_0 : _GEN_3766; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4030 = _GEN_3059 | _GEN_3187 ? valid_60_0 : _GEN_3767; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4031 = _GEN_3059 | _GEN_3187 ? valid_61_0 : _GEN_3768; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4032 = _GEN_3059 | _GEN_3187 ? valid_62_0 : _GEN_3769; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4033 = _GEN_3059 | _GEN_3187 ? valid_63_0 : _GEN_3770; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4034 = _GEN_3059 | _GEN_3187 ? valid_64_0 : _GEN_3771; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4035 = _GEN_3059 | _GEN_3187 ? valid_65_0 : _GEN_3772; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4036 = _GEN_3059 | _GEN_3187 ? valid_66_0 : _GEN_3773; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4037 = _GEN_3059 | _GEN_3187 ? valid_67_0 : _GEN_3774; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4038 = _GEN_3059 | _GEN_3187 ? valid_68_0 : _GEN_3775; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4039 = _GEN_3059 | _GEN_3187 ? valid_69_0 : _GEN_3776; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4040 = _GEN_3059 | _GEN_3187 ? valid_70_0 : _GEN_3777; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4041 = _GEN_3059 | _GEN_3187 ? valid_71_0 : _GEN_3778; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4042 = _GEN_3059 | _GEN_3187 ? valid_72_0 : _GEN_3779; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4043 = _GEN_3059 | _GEN_3187 ? valid_73_0 : _GEN_3780; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4044 = _GEN_3059 | _GEN_3187 ? valid_74_0 : _GEN_3781; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4045 = _GEN_3059 | _GEN_3187 ? valid_75_0 : _GEN_3782; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4046 = _GEN_3059 | _GEN_3187 ? valid_76_0 : _GEN_3783; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4047 = _GEN_3059 | _GEN_3187 ? valid_77_0 : _GEN_3784; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4048 = _GEN_3059 | _GEN_3187 ? valid_78_0 : _GEN_3785; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4049 = _GEN_3059 | _GEN_3187 ? valid_79_0 : _GEN_3786; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4050 = _GEN_3059 | _GEN_3187 ? valid_80_0 : _GEN_3787; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4051 = _GEN_3059 | _GEN_3187 ? valid_81_0 : _GEN_3788; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4052 = _GEN_3059 | _GEN_3187 ? valid_82_0 : _GEN_3789; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4053 = _GEN_3059 | _GEN_3187 ? valid_83_0 : _GEN_3790; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4054 = _GEN_3059 | _GEN_3187 ? valid_84_0 : _GEN_3791; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4055 = _GEN_3059 | _GEN_3187 ? valid_85_0 : _GEN_3792; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4056 = _GEN_3059 | _GEN_3187 ? valid_86_0 : _GEN_3793; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4057 = _GEN_3059 | _GEN_3187 ? valid_87_0 : _GEN_3794; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4058 = _GEN_3059 | _GEN_3187 ? valid_88_0 : _GEN_3795; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4059 = _GEN_3059 | _GEN_3187 ? valid_89_0 : _GEN_3796; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4060 = _GEN_3059 | _GEN_3187 ? valid_90_0 : _GEN_3797; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4061 = _GEN_3059 | _GEN_3187 ? valid_91_0 : _GEN_3798; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4062 = _GEN_3059 | _GEN_3187 ? valid_92_0 : _GEN_3799; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4063 = _GEN_3059 | _GEN_3187 ? valid_93_0 : _GEN_3800; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4064 = _GEN_3059 | _GEN_3187 ? valid_94_0 : _GEN_3801; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4065 = _GEN_3059 | _GEN_3187 ? valid_95_0 : _GEN_3802; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4066 = _GEN_3059 | _GEN_3187 ? valid_96_0 : _GEN_3803; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4067 = _GEN_3059 | _GEN_3187 ? valid_97_0 : _GEN_3804; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4068 = _GEN_3059 | _GEN_3187 ? valid_98_0 : _GEN_3805; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4069 = _GEN_3059 | _GEN_3187 ? valid_99_0 : _GEN_3806; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4070 = _GEN_3059 | _GEN_3187 ? valid_100_0 : _GEN_3807; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4071 = _GEN_3059 | _GEN_3187 ? valid_101_0 : _GEN_3808; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4072 = _GEN_3059 | _GEN_3187 ? valid_102_0 : _GEN_3809; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4073 = _GEN_3059 | _GEN_3187 ? valid_103_0 : _GEN_3810; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4074 = _GEN_3059 | _GEN_3187 ? valid_104_0 : _GEN_3811; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4075 = _GEN_3059 | _GEN_3187 ? valid_105_0 : _GEN_3812; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4076 = _GEN_3059 | _GEN_3187 ? valid_106_0 : _GEN_3813; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4077 = _GEN_3059 | _GEN_3187 ? valid_107_0 : _GEN_3814; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4078 = _GEN_3059 | _GEN_3187 ? valid_108_0 : _GEN_3815; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4079 = _GEN_3059 | _GEN_3187 ? valid_109_0 : _GEN_3816; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4080 = _GEN_3059 | _GEN_3187 ? valid_110_0 : _GEN_3817; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4081 = _GEN_3059 | _GEN_3187 ? valid_111_0 : _GEN_3818; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4082 = _GEN_3059 | _GEN_3187 ? valid_112_0 : _GEN_3819; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4083 = _GEN_3059 | _GEN_3187 ? valid_113_0 : _GEN_3820; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4084 = _GEN_3059 | _GEN_3187 ? valid_114_0 : _GEN_3821; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4085 = _GEN_3059 | _GEN_3187 ? valid_115_0 : _GEN_3822; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4086 = _GEN_3059 | _GEN_3187 ? valid_116_0 : _GEN_3823; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4087 = _GEN_3059 | _GEN_3187 ? valid_117_0 : _GEN_3824; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4088 = _GEN_3059 | _GEN_3187 ? valid_118_0 : _GEN_3825; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4089 = _GEN_3059 | _GEN_3187 ? valid_119_0 : _GEN_3826; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4090 = _GEN_3059 | _GEN_3187 ? valid_120_0 : _GEN_3827; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4091 = _GEN_3059 | _GEN_3187 ? valid_121_0 : _GEN_3828; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4092 = _GEN_3059 | _GEN_3187 ? valid_122_0 : _GEN_3829; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4093 = _GEN_3059 | _GEN_3187 ? valid_123_0 : _GEN_3830; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4094 = _GEN_3059 | _GEN_3187 ? valid_124_0 : _GEN_3831; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4095 = _GEN_3059 | _GEN_3187 ? valid_125_0 : _GEN_3832; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4096 = _GEN_3059 | _GEN_3187 ? valid_126_0 : _GEN_3833; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4097 = _GEN_3059 | _GEN_3187 ? valid_127_0 : _GEN_3834; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4098 = _GEN_3059 | _GEN_3187 ? valid_0_1 : _GEN_3835; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4099 = _GEN_3059 | _GEN_3187 ? valid_1_1 : _GEN_3836; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4100 = _GEN_3059 | _GEN_3187 ? valid_2_1 : _GEN_3837; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4101 = _GEN_3059 | _GEN_3187 ? valid_3_1 : _GEN_3838; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4102 = _GEN_3059 | _GEN_3187 ? valid_4_1 : _GEN_3839; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4103 = _GEN_3059 | _GEN_3187 ? valid_5_1 : _GEN_3840; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4104 = _GEN_3059 | _GEN_3187 ? valid_6_1 : _GEN_3841; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4105 = _GEN_3059 | _GEN_3187 ? valid_7_1 : _GEN_3842; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4106 = _GEN_3059 | _GEN_3187 ? valid_8_1 : _GEN_3843; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4107 = _GEN_3059 | _GEN_3187 ? valid_9_1 : _GEN_3844; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4108 = _GEN_3059 | _GEN_3187 ? valid_10_1 : _GEN_3845; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4109 = _GEN_3059 | _GEN_3187 ? valid_11_1 : _GEN_3846; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4110 = _GEN_3059 | _GEN_3187 ? valid_12_1 : _GEN_3847; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4111 = _GEN_3059 | _GEN_3187 ? valid_13_1 : _GEN_3848; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4112 = _GEN_3059 | _GEN_3187 ? valid_14_1 : _GEN_3849; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4113 = _GEN_3059 | _GEN_3187 ? valid_15_1 : _GEN_3850; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4114 = _GEN_3059 | _GEN_3187 ? valid_16_1 : _GEN_3851; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4115 = _GEN_3059 | _GEN_3187 ? valid_17_1 : _GEN_3852; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4116 = _GEN_3059 | _GEN_3187 ? valid_18_1 : _GEN_3853; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4117 = _GEN_3059 | _GEN_3187 ? valid_19_1 : _GEN_3854; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4118 = _GEN_3059 | _GEN_3187 ? valid_20_1 : _GEN_3855; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4119 = _GEN_3059 | _GEN_3187 ? valid_21_1 : _GEN_3856; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4120 = _GEN_3059 | _GEN_3187 ? valid_22_1 : _GEN_3857; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4121 = _GEN_3059 | _GEN_3187 ? valid_23_1 : _GEN_3858; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4122 = _GEN_3059 | _GEN_3187 ? valid_24_1 : _GEN_3859; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4123 = _GEN_3059 | _GEN_3187 ? valid_25_1 : _GEN_3860; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4124 = _GEN_3059 | _GEN_3187 ? valid_26_1 : _GEN_3861; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4125 = _GEN_3059 | _GEN_3187 ? valid_27_1 : _GEN_3862; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4126 = _GEN_3059 | _GEN_3187 ? valid_28_1 : _GEN_3863; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4127 = _GEN_3059 | _GEN_3187 ? valid_29_1 : _GEN_3864; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4128 = _GEN_3059 | _GEN_3187 ? valid_30_1 : _GEN_3865; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4129 = _GEN_3059 | _GEN_3187 ? valid_31_1 : _GEN_3866; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4130 = _GEN_3059 | _GEN_3187 ? valid_32_1 : _GEN_3867; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4131 = _GEN_3059 | _GEN_3187 ? valid_33_1 : _GEN_3868; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4132 = _GEN_3059 | _GEN_3187 ? valid_34_1 : _GEN_3869; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4133 = _GEN_3059 | _GEN_3187 ? valid_35_1 : _GEN_3870; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4134 = _GEN_3059 | _GEN_3187 ? valid_36_1 : _GEN_3871; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4135 = _GEN_3059 | _GEN_3187 ? valid_37_1 : _GEN_3872; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4136 = _GEN_3059 | _GEN_3187 ? valid_38_1 : _GEN_3873; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4137 = _GEN_3059 | _GEN_3187 ? valid_39_1 : _GEN_3874; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4138 = _GEN_3059 | _GEN_3187 ? valid_40_1 : _GEN_3875; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4139 = _GEN_3059 | _GEN_3187 ? valid_41_1 : _GEN_3876; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4140 = _GEN_3059 | _GEN_3187 ? valid_42_1 : _GEN_3877; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4141 = _GEN_3059 | _GEN_3187 ? valid_43_1 : _GEN_3878; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4142 = _GEN_3059 | _GEN_3187 ? valid_44_1 : _GEN_3879; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4143 = _GEN_3059 | _GEN_3187 ? valid_45_1 : _GEN_3880; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4144 = _GEN_3059 | _GEN_3187 ? valid_46_1 : _GEN_3881; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4145 = _GEN_3059 | _GEN_3187 ? valid_47_1 : _GEN_3882; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4146 = _GEN_3059 | _GEN_3187 ? valid_48_1 : _GEN_3883; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4147 = _GEN_3059 | _GEN_3187 ? valid_49_1 : _GEN_3884; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4148 = _GEN_3059 | _GEN_3187 ? valid_50_1 : _GEN_3885; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4149 = _GEN_3059 | _GEN_3187 ? valid_51_1 : _GEN_3886; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4150 = _GEN_3059 | _GEN_3187 ? valid_52_1 : _GEN_3887; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4151 = _GEN_3059 | _GEN_3187 ? valid_53_1 : _GEN_3888; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4152 = _GEN_3059 | _GEN_3187 ? valid_54_1 : _GEN_3889; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4153 = _GEN_3059 | _GEN_3187 ? valid_55_1 : _GEN_3890; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4154 = _GEN_3059 | _GEN_3187 ? valid_56_1 : _GEN_3891; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4155 = _GEN_3059 | _GEN_3187 ? valid_57_1 : _GEN_3892; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4156 = _GEN_3059 | _GEN_3187 ? valid_58_1 : _GEN_3893; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4157 = _GEN_3059 | _GEN_3187 ? valid_59_1 : _GEN_3894; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4158 = _GEN_3059 | _GEN_3187 ? valid_60_1 : _GEN_3895; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4159 = _GEN_3059 | _GEN_3187 ? valid_61_1 : _GEN_3896; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4160 = _GEN_3059 | _GEN_3187 ? valid_62_1 : _GEN_3897; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4161 = _GEN_3059 | _GEN_3187 ? valid_63_1 : _GEN_3898; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4162 = _GEN_3059 | _GEN_3187 ? valid_64_1 : _GEN_3899; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4163 = _GEN_3059 | _GEN_3187 ? valid_65_1 : _GEN_3900; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4164 = _GEN_3059 | _GEN_3187 ? valid_66_1 : _GEN_3901; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4165 = _GEN_3059 | _GEN_3187 ? valid_67_1 : _GEN_3902; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4166 = _GEN_3059 | _GEN_3187 ? valid_68_1 : _GEN_3903; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4167 = _GEN_3059 | _GEN_3187 ? valid_69_1 : _GEN_3904; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4168 = _GEN_3059 | _GEN_3187 ? valid_70_1 : _GEN_3905; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4169 = _GEN_3059 | _GEN_3187 ? valid_71_1 : _GEN_3906; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4170 = _GEN_3059 | _GEN_3187 ? valid_72_1 : _GEN_3907; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4171 = _GEN_3059 | _GEN_3187 ? valid_73_1 : _GEN_3908; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4172 = _GEN_3059 | _GEN_3187 ? valid_74_1 : _GEN_3909; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4173 = _GEN_3059 | _GEN_3187 ? valid_75_1 : _GEN_3910; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4174 = _GEN_3059 | _GEN_3187 ? valid_76_1 : _GEN_3911; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4175 = _GEN_3059 | _GEN_3187 ? valid_77_1 : _GEN_3912; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4176 = _GEN_3059 | _GEN_3187 ? valid_78_1 : _GEN_3913; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4177 = _GEN_3059 | _GEN_3187 ? valid_79_1 : _GEN_3914; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4178 = _GEN_3059 | _GEN_3187 ? valid_80_1 : _GEN_3915; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4179 = _GEN_3059 | _GEN_3187 ? valid_81_1 : _GEN_3916; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4180 = _GEN_3059 | _GEN_3187 ? valid_82_1 : _GEN_3917; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4181 = _GEN_3059 | _GEN_3187 ? valid_83_1 : _GEN_3918; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4182 = _GEN_3059 | _GEN_3187 ? valid_84_1 : _GEN_3919; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4183 = _GEN_3059 | _GEN_3187 ? valid_85_1 : _GEN_3920; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4184 = _GEN_3059 | _GEN_3187 ? valid_86_1 : _GEN_3921; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4185 = _GEN_3059 | _GEN_3187 ? valid_87_1 : _GEN_3922; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4186 = _GEN_3059 | _GEN_3187 ? valid_88_1 : _GEN_3923; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4187 = _GEN_3059 | _GEN_3187 ? valid_89_1 : _GEN_3924; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4188 = _GEN_3059 | _GEN_3187 ? valid_90_1 : _GEN_3925; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4189 = _GEN_3059 | _GEN_3187 ? valid_91_1 : _GEN_3926; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4190 = _GEN_3059 | _GEN_3187 ? valid_92_1 : _GEN_3927; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4191 = _GEN_3059 | _GEN_3187 ? valid_93_1 : _GEN_3928; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4192 = _GEN_3059 | _GEN_3187 ? valid_94_1 : _GEN_3929; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4193 = _GEN_3059 | _GEN_3187 ? valid_95_1 : _GEN_3930; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4194 = _GEN_3059 | _GEN_3187 ? valid_96_1 : _GEN_3931; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4195 = _GEN_3059 | _GEN_3187 ? valid_97_1 : _GEN_3932; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4196 = _GEN_3059 | _GEN_3187 ? valid_98_1 : _GEN_3933; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4197 = _GEN_3059 | _GEN_3187 ? valid_99_1 : _GEN_3934; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4198 = _GEN_3059 | _GEN_3187 ? valid_100_1 : _GEN_3935; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4199 = _GEN_3059 | _GEN_3187 ? valid_101_1 : _GEN_3936; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4200 = _GEN_3059 | _GEN_3187 ? valid_102_1 : _GEN_3937; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4201 = _GEN_3059 | _GEN_3187 ? valid_103_1 : _GEN_3938; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4202 = _GEN_3059 | _GEN_3187 ? valid_104_1 : _GEN_3939; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4203 = _GEN_3059 | _GEN_3187 ? valid_105_1 : _GEN_3940; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4204 = _GEN_3059 | _GEN_3187 ? valid_106_1 : _GEN_3941; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4205 = _GEN_3059 | _GEN_3187 ? valid_107_1 : _GEN_3942; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4206 = _GEN_3059 | _GEN_3187 ? valid_108_1 : _GEN_3943; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4207 = _GEN_3059 | _GEN_3187 ? valid_109_1 : _GEN_3944; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4208 = _GEN_3059 | _GEN_3187 ? valid_110_1 : _GEN_3945; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4209 = _GEN_3059 | _GEN_3187 ? valid_111_1 : _GEN_3946; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4210 = _GEN_3059 | _GEN_3187 ? valid_112_1 : _GEN_3947; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4211 = _GEN_3059 | _GEN_3187 ? valid_113_1 : _GEN_3948; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4212 = _GEN_3059 | _GEN_3187 ? valid_114_1 : _GEN_3949; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4213 = _GEN_3059 | _GEN_3187 ? valid_115_1 : _GEN_3950; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4214 = _GEN_3059 | _GEN_3187 ? valid_116_1 : _GEN_3951; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4215 = _GEN_3059 | _GEN_3187 ? valid_117_1 : _GEN_3952; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4216 = _GEN_3059 | _GEN_3187 ? valid_118_1 : _GEN_3953; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4217 = _GEN_3059 | _GEN_3187 ? valid_119_1 : _GEN_3954; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4218 = _GEN_3059 | _GEN_3187 ? valid_120_1 : _GEN_3955; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4219 = _GEN_3059 | _GEN_3187 ? valid_121_1 : _GEN_3956; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4220 = _GEN_3059 | _GEN_3187 ? valid_122_1 : _GEN_3957; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4221 = _GEN_3059 | _GEN_3187 ? valid_123_1 : _GEN_3958; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4222 = _GEN_3059 | _GEN_3187 ? valid_124_1 : _GEN_3959; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4223 = _GEN_3059 | _GEN_3187 ? valid_125_1 : _GEN_3960; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4224 = _GEN_3059 | _GEN_3187 ? valid_126_1 : _GEN_3961; // @[DCache.scala 323:55 68:22]
  wire  _GEN_4225 = _GEN_3059 | _GEN_3187 ? valid_127_1 : _GEN_3962; // @[DCache.scala 323:55 68:22]
  wire [19:0] _GEN_4491 = io_cpu_M_mem_en ? _GEN_2527 : {{1'd0}, tlb2_vpn}; // @[DCache.scala 245:21 262:22]
  wire  _GEN_4492 = io_cpu_M_mem_en & _GEN_2528; // @[DCache.scala 262:22 83:29]
  wire [31:0] _GEN_4493 = io_cpu_M_mem_en ? _GEN_2529 : 32'h0; // @[DCache.scala 262:22 84:29]
  wire [1:0] _GEN_4494 = io_cpu_M_mem_en ? _GEN_2530 : 2'h0; // @[DCache.scala 262:22 84:29]
  wire [3:0] _GEN_4495 = io_cpu_M_mem_en ? _GEN_2531 : 4'h0; // @[DCache.scala 262:22 84:29]
  wire [31:0] _GEN_4496 = io_cpu_M_mem_en ? _GEN_2532 : 32'h0; // @[DCache.scala 262:22 84:29]
  wire [19:0] _GEN_5153 = data_vpn[0] ? io_cpu_tlb_entry_pfn_1 : io_cpu_tlb_entry_pfn_0; // @[DCache.scala 346:{24,24}]
  wire  _GEN_5155 = data_vpn[0] ? io_cpu_tlb_entry_c_1 : io_cpu_tlb_entry_c_0; // @[DCache.scala 347:{27,27}]
  wire  _GEN_5157 = data_vpn[0] ? io_cpu_tlb_entry_d_1 : io_cpu_tlb_entry_d_0; // @[DCache.scala 348:{24,24}]
  wire [19:0] _GEN_5158 = data_vpn[0] & io_cpu_tlb_entry_v_1 | ~data_vpn[0] & io_cpu_tlb_entry_v_0 ? data_vpn : tlb_vpn; // @[DCache.scala 344:94 345:24 46:20]
  wire [19:0] _GEN_5159 = data_vpn[0] & io_cpu_tlb_entry_v_1 | ~data_vpn[0] & io_cpu_tlb_entry_v_0 ? _GEN_5153 : tlb_ppn
    ; // @[DCache.scala 344:94 346:24 46:20]
  wire  _GEN_5160 = data_vpn[0] & io_cpu_tlb_entry_v_1 | ~data_vpn[0] & io_cpu_tlb_entry_v_0 ? ~_GEN_5155 : tlb_uncached
    ; // @[DCache.scala 344:94 347:24 46:20]
  wire  _GEN_5161 = data_vpn[0] & io_cpu_tlb_entry_v_1 | ~data_vpn[0] & io_cpu_tlb_entry_v_0 ? _GEN_5157 : tlb_dirty; // @[DCache.scala 344:94 348:24 46:20]
  wire  _GEN_5162 = data_vpn[0] & io_cpu_tlb_entry_v_1 | ~data_vpn[0] & io_cpu_tlb_entry_v_0 | tlb_valid; // @[DCache.scala 344:94 349:24 46:20]
  wire [2:0] _GEN_5163 = data_vpn[0] & io_cpu_tlb_entry_v_1 | ~data_vpn[0] & io_cpu_tlb_entry_v_0 ? 3'h0 : 3'h5; // @[DCache.scala 344:94 350:24 352:28]
  wire  _GEN_5164 = data_vpn[0] & io_cpu_tlb_entry_v_1 | ~data_vpn[0] & io_cpu_tlb_entry_v_0 ? data_tlb_invalid : 1'h1; // @[DCache.scala 250:25 344:94 353:28]
  wire  _GEN_5169 = io_cpu_tlb_found ? _GEN_5162 : tlb_valid; // @[DCache.scala 343:30 46:20]
  wire  _GEN_5173 = arvalid & io_axi_ar_ready ? 1'h0 : arvalid; // @[DCache.scala 361:40 362:17 200:24]
  wire [31:0] _GEN_5174 = io_axi_r_valid ? io_axi_r_bits_data : saved_rdata; // @[DCache.scala 364:28 365:21 141:28]
  wire [2:0] _GEN_5175 = io_axi_r_valid ? 3'h5 : state; // @[DCache.scala 364:28 366:21 65:96]
  wire [9:0] _bram_replace_addr_T_4 = bram_replace_addr + 10'h1; // @[DCache.scala 372:50]
  wire [9:0] _GEN_5176 = bram_replace_addr[3:0] != 4'hf ? _bram_replace_addr_T_4 : bram_replace_addr; // @[DCache.scala 371:48 372:29 90:40]
  wire [31:0] _GEN_5194 = _GEN_3187 ? cache_data_1 : cache_data_0; // @[DCache.scala 375:{51,51}]
  wire [31:0] _GEN_5177 = 4'h0 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_0; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5178 = 4'h1 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_1; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5179 = 4'h2 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_2; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5180 = 4'h3 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_3; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5181 = 4'h4 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_4; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5182 = 4'h5 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_5; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5183 = 4'h6 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_6; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5184 = 4'h7 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_7; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5185 = 4'h8 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_8; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5186 = 4'h9 == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_9; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5187 = 4'ha == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_10; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5188 = 4'hb == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_11; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5189 = 4'hc == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_12; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5190 = 4'hd == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_13; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5191 = 4'he == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_14; // @[DCache.scala 375:{51,51} 94:40]
  wire [31:0] _GEN_5192 = 4'hf == bram_read_ready_addr[3:0] ? _GEN_5194 : bram_r_buffer_15; // @[DCache.scala 375:{51,51} 94:40]
  wire  _T_38 = ~aw_handshake; // @[DCache.scala 376:14]
  wire [19:0] _GEN_5196 = _GEN_3187 ? cache_tag_1 : cache_tag_0; // @[Cat.scala 33:{92,92}]
  wire [31:0] _aw_addr_T = {_GEN_5196,fence_line_addr,6'h0}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_5199 = ~aw_handshake ? _aw_addr_T : _GEN_281; // @[DCache.scala 376:29 377:24]
  wire [7:0] _GEN_5200 = ~aw_handshake ? 8'hf : _GEN_285; // @[DCache.scala 376:29 378:24]
  wire [2:0] _GEN_5201 = ~aw_handshake ? 3'h2 : _GEN_282; // @[DCache.scala 376:29 379:24]
  wire  _GEN_5202 = ~aw_handshake | _GEN_276; // @[DCache.scala 376:29 380:24]
  wire [31:0] _GEN_5203 = ~aw_handshake ? _GEN_5194 : _GEN_283; // @[DCache.scala 376:29 381:24]
  wire [3:0] _GEN_5204 = ~aw_handshake ? 4'hf : _GEN_284; // @[DCache.scala 376:29 382:24]
  wire  _GEN_5205 = ~aw_handshake ? 1'h0 : _GEN_278; // @[DCache.scala 376:29 383:24]
  wire  _GEN_5206 = ~aw_handshake | _GEN_277; // @[DCache.scala 376:29 384:24]
  wire  _GEN_5207 = ~aw_handshake | aw_handshake; // @[DCache.scala 376:29 385:24 100:40]
  wire  _GEN_5208 = _T ? 1'h0 : _GEN_5202; // @[DCache.scala 387:30 388:19]
  wire [3:0] _w_data_T_1 = axi_wcnt + 4'h1; // @[DCache.scala 395:26]
  wire  _w_data_T_3 = _w_data_T_1 == bram_read_ready_addr[3:0]; // @[DCache.scala 395:33]
  wire [31:0] _GEN_5212 = 4'h1 == _w_data_T_1 ? bram_r_buffer_1 : bram_r_buffer_0; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5213 = 4'h2 == _w_data_T_1 ? bram_r_buffer_2 : _GEN_5212; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5214 = 4'h3 == _w_data_T_1 ? bram_r_buffer_3 : _GEN_5213; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5215 = 4'h4 == _w_data_T_1 ? bram_r_buffer_4 : _GEN_5214; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5216 = 4'h5 == _w_data_T_1 ? bram_r_buffer_5 : _GEN_5215; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5217 = 4'h6 == _w_data_T_1 ? bram_r_buffer_6 : _GEN_5216; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5218 = 4'h7 == _w_data_T_1 ? bram_r_buffer_7 : _GEN_5217; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5219 = 4'h8 == _w_data_T_1 ? bram_r_buffer_8 : _GEN_5218; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5220 = 4'h9 == _w_data_T_1 ? bram_r_buffer_9 : _GEN_5219; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5221 = 4'ha == _w_data_T_1 ? bram_r_buffer_10 : _GEN_5220; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5222 = 4'hb == _w_data_T_1 ? bram_r_buffer_11 : _GEN_5221; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5223 = 4'hc == _w_data_T_1 ? bram_r_buffer_12 : _GEN_5222; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5224 = 4'hd == _w_data_T_1 ? bram_r_buffer_13 : _GEN_5223; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5225 = 4'he == _w_data_T_1 ? bram_r_buffer_14 : _GEN_5224; // @[DCache.scala 394:{26,26}]
  wire [31:0] _GEN_5226 = 4'hf == _w_data_T_1 ? bram_r_buffer_15 : _GEN_5225; // @[DCache.scala 394:{26,26}]
  wire [31:0] _w_data_T_6 = _w_data_T_3 ? _GEN_5194 : _GEN_5226; // @[DCache.scala 394:26]
  wire  _GEN_5227 = _w_data_T_1 == 4'hf | _GEN_5205; // @[DCache.scala 400:43 401:22]
  wire  _GEN_5228 = w_last ? 1'h0 : _GEN_5206; // @[DCache.scala 391:24 392:20]
  wire [31:0] _GEN_5229 = w_last ? _GEN_5203 : _w_data_T_6; // @[DCache.scala 391:24 394:20]
  wire [3:0] _GEN_5230 = w_last ? axi_wcnt : _w_data_T_1; // @[DCache.scala 391:24 399:22 89:40]
  wire  _GEN_5231 = w_last ? _GEN_5205 : _GEN_5227; // @[DCache.scala 391:24]
  wire  _GEN_5232 = _T_1 ? _GEN_5228 : _GEN_5206; // @[DCache.scala 390:29]
  wire [31:0] _GEN_5233 = _T_1 ? _GEN_5229 : _GEN_5203; // @[DCache.scala 390:29]
  wire [3:0] _GEN_5234 = _T_1 ? _GEN_5230 : axi_wcnt; // @[DCache.scala 390:29 89:40]
  wire  _GEN_5235 = _T_1 ? _GEN_5231 : _GEN_5205; // @[DCache.scala 390:29]
  wire  _GEN_5236 = 6'h0 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_0_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5237 = 6'h0 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_0_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5238 = 6'h1 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_1_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5239 = 6'h1 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_1_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5240 = 6'h2 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_2_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5241 = 6'h2 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_2_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5242 = 6'h3 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_3_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5243 = 6'h3 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_3_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5244 = 6'h4 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_4_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5245 = 6'h4 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_4_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5246 = 6'h5 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_5_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5247 = 6'h5 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_5_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5248 = 6'h6 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_6_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5249 = 6'h6 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_6_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5250 = 6'h7 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_7_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5251 = 6'h7 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_7_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5252 = 6'h8 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_8_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5253 = 6'h8 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_8_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5254 = 6'h9 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_9_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5255 = 6'h9 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_9_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5256 = 6'ha == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_10_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5257 = 6'ha == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_10_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5258 = 6'hb == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_11_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5259 = 6'hb == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_11_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5260 = 6'hc == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_12_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5261 = 6'hc == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_12_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5262 = 6'hd == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_13_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5263 = 6'hd == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_13_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5264 = 6'he == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_14_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5265 = 6'he == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_14_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5266 = 6'hf == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_15_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5267 = 6'hf == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_15_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5268 = 6'h10 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_16_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5269 = 6'h10 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_16_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5270 = 6'h11 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_17_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5271 = 6'h11 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_17_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5272 = 6'h12 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_18_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5273 = 6'h12 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_18_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5274 = 6'h13 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_19_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5275 = 6'h13 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_19_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5276 = 6'h14 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_20_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5277 = 6'h14 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_20_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5278 = 6'h15 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_21_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5279 = 6'h15 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_21_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5280 = 6'h16 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_22_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5281 = 6'h16 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_22_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5282 = 6'h17 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_23_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5283 = 6'h17 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_23_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5284 = 6'h18 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_24_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5285 = 6'h18 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_24_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5286 = 6'h19 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_25_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5287 = 6'h19 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_25_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5288 = 6'h1a == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_26_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5289 = 6'h1a == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_26_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5290 = 6'h1b == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_27_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5291 = 6'h1b == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_27_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5292 = 6'h1c == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_28_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5293 = 6'h1c == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_28_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5294 = 6'h1d == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_29_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5295 = 6'h1d == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_29_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5296 = 6'h1e == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_30_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5297 = 6'h1e == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_30_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5298 = 6'h1f == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_31_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5299 = 6'h1f == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_31_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5300 = 6'h20 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_32_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5301 = 6'h20 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_32_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5302 = 6'h21 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_33_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5303 = 6'h21 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_33_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5304 = 6'h22 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_34_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5305 = 6'h22 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_34_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5306 = 6'h23 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_35_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5307 = 6'h23 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_35_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5308 = 6'h24 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_36_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5309 = 6'h24 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_36_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5310 = 6'h25 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_37_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5311 = 6'h25 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_37_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5312 = 6'h26 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_38_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5313 = 6'h26 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_38_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5314 = 6'h27 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_39_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5315 = 6'h27 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_39_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5316 = 6'h28 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_40_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5317 = 6'h28 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_40_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5318 = 6'h29 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_41_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5319 = 6'h29 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_41_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5320 = 6'h2a == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_42_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5321 = 6'h2a == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_42_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5322 = 6'h2b == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_43_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5323 = 6'h2b == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_43_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5324 = 6'h2c == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_44_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5325 = 6'h2c == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_44_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5326 = 6'h2d == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_45_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5327 = 6'h2d == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_45_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5328 = 6'h2e == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_46_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5329 = 6'h2e == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_46_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5330 = 6'h2f == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_47_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5331 = 6'h2f == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_47_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5332 = 6'h30 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_48_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5333 = 6'h30 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_48_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5334 = 6'h31 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_49_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5335 = 6'h31 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_49_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5336 = 6'h32 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_50_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5337 = 6'h32 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_50_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5338 = 6'h33 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_51_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5339 = 6'h33 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_51_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5340 = 6'h34 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_52_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5341 = 6'h34 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_52_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5342 = 6'h35 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_53_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5343 = 6'h35 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_53_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5344 = 6'h36 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_54_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5345 = 6'h36 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_54_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5346 = 6'h37 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_55_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5347 = 6'h37 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_55_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5348 = 6'h38 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_56_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5349 = 6'h38 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_56_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5350 = 6'h39 == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_57_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5351 = 6'h39 == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_57_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5352 = 6'h3a == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_58_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5353 = 6'h3a == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_58_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5354 = 6'h3b == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_59_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5355 = 6'h3b == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_59_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5356 = 6'h3c == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_60_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5357 = 6'h3c == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_60_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5358 = 6'h3d == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_61_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5359 = 6'h3d == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_61_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5360 = 6'h3e == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_62_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5361 = 6'h3e == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_62_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5362 = 6'h3f == fence_line_addr & ~_GEN_3187 ? 1'h0 : dirty_63_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5363 = 6'h3f == fence_line_addr & _GEN_3187 ? 1'h0 : dirty_63_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5364 = 7'h40 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_64_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5365 = 7'h40 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_64_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5366 = 7'h41 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_65_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5367 = 7'h41 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_65_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5368 = 7'h42 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_66_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5369 = 7'h42 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_66_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5370 = 7'h43 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_67_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5371 = 7'h43 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_67_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5372 = 7'h44 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_68_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5373 = 7'h44 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_68_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5374 = 7'h45 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_69_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5375 = 7'h45 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_69_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5376 = 7'h46 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_70_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5377 = 7'h46 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_70_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5378 = 7'h47 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_71_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5379 = 7'h47 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_71_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5380 = 7'h48 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_72_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5381 = 7'h48 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_72_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5382 = 7'h49 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_73_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5383 = 7'h49 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_73_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5384 = 7'h4a == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_74_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5385 = 7'h4a == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_74_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5386 = 7'h4b == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_75_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5387 = 7'h4b == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_75_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5388 = 7'h4c == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_76_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5389 = 7'h4c == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_76_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5390 = 7'h4d == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_77_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5391 = 7'h4d == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_77_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5392 = 7'h4e == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_78_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5393 = 7'h4e == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_78_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5394 = 7'h4f == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_79_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5395 = 7'h4f == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_79_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5396 = 7'h50 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_80_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5397 = 7'h50 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_80_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5398 = 7'h51 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_81_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5399 = 7'h51 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_81_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5400 = 7'h52 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_82_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5401 = 7'h52 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_82_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5402 = 7'h53 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_83_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5403 = 7'h53 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_83_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5404 = 7'h54 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_84_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5405 = 7'h54 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_84_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5406 = 7'h55 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_85_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5407 = 7'h55 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_85_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5408 = 7'h56 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_86_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5409 = 7'h56 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_86_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5410 = 7'h57 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_87_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5411 = 7'h57 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_87_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5412 = 7'h58 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_88_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5413 = 7'h58 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_88_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5414 = 7'h59 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_89_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5415 = 7'h59 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_89_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5416 = 7'h5a == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_90_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5417 = 7'h5a == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_90_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5418 = 7'h5b == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_91_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5419 = 7'h5b == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_91_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5420 = 7'h5c == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_92_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5421 = 7'h5c == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_92_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5422 = 7'h5d == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_93_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5423 = 7'h5d == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_93_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5424 = 7'h5e == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_94_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5425 = 7'h5e == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_94_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5426 = 7'h5f == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_95_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5427 = 7'h5f == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_95_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5428 = 7'h60 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_96_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5429 = 7'h60 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_96_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5430 = 7'h61 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_97_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5431 = 7'h61 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_97_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5432 = 7'h62 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_98_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5433 = 7'h62 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_98_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5434 = 7'h63 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_99_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5435 = 7'h63 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_99_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5436 = 7'h64 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_100_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5437 = 7'h64 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_100_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5438 = 7'h65 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_101_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5439 = 7'h65 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_101_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5440 = 7'h66 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_102_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5441 = 7'h66 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_102_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5442 = 7'h67 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_103_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5443 = 7'h67 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_103_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5444 = 7'h68 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_104_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5445 = 7'h68 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_104_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5446 = 7'h69 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_105_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5447 = 7'h69 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_105_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5448 = 7'h6a == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_106_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5449 = 7'h6a == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_106_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5450 = 7'h6b == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_107_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5451 = 7'h6b == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_107_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5452 = 7'h6c == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_108_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5453 = 7'h6c == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_108_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5454 = 7'h6d == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_109_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5455 = 7'h6d == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_109_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5456 = 7'h6e == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_110_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5457 = 7'h6e == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_110_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5458 = 7'h6f == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_111_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5459 = 7'h6f == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_111_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5460 = 7'h70 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_112_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5461 = 7'h70 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_112_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5462 = 7'h71 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_113_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5463 = 7'h71 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_113_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5464 = 7'h72 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_114_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5465 = 7'h72 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_114_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5466 = 7'h73 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_115_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5467 = 7'h73 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_115_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5468 = 7'h74 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_116_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5469 = 7'h74 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_116_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5470 = 7'h75 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_117_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5471 = 7'h75 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_117_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5472 = 7'h76 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_118_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5473 = 7'h76 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_118_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5474 = 7'h77 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_119_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5475 = 7'h77 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_119_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5476 = 7'h78 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_120_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5477 = 7'h78 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_120_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5478 = 7'h79 == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_121_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5479 = 7'h79 == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_121_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5480 = 7'h7a == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_122_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5481 = 7'h7a == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_122_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5482 = 7'h7b == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_123_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5483 = 7'h7b == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_123_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5484 = 7'h7c == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_124_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5485 = 7'h7c == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_124_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5486 = 7'h7d == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_125_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5487 = 7'h7d == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_125_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5488 = 7'h7e == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_126_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5489 = 7'h7e == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_126_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5490 = 7'h7f == _GEN_13029 & ~_GEN_3187 ? 1'h0 : dirty_127_0; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5491 = 7'h7f == _GEN_13029 & _GEN_3187 ? 1'h0 : dirty_127_1; // @[DCache.scala 406:{45,45} 69:22]
  wire  _GEN_5492 = io_axi_b_valid ? _GEN_5236 : dirty_0_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5493 = io_axi_b_valid ? _GEN_5237 : dirty_0_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5494 = io_axi_b_valid ? _GEN_5238 : dirty_1_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5495 = io_axi_b_valid ? _GEN_5239 : dirty_1_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5496 = io_axi_b_valid ? _GEN_5240 : dirty_2_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5497 = io_axi_b_valid ? _GEN_5241 : dirty_2_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5498 = io_axi_b_valid ? _GEN_5242 : dirty_3_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5499 = io_axi_b_valid ? _GEN_5243 : dirty_3_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5500 = io_axi_b_valid ? _GEN_5244 : dirty_4_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5501 = io_axi_b_valid ? _GEN_5245 : dirty_4_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5502 = io_axi_b_valid ? _GEN_5246 : dirty_5_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5503 = io_axi_b_valid ? _GEN_5247 : dirty_5_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5504 = io_axi_b_valid ? _GEN_5248 : dirty_6_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5505 = io_axi_b_valid ? _GEN_5249 : dirty_6_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5506 = io_axi_b_valid ? _GEN_5250 : dirty_7_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5507 = io_axi_b_valid ? _GEN_5251 : dirty_7_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5508 = io_axi_b_valid ? _GEN_5252 : dirty_8_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5509 = io_axi_b_valid ? _GEN_5253 : dirty_8_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5510 = io_axi_b_valid ? _GEN_5254 : dirty_9_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5511 = io_axi_b_valid ? _GEN_5255 : dirty_9_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5512 = io_axi_b_valid ? _GEN_5256 : dirty_10_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5513 = io_axi_b_valid ? _GEN_5257 : dirty_10_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5514 = io_axi_b_valid ? _GEN_5258 : dirty_11_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5515 = io_axi_b_valid ? _GEN_5259 : dirty_11_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5516 = io_axi_b_valid ? _GEN_5260 : dirty_12_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5517 = io_axi_b_valid ? _GEN_5261 : dirty_12_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5518 = io_axi_b_valid ? _GEN_5262 : dirty_13_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5519 = io_axi_b_valid ? _GEN_5263 : dirty_13_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5520 = io_axi_b_valid ? _GEN_5264 : dirty_14_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5521 = io_axi_b_valid ? _GEN_5265 : dirty_14_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5522 = io_axi_b_valid ? _GEN_5266 : dirty_15_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5523 = io_axi_b_valid ? _GEN_5267 : dirty_15_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5524 = io_axi_b_valid ? _GEN_5268 : dirty_16_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5525 = io_axi_b_valid ? _GEN_5269 : dirty_16_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5526 = io_axi_b_valid ? _GEN_5270 : dirty_17_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5527 = io_axi_b_valid ? _GEN_5271 : dirty_17_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5528 = io_axi_b_valid ? _GEN_5272 : dirty_18_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5529 = io_axi_b_valid ? _GEN_5273 : dirty_18_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5530 = io_axi_b_valid ? _GEN_5274 : dirty_19_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5531 = io_axi_b_valid ? _GEN_5275 : dirty_19_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5532 = io_axi_b_valid ? _GEN_5276 : dirty_20_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5533 = io_axi_b_valid ? _GEN_5277 : dirty_20_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5534 = io_axi_b_valid ? _GEN_5278 : dirty_21_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5535 = io_axi_b_valid ? _GEN_5279 : dirty_21_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5536 = io_axi_b_valid ? _GEN_5280 : dirty_22_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5537 = io_axi_b_valid ? _GEN_5281 : dirty_22_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5538 = io_axi_b_valid ? _GEN_5282 : dirty_23_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5539 = io_axi_b_valid ? _GEN_5283 : dirty_23_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5540 = io_axi_b_valid ? _GEN_5284 : dirty_24_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5541 = io_axi_b_valid ? _GEN_5285 : dirty_24_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5542 = io_axi_b_valid ? _GEN_5286 : dirty_25_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5543 = io_axi_b_valid ? _GEN_5287 : dirty_25_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5544 = io_axi_b_valid ? _GEN_5288 : dirty_26_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5545 = io_axi_b_valid ? _GEN_5289 : dirty_26_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5546 = io_axi_b_valid ? _GEN_5290 : dirty_27_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5547 = io_axi_b_valid ? _GEN_5291 : dirty_27_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5548 = io_axi_b_valid ? _GEN_5292 : dirty_28_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5549 = io_axi_b_valid ? _GEN_5293 : dirty_28_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5550 = io_axi_b_valid ? _GEN_5294 : dirty_29_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5551 = io_axi_b_valid ? _GEN_5295 : dirty_29_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5552 = io_axi_b_valid ? _GEN_5296 : dirty_30_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5553 = io_axi_b_valid ? _GEN_5297 : dirty_30_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5554 = io_axi_b_valid ? _GEN_5298 : dirty_31_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5555 = io_axi_b_valid ? _GEN_5299 : dirty_31_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5556 = io_axi_b_valid ? _GEN_5300 : dirty_32_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5557 = io_axi_b_valid ? _GEN_5301 : dirty_32_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5558 = io_axi_b_valid ? _GEN_5302 : dirty_33_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5559 = io_axi_b_valid ? _GEN_5303 : dirty_33_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5560 = io_axi_b_valid ? _GEN_5304 : dirty_34_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5561 = io_axi_b_valid ? _GEN_5305 : dirty_34_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5562 = io_axi_b_valid ? _GEN_5306 : dirty_35_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5563 = io_axi_b_valid ? _GEN_5307 : dirty_35_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5564 = io_axi_b_valid ? _GEN_5308 : dirty_36_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5565 = io_axi_b_valid ? _GEN_5309 : dirty_36_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5566 = io_axi_b_valid ? _GEN_5310 : dirty_37_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5567 = io_axi_b_valid ? _GEN_5311 : dirty_37_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5568 = io_axi_b_valid ? _GEN_5312 : dirty_38_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5569 = io_axi_b_valid ? _GEN_5313 : dirty_38_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5570 = io_axi_b_valid ? _GEN_5314 : dirty_39_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5571 = io_axi_b_valid ? _GEN_5315 : dirty_39_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5572 = io_axi_b_valid ? _GEN_5316 : dirty_40_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5573 = io_axi_b_valid ? _GEN_5317 : dirty_40_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5574 = io_axi_b_valid ? _GEN_5318 : dirty_41_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5575 = io_axi_b_valid ? _GEN_5319 : dirty_41_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5576 = io_axi_b_valid ? _GEN_5320 : dirty_42_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5577 = io_axi_b_valid ? _GEN_5321 : dirty_42_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5578 = io_axi_b_valid ? _GEN_5322 : dirty_43_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5579 = io_axi_b_valid ? _GEN_5323 : dirty_43_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5580 = io_axi_b_valid ? _GEN_5324 : dirty_44_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5581 = io_axi_b_valid ? _GEN_5325 : dirty_44_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5582 = io_axi_b_valid ? _GEN_5326 : dirty_45_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5583 = io_axi_b_valid ? _GEN_5327 : dirty_45_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5584 = io_axi_b_valid ? _GEN_5328 : dirty_46_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5585 = io_axi_b_valid ? _GEN_5329 : dirty_46_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5586 = io_axi_b_valid ? _GEN_5330 : dirty_47_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5587 = io_axi_b_valid ? _GEN_5331 : dirty_47_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5588 = io_axi_b_valid ? _GEN_5332 : dirty_48_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5589 = io_axi_b_valid ? _GEN_5333 : dirty_48_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5590 = io_axi_b_valid ? _GEN_5334 : dirty_49_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5591 = io_axi_b_valid ? _GEN_5335 : dirty_49_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5592 = io_axi_b_valid ? _GEN_5336 : dirty_50_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5593 = io_axi_b_valid ? _GEN_5337 : dirty_50_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5594 = io_axi_b_valid ? _GEN_5338 : dirty_51_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5595 = io_axi_b_valid ? _GEN_5339 : dirty_51_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5596 = io_axi_b_valid ? _GEN_5340 : dirty_52_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5597 = io_axi_b_valid ? _GEN_5341 : dirty_52_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5598 = io_axi_b_valid ? _GEN_5342 : dirty_53_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5599 = io_axi_b_valid ? _GEN_5343 : dirty_53_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5600 = io_axi_b_valid ? _GEN_5344 : dirty_54_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5601 = io_axi_b_valid ? _GEN_5345 : dirty_54_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5602 = io_axi_b_valid ? _GEN_5346 : dirty_55_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5603 = io_axi_b_valid ? _GEN_5347 : dirty_55_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5604 = io_axi_b_valid ? _GEN_5348 : dirty_56_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5605 = io_axi_b_valid ? _GEN_5349 : dirty_56_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5606 = io_axi_b_valid ? _GEN_5350 : dirty_57_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5607 = io_axi_b_valid ? _GEN_5351 : dirty_57_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5608 = io_axi_b_valid ? _GEN_5352 : dirty_58_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5609 = io_axi_b_valid ? _GEN_5353 : dirty_58_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5610 = io_axi_b_valid ? _GEN_5354 : dirty_59_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5611 = io_axi_b_valid ? _GEN_5355 : dirty_59_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5612 = io_axi_b_valid ? _GEN_5356 : dirty_60_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5613 = io_axi_b_valid ? _GEN_5357 : dirty_60_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5614 = io_axi_b_valid ? _GEN_5358 : dirty_61_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5615 = io_axi_b_valid ? _GEN_5359 : dirty_61_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5616 = io_axi_b_valid ? _GEN_5360 : dirty_62_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5617 = io_axi_b_valid ? _GEN_5361 : dirty_62_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5618 = io_axi_b_valid ? _GEN_5362 : dirty_63_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5619 = io_axi_b_valid ? _GEN_5363 : dirty_63_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5620 = io_axi_b_valid ? _GEN_5364 : dirty_64_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5621 = io_axi_b_valid ? _GEN_5365 : dirty_64_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5622 = io_axi_b_valid ? _GEN_5366 : dirty_65_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5623 = io_axi_b_valid ? _GEN_5367 : dirty_65_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5624 = io_axi_b_valid ? _GEN_5368 : dirty_66_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5625 = io_axi_b_valid ? _GEN_5369 : dirty_66_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5626 = io_axi_b_valid ? _GEN_5370 : dirty_67_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5627 = io_axi_b_valid ? _GEN_5371 : dirty_67_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5628 = io_axi_b_valid ? _GEN_5372 : dirty_68_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5629 = io_axi_b_valid ? _GEN_5373 : dirty_68_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5630 = io_axi_b_valid ? _GEN_5374 : dirty_69_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5631 = io_axi_b_valid ? _GEN_5375 : dirty_69_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5632 = io_axi_b_valid ? _GEN_5376 : dirty_70_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5633 = io_axi_b_valid ? _GEN_5377 : dirty_70_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5634 = io_axi_b_valid ? _GEN_5378 : dirty_71_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5635 = io_axi_b_valid ? _GEN_5379 : dirty_71_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5636 = io_axi_b_valid ? _GEN_5380 : dirty_72_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5637 = io_axi_b_valid ? _GEN_5381 : dirty_72_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5638 = io_axi_b_valid ? _GEN_5382 : dirty_73_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5639 = io_axi_b_valid ? _GEN_5383 : dirty_73_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5640 = io_axi_b_valid ? _GEN_5384 : dirty_74_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5641 = io_axi_b_valid ? _GEN_5385 : dirty_74_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5642 = io_axi_b_valid ? _GEN_5386 : dirty_75_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5643 = io_axi_b_valid ? _GEN_5387 : dirty_75_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5644 = io_axi_b_valid ? _GEN_5388 : dirty_76_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5645 = io_axi_b_valid ? _GEN_5389 : dirty_76_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5646 = io_axi_b_valid ? _GEN_5390 : dirty_77_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5647 = io_axi_b_valid ? _GEN_5391 : dirty_77_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5648 = io_axi_b_valid ? _GEN_5392 : dirty_78_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5649 = io_axi_b_valid ? _GEN_5393 : dirty_78_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5650 = io_axi_b_valid ? _GEN_5394 : dirty_79_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5651 = io_axi_b_valid ? _GEN_5395 : dirty_79_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5652 = io_axi_b_valid ? _GEN_5396 : dirty_80_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5653 = io_axi_b_valid ? _GEN_5397 : dirty_80_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5654 = io_axi_b_valid ? _GEN_5398 : dirty_81_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5655 = io_axi_b_valid ? _GEN_5399 : dirty_81_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5656 = io_axi_b_valid ? _GEN_5400 : dirty_82_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5657 = io_axi_b_valid ? _GEN_5401 : dirty_82_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5658 = io_axi_b_valid ? _GEN_5402 : dirty_83_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5659 = io_axi_b_valid ? _GEN_5403 : dirty_83_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5660 = io_axi_b_valid ? _GEN_5404 : dirty_84_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5661 = io_axi_b_valid ? _GEN_5405 : dirty_84_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5662 = io_axi_b_valid ? _GEN_5406 : dirty_85_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5663 = io_axi_b_valid ? _GEN_5407 : dirty_85_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5664 = io_axi_b_valid ? _GEN_5408 : dirty_86_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5665 = io_axi_b_valid ? _GEN_5409 : dirty_86_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5666 = io_axi_b_valid ? _GEN_5410 : dirty_87_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5667 = io_axi_b_valid ? _GEN_5411 : dirty_87_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5668 = io_axi_b_valid ? _GEN_5412 : dirty_88_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5669 = io_axi_b_valid ? _GEN_5413 : dirty_88_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5670 = io_axi_b_valid ? _GEN_5414 : dirty_89_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5671 = io_axi_b_valid ? _GEN_5415 : dirty_89_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5672 = io_axi_b_valid ? _GEN_5416 : dirty_90_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5673 = io_axi_b_valid ? _GEN_5417 : dirty_90_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5674 = io_axi_b_valid ? _GEN_5418 : dirty_91_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5675 = io_axi_b_valid ? _GEN_5419 : dirty_91_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5676 = io_axi_b_valid ? _GEN_5420 : dirty_92_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5677 = io_axi_b_valid ? _GEN_5421 : dirty_92_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5678 = io_axi_b_valid ? _GEN_5422 : dirty_93_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5679 = io_axi_b_valid ? _GEN_5423 : dirty_93_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5680 = io_axi_b_valid ? _GEN_5424 : dirty_94_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5681 = io_axi_b_valid ? _GEN_5425 : dirty_94_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5682 = io_axi_b_valid ? _GEN_5426 : dirty_95_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5683 = io_axi_b_valid ? _GEN_5427 : dirty_95_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5684 = io_axi_b_valid ? _GEN_5428 : dirty_96_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5685 = io_axi_b_valid ? _GEN_5429 : dirty_96_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5686 = io_axi_b_valid ? _GEN_5430 : dirty_97_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5687 = io_axi_b_valid ? _GEN_5431 : dirty_97_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5688 = io_axi_b_valid ? _GEN_5432 : dirty_98_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5689 = io_axi_b_valid ? _GEN_5433 : dirty_98_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5690 = io_axi_b_valid ? _GEN_5434 : dirty_99_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5691 = io_axi_b_valid ? _GEN_5435 : dirty_99_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5692 = io_axi_b_valid ? _GEN_5436 : dirty_100_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5693 = io_axi_b_valid ? _GEN_5437 : dirty_100_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5694 = io_axi_b_valid ? _GEN_5438 : dirty_101_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5695 = io_axi_b_valid ? _GEN_5439 : dirty_101_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5696 = io_axi_b_valid ? _GEN_5440 : dirty_102_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5697 = io_axi_b_valid ? _GEN_5441 : dirty_102_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5698 = io_axi_b_valid ? _GEN_5442 : dirty_103_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5699 = io_axi_b_valid ? _GEN_5443 : dirty_103_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5700 = io_axi_b_valid ? _GEN_5444 : dirty_104_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5701 = io_axi_b_valid ? _GEN_5445 : dirty_104_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5702 = io_axi_b_valid ? _GEN_5446 : dirty_105_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5703 = io_axi_b_valid ? _GEN_5447 : dirty_105_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5704 = io_axi_b_valid ? _GEN_5448 : dirty_106_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5705 = io_axi_b_valid ? _GEN_5449 : dirty_106_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5706 = io_axi_b_valid ? _GEN_5450 : dirty_107_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5707 = io_axi_b_valid ? _GEN_5451 : dirty_107_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5708 = io_axi_b_valid ? _GEN_5452 : dirty_108_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5709 = io_axi_b_valid ? _GEN_5453 : dirty_108_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5710 = io_axi_b_valid ? _GEN_5454 : dirty_109_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5711 = io_axi_b_valid ? _GEN_5455 : dirty_109_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5712 = io_axi_b_valid ? _GEN_5456 : dirty_110_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5713 = io_axi_b_valid ? _GEN_5457 : dirty_110_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5714 = io_axi_b_valid ? _GEN_5458 : dirty_111_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5715 = io_axi_b_valid ? _GEN_5459 : dirty_111_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5716 = io_axi_b_valid ? _GEN_5460 : dirty_112_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5717 = io_axi_b_valid ? _GEN_5461 : dirty_112_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5718 = io_axi_b_valid ? _GEN_5462 : dirty_113_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5719 = io_axi_b_valid ? _GEN_5463 : dirty_113_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5720 = io_axi_b_valid ? _GEN_5464 : dirty_114_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5721 = io_axi_b_valid ? _GEN_5465 : dirty_114_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5722 = io_axi_b_valid ? _GEN_5466 : dirty_115_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5723 = io_axi_b_valid ? _GEN_5467 : dirty_115_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5724 = io_axi_b_valid ? _GEN_5468 : dirty_116_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5725 = io_axi_b_valid ? _GEN_5469 : dirty_116_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5726 = io_axi_b_valid ? _GEN_5470 : dirty_117_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5727 = io_axi_b_valid ? _GEN_5471 : dirty_117_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5728 = io_axi_b_valid ? _GEN_5472 : dirty_118_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5729 = io_axi_b_valid ? _GEN_5473 : dirty_118_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5730 = io_axi_b_valid ? _GEN_5474 : dirty_119_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5731 = io_axi_b_valid ? _GEN_5475 : dirty_119_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5732 = io_axi_b_valid ? _GEN_5476 : dirty_120_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5733 = io_axi_b_valid ? _GEN_5477 : dirty_120_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5734 = io_axi_b_valid ? _GEN_5478 : dirty_121_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5735 = io_axi_b_valid ? _GEN_5479 : dirty_121_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5736 = io_axi_b_valid ? _GEN_5480 : dirty_122_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5737 = io_axi_b_valid ? _GEN_5481 : dirty_122_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5738 = io_axi_b_valid ? _GEN_5482 : dirty_123_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5739 = io_axi_b_valid ? _GEN_5483 : dirty_123_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5740 = io_axi_b_valid ? _GEN_5484 : dirty_124_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5741 = io_axi_b_valid ? _GEN_5485 : dirty_124_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5742 = io_axi_b_valid ? _GEN_5486 : dirty_125_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5743 = io_axi_b_valid ? _GEN_5487 : dirty_125_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5744 = io_axi_b_valid ? _GEN_5488 : dirty_126_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5745 = io_axi_b_valid ? _GEN_5489 : dirty_126_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5746 = io_axi_b_valid ? _GEN_5490 : dirty_127_0; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5747 = io_axi_b_valid ? _GEN_5491 : dirty_127_1; // @[DCache.scala 405:30 69:22]
  wire  _GEN_5748 = io_axi_b_valid ? 1'h0 : fence_working; // @[DCache.scala 405:30 407:45 97:40]
  wire  _GEN_5749 = io_axi_b_valid ? 1'h0 : bram_use_replace_addr; // @[DCache.scala 405:30 408:45 95:40]
  wire [2:0] _GEN_5750 = io_axi_b_valid ? 3'h0 : state; // @[DCache.scala 405:30 409:45 65:96]
  wire [9:0] _GEN_5751 = fence_working ? _GEN_5176 : _bram_replace_addr_T_4; // @[DCache.scala 370:27 414:27]
  wire [9:0] _GEN_5752 = fence_working ? bram_replace_addr : bram_read_ready_addr; // @[DCache.scala 370:27 374:51 91:40]
  wire [31:0] _GEN_5753 = fence_working ? _GEN_5177 : bram_r_buffer_0; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5754 = fence_working ? _GEN_5178 : bram_r_buffer_1; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5755 = fence_working ? _GEN_5179 : bram_r_buffer_2; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5756 = fence_working ? _GEN_5180 : bram_r_buffer_3; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5757 = fence_working ? _GEN_5181 : bram_r_buffer_4; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5758 = fence_working ? _GEN_5182 : bram_r_buffer_5; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5759 = fence_working ? _GEN_5183 : bram_r_buffer_6; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5760 = fence_working ? _GEN_5184 : bram_r_buffer_7; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5761 = fence_working ? _GEN_5185 : bram_r_buffer_8; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5762 = fence_working ? _GEN_5186 : bram_r_buffer_9; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5763 = fence_working ? _GEN_5187 : bram_r_buffer_10; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5764 = fence_working ? _GEN_5188 : bram_r_buffer_11; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5765 = fence_working ? _GEN_5189 : bram_r_buffer_12; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5766 = fence_working ? _GEN_5190 : bram_r_buffer_13; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5767 = fence_working ? _GEN_5191 : bram_r_buffer_14; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5768 = fence_working ? _GEN_5192 : bram_r_buffer_15; // @[DCache.scala 370:27 94:40]
  wire [31:0] _GEN_5769 = fence_working ? _GEN_5199 : _GEN_281; // @[DCache.scala 370:27]
  wire [7:0] _GEN_5770 = fence_working ? _GEN_5200 : _GEN_285; // @[DCache.scala 370:27]
  wire [2:0] _GEN_5771 = fence_working ? _GEN_5201 : _GEN_282; // @[DCache.scala 370:27]
  wire  _GEN_5772 = fence_working ? _GEN_5208 : _GEN_276; // @[DCache.scala 370:27]
  wire [31:0] _GEN_5773 = fence_working ? _GEN_5233 : _GEN_283; // @[DCache.scala 370:27]
  wire [3:0] _GEN_5774 = fence_working ? _GEN_5204 : _GEN_284; // @[DCache.scala 370:27]
  wire  _GEN_5775 = fence_working ? _GEN_5235 : _GEN_278; // @[DCache.scala 370:27]
  wire  _GEN_5776 = fence_working ? _GEN_5232 : _GEN_277; // @[DCache.scala 370:27]
  wire  _GEN_5777 = fence_working & _GEN_5207; // @[DCache.scala 370:27 412:27]
  wire [3:0] _GEN_5778 = fence_working ? _GEN_5234 : axi_wcnt; // @[DCache.scala 370:27 89:40]
  wire  _GEN_5779 = fence_working ? _GEN_5492 : dirty_0_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5780 = fence_working ? _GEN_5493 : dirty_0_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5781 = fence_working ? _GEN_5494 : dirty_1_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5782 = fence_working ? _GEN_5495 : dirty_1_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5783 = fence_working ? _GEN_5496 : dirty_2_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5784 = fence_working ? _GEN_5497 : dirty_2_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5785 = fence_working ? _GEN_5498 : dirty_3_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5786 = fence_working ? _GEN_5499 : dirty_3_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5787 = fence_working ? _GEN_5500 : dirty_4_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5788 = fence_working ? _GEN_5501 : dirty_4_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5789 = fence_working ? _GEN_5502 : dirty_5_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5790 = fence_working ? _GEN_5503 : dirty_5_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5791 = fence_working ? _GEN_5504 : dirty_6_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5792 = fence_working ? _GEN_5505 : dirty_6_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5793 = fence_working ? _GEN_5506 : dirty_7_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5794 = fence_working ? _GEN_5507 : dirty_7_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5795 = fence_working ? _GEN_5508 : dirty_8_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5796 = fence_working ? _GEN_5509 : dirty_8_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5797 = fence_working ? _GEN_5510 : dirty_9_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5798 = fence_working ? _GEN_5511 : dirty_9_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5799 = fence_working ? _GEN_5512 : dirty_10_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5800 = fence_working ? _GEN_5513 : dirty_10_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5801 = fence_working ? _GEN_5514 : dirty_11_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5802 = fence_working ? _GEN_5515 : dirty_11_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5803 = fence_working ? _GEN_5516 : dirty_12_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5804 = fence_working ? _GEN_5517 : dirty_12_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5805 = fence_working ? _GEN_5518 : dirty_13_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5806 = fence_working ? _GEN_5519 : dirty_13_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5807 = fence_working ? _GEN_5520 : dirty_14_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5808 = fence_working ? _GEN_5521 : dirty_14_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5809 = fence_working ? _GEN_5522 : dirty_15_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5810 = fence_working ? _GEN_5523 : dirty_15_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5811 = fence_working ? _GEN_5524 : dirty_16_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5812 = fence_working ? _GEN_5525 : dirty_16_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5813 = fence_working ? _GEN_5526 : dirty_17_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5814 = fence_working ? _GEN_5527 : dirty_17_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5815 = fence_working ? _GEN_5528 : dirty_18_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5816 = fence_working ? _GEN_5529 : dirty_18_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5817 = fence_working ? _GEN_5530 : dirty_19_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5818 = fence_working ? _GEN_5531 : dirty_19_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5819 = fence_working ? _GEN_5532 : dirty_20_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5820 = fence_working ? _GEN_5533 : dirty_20_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5821 = fence_working ? _GEN_5534 : dirty_21_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5822 = fence_working ? _GEN_5535 : dirty_21_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5823 = fence_working ? _GEN_5536 : dirty_22_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5824 = fence_working ? _GEN_5537 : dirty_22_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5825 = fence_working ? _GEN_5538 : dirty_23_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5826 = fence_working ? _GEN_5539 : dirty_23_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5827 = fence_working ? _GEN_5540 : dirty_24_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5828 = fence_working ? _GEN_5541 : dirty_24_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5829 = fence_working ? _GEN_5542 : dirty_25_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5830 = fence_working ? _GEN_5543 : dirty_25_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5831 = fence_working ? _GEN_5544 : dirty_26_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5832 = fence_working ? _GEN_5545 : dirty_26_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5833 = fence_working ? _GEN_5546 : dirty_27_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5834 = fence_working ? _GEN_5547 : dirty_27_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5835 = fence_working ? _GEN_5548 : dirty_28_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5836 = fence_working ? _GEN_5549 : dirty_28_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5837 = fence_working ? _GEN_5550 : dirty_29_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5838 = fence_working ? _GEN_5551 : dirty_29_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5839 = fence_working ? _GEN_5552 : dirty_30_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5840 = fence_working ? _GEN_5553 : dirty_30_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5841 = fence_working ? _GEN_5554 : dirty_31_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5842 = fence_working ? _GEN_5555 : dirty_31_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5843 = fence_working ? _GEN_5556 : dirty_32_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5844 = fence_working ? _GEN_5557 : dirty_32_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5845 = fence_working ? _GEN_5558 : dirty_33_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5846 = fence_working ? _GEN_5559 : dirty_33_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5847 = fence_working ? _GEN_5560 : dirty_34_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5848 = fence_working ? _GEN_5561 : dirty_34_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5849 = fence_working ? _GEN_5562 : dirty_35_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5850 = fence_working ? _GEN_5563 : dirty_35_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5851 = fence_working ? _GEN_5564 : dirty_36_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5852 = fence_working ? _GEN_5565 : dirty_36_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5853 = fence_working ? _GEN_5566 : dirty_37_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5854 = fence_working ? _GEN_5567 : dirty_37_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5855 = fence_working ? _GEN_5568 : dirty_38_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5856 = fence_working ? _GEN_5569 : dirty_38_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5857 = fence_working ? _GEN_5570 : dirty_39_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5858 = fence_working ? _GEN_5571 : dirty_39_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5859 = fence_working ? _GEN_5572 : dirty_40_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5860 = fence_working ? _GEN_5573 : dirty_40_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5861 = fence_working ? _GEN_5574 : dirty_41_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5862 = fence_working ? _GEN_5575 : dirty_41_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5863 = fence_working ? _GEN_5576 : dirty_42_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5864 = fence_working ? _GEN_5577 : dirty_42_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5865 = fence_working ? _GEN_5578 : dirty_43_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5866 = fence_working ? _GEN_5579 : dirty_43_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5867 = fence_working ? _GEN_5580 : dirty_44_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5868 = fence_working ? _GEN_5581 : dirty_44_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5869 = fence_working ? _GEN_5582 : dirty_45_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5870 = fence_working ? _GEN_5583 : dirty_45_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5871 = fence_working ? _GEN_5584 : dirty_46_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5872 = fence_working ? _GEN_5585 : dirty_46_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5873 = fence_working ? _GEN_5586 : dirty_47_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5874 = fence_working ? _GEN_5587 : dirty_47_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5875 = fence_working ? _GEN_5588 : dirty_48_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5876 = fence_working ? _GEN_5589 : dirty_48_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5877 = fence_working ? _GEN_5590 : dirty_49_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5878 = fence_working ? _GEN_5591 : dirty_49_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5879 = fence_working ? _GEN_5592 : dirty_50_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5880 = fence_working ? _GEN_5593 : dirty_50_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5881 = fence_working ? _GEN_5594 : dirty_51_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5882 = fence_working ? _GEN_5595 : dirty_51_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5883 = fence_working ? _GEN_5596 : dirty_52_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5884 = fence_working ? _GEN_5597 : dirty_52_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5885 = fence_working ? _GEN_5598 : dirty_53_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5886 = fence_working ? _GEN_5599 : dirty_53_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5887 = fence_working ? _GEN_5600 : dirty_54_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5888 = fence_working ? _GEN_5601 : dirty_54_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5889 = fence_working ? _GEN_5602 : dirty_55_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5890 = fence_working ? _GEN_5603 : dirty_55_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5891 = fence_working ? _GEN_5604 : dirty_56_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5892 = fence_working ? _GEN_5605 : dirty_56_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5893 = fence_working ? _GEN_5606 : dirty_57_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5894 = fence_working ? _GEN_5607 : dirty_57_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5895 = fence_working ? _GEN_5608 : dirty_58_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5896 = fence_working ? _GEN_5609 : dirty_58_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5897 = fence_working ? _GEN_5610 : dirty_59_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5898 = fence_working ? _GEN_5611 : dirty_59_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5899 = fence_working ? _GEN_5612 : dirty_60_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5900 = fence_working ? _GEN_5613 : dirty_60_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5901 = fence_working ? _GEN_5614 : dirty_61_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5902 = fence_working ? _GEN_5615 : dirty_61_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5903 = fence_working ? _GEN_5616 : dirty_62_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5904 = fence_working ? _GEN_5617 : dirty_62_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5905 = fence_working ? _GEN_5618 : dirty_63_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5906 = fence_working ? _GEN_5619 : dirty_63_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5907 = fence_working ? _GEN_5620 : dirty_64_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5908 = fence_working ? _GEN_5621 : dirty_64_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5909 = fence_working ? _GEN_5622 : dirty_65_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5910 = fence_working ? _GEN_5623 : dirty_65_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5911 = fence_working ? _GEN_5624 : dirty_66_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5912 = fence_working ? _GEN_5625 : dirty_66_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5913 = fence_working ? _GEN_5626 : dirty_67_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5914 = fence_working ? _GEN_5627 : dirty_67_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5915 = fence_working ? _GEN_5628 : dirty_68_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5916 = fence_working ? _GEN_5629 : dirty_68_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5917 = fence_working ? _GEN_5630 : dirty_69_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5918 = fence_working ? _GEN_5631 : dirty_69_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5919 = fence_working ? _GEN_5632 : dirty_70_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5920 = fence_working ? _GEN_5633 : dirty_70_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5921 = fence_working ? _GEN_5634 : dirty_71_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5922 = fence_working ? _GEN_5635 : dirty_71_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5923 = fence_working ? _GEN_5636 : dirty_72_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5924 = fence_working ? _GEN_5637 : dirty_72_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5925 = fence_working ? _GEN_5638 : dirty_73_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5926 = fence_working ? _GEN_5639 : dirty_73_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5927 = fence_working ? _GEN_5640 : dirty_74_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5928 = fence_working ? _GEN_5641 : dirty_74_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5929 = fence_working ? _GEN_5642 : dirty_75_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5930 = fence_working ? _GEN_5643 : dirty_75_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5931 = fence_working ? _GEN_5644 : dirty_76_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5932 = fence_working ? _GEN_5645 : dirty_76_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5933 = fence_working ? _GEN_5646 : dirty_77_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5934 = fence_working ? _GEN_5647 : dirty_77_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5935 = fence_working ? _GEN_5648 : dirty_78_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5936 = fence_working ? _GEN_5649 : dirty_78_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5937 = fence_working ? _GEN_5650 : dirty_79_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5938 = fence_working ? _GEN_5651 : dirty_79_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5939 = fence_working ? _GEN_5652 : dirty_80_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5940 = fence_working ? _GEN_5653 : dirty_80_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5941 = fence_working ? _GEN_5654 : dirty_81_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5942 = fence_working ? _GEN_5655 : dirty_81_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5943 = fence_working ? _GEN_5656 : dirty_82_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5944 = fence_working ? _GEN_5657 : dirty_82_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5945 = fence_working ? _GEN_5658 : dirty_83_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5946 = fence_working ? _GEN_5659 : dirty_83_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5947 = fence_working ? _GEN_5660 : dirty_84_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5948 = fence_working ? _GEN_5661 : dirty_84_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5949 = fence_working ? _GEN_5662 : dirty_85_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5950 = fence_working ? _GEN_5663 : dirty_85_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5951 = fence_working ? _GEN_5664 : dirty_86_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5952 = fence_working ? _GEN_5665 : dirty_86_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5953 = fence_working ? _GEN_5666 : dirty_87_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5954 = fence_working ? _GEN_5667 : dirty_87_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5955 = fence_working ? _GEN_5668 : dirty_88_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5956 = fence_working ? _GEN_5669 : dirty_88_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5957 = fence_working ? _GEN_5670 : dirty_89_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5958 = fence_working ? _GEN_5671 : dirty_89_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5959 = fence_working ? _GEN_5672 : dirty_90_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5960 = fence_working ? _GEN_5673 : dirty_90_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5961 = fence_working ? _GEN_5674 : dirty_91_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5962 = fence_working ? _GEN_5675 : dirty_91_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5963 = fence_working ? _GEN_5676 : dirty_92_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5964 = fence_working ? _GEN_5677 : dirty_92_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5965 = fence_working ? _GEN_5678 : dirty_93_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5966 = fence_working ? _GEN_5679 : dirty_93_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5967 = fence_working ? _GEN_5680 : dirty_94_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5968 = fence_working ? _GEN_5681 : dirty_94_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5969 = fence_working ? _GEN_5682 : dirty_95_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5970 = fence_working ? _GEN_5683 : dirty_95_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5971 = fence_working ? _GEN_5684 : dirty_96_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5972 = fence_working ? _GEN_5685 : dirty_96_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5973 = fence_working ? _GEN_5686 : dirty_97_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5974 = fence_working ? _GEN_5687 : dirty_97_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5975 = fence_working ? _GEN_5688 : dirty_98_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5976 = fence_working ? _GEN_5689 : dirty_98_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5977 = fence_working ? _GEN_5690 : dirty_99_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5978 = fence_working ? _GEN_5691 : dirty_99_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5979 = fence_working ? _GEN_5692 : dirty_100_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5980 = fence_working ? _GEN_5693 : dirty_100_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5981 = fence_working ? _GEN_5694 : dirty_101_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5982 = fence_working ? _GEN_5695 : dirty_101_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5983 = fence_working ? _GEN_5696 : dirty_102_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5984 = fence_working ? _GEN_5697 : dirty_102_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5985 = fence_working ? _GEN_5698 : dirty_103_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5986 = fence_working ? _GEN_5699 : dirty_103_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5987 = fence_working ? _GEN_5700 : dirty_104_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5988 = fence_working ? _GEN_5701 : dirty_104_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5989 = fence_working ? _GEN_5702 : dirty_105_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5990 = fence_working ? _GEN_5703 : dirty_105_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5991 = fence_working ? _GEN_5704 : dirty_106_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5992 = fence_working ? _GEN_5705 : dirty_106_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5993 = fence_working ? _GEN_5706 : dirty_107_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5994 = fence_working ? _GEN_5707 : dirty_107_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5995 = fence_working ? _GEN_5708 : dirty_108_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5996 = fence_working ? _GEN_5709 : dirty_108_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5997 = fence_working ? _GEN_5710 : dirty_109_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5998 = fence_working ? _GEN_5711 : dirty_109_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_5999 = fence_working ? _GEN_5712 : dirty_110_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6000 = fence_working ? _GEN_5713 : dirty_110_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6001 = fence_working ? _GEN_5714 : dirty_111_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6002 = fence_working ? _GEN_5715 : dirty_111_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6003 = fence_working ? _GEN_5716 : dirty_112_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6004 = fence_working ? _GEN_5717 : dirty_112_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6005 = fence_working ? _GEN_5718 : dirty_113_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6006 = fence_working ? _GEN_5719 : dirty_113_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6007 = fence_working ? _GEN_5720 : dirty_114_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6008 = fence_working ? _GEN_5721 : dirty_114_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6009 = fence_working ? _GEN_5722 : dirty_115_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6010 = fence_working ? _GEN_5723 : dirty_115_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6011 = fence_working ? _GEN_5724 : dirty_116_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6012 = fence_working ? _GEN_5725 : dirty_116_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6013 = fence_working ? _GEN_5726 : dirty_117_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6014 = fence_working ? _GEN_5727 : dirty_117_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6015 = fence_working ? _GEN_5728 : dirty_118_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6016 = fence_working ? _GEN_5729 : dirty_118_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6017 = fence_working ? _GEN_5730 : dirty_119_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6018 = fence_working ? _GEN_5731 : dirty_119_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6019 = fence_working ? _GEN_5732 : dirty_120_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6020 = fence_working ? _GEN_5733 : dirty_120_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6021 = fence_working ? _GEN_5734 : dirty_121_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6022 = fence_working ? _GEN_5735 : dirty_121_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6023 = fence_working ? _GEN_5736 : dirty_122_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6024 = fence_working ? _GEN_5737 : dirty_122_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6025 = fence_working ? _GEN_5738 : dirty_123_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6026 = fence_working ? _GEN_5739 : dirty_123_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6027 = fence_working ? _GEN_5740 : dirty_124_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6028 = fence_working ? _GEN_5741 : dirty_124_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6029 = fence_working ? _GEN_5742 : dirty_125_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6030 = fence_working ? _GEN_5743 : dirty_125_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6031 = fence_working ? _GEN_5744 : dirty_126_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6032 = fence_working ? _GEN_5745 : dirty_126_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6033 = fence_working ? _GEN_5746 : dirty_127_0; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6034 = fence_working ? _GEN_5747 : dirty_127_1; // @[DCache.scala 370:27 69:22]
  wire  _GEN_6035 = fence_working ? _GEN_5748 : 1'h1; // @[DCache.scala 370:27 413:27]
  wire  _GEN_6036 = fence_working ? _GEN_5749 : bram_use_replace_addr; // @[DCache.scala 370:27 95:40]
  wire [2:0] _GEN_6037 = fence_working ? _GEN_5750 : state; // @[DCache.scala 370:27 65:96]
  wire [31:0] _GEN_6056 = _GEN_441 ? cache_data_1 : cache_data_0; // @[DCache.scala 425:{55,55}]
  wire [31:0] _GEN_6039 = 4'h0 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_0; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6040 = 4'h1 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_1; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6041 = 4'h2 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_2; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6042 = 4'h3 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_3; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6043 = 4'h4 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_4; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6044 = 4'h5 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_5; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6045 = 4'h6 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_6; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6046 = 4'h7 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_7; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6047 = 4'h8 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_8; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6048 = 4'h9 == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_9; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6049 = 4'ha == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_10; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6050 = 4'hb == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_11; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6051 = 4'hc == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_12; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6052 = 4'hd == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_13; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6053 = 4'he == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_14; // @[DCache.scala 425:{55,55} 94:40]
  wire [31:0] _GEN_6054 = 4'hf == bram_read_ready_addr[3:0] ? _GEN_6056 : bram_r_buffer_15; // @[DCache.scala 425:{55,55} 94:40]
  wire [19:0] _GEN_6058 = _GEN_441 ? cache_tag_1 : cache_tag_0; // @[Cat.scala 33:{92,92}]
  wire [31:0] _aw_addr_T_1 = {_GEN_6058,io_cpu_M_mem_va[11:6],6'h0}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_6061 = _T_38 ? _aw_addr_T_1 : _GEN_281; // @[DCache.scala 426:33 427:28]
  wire [31:0] _GEN_6065 = _T_38 ? _GEN_6056 : _GEN_283; // @[DCache.scala 426:33 431:28]
  wire [31:0] _w_data_T_13 = _w_data_T_3 ? _GEN_6056 : _GEN_5226; // @[DCache.scala 444:30]
  wire [31:0] _GEN_6091 = w_last ? _GEN_6065 : _w_data_T_13; // @[DCache.scala 441:28 444:24]
  wire [31:0] _GEN_6095 = _T_1 ? _GEN_6091 : _GEN_6065; // @[DCache.scala 440:33]
  wire  _GEN_6098 = _GEN_11687 & _GEN_11689 ? 1'h0 : dirty_0_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6099 = _GEN_11687 & _GEN_441 ? 1'h0 : dirty_0_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6100 = _GEN_11688 & _GEN_11689 ? 1'h0 : dirty_1_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6101 = _GEN_11688 & _GEN_441 ? 1'h0 : dirty_1_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6102 = _GEN_11691 & _GEN_11689 ? 1'h0 : dirty_2_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6103 = _GEN_11691 & _GEN_441 ? 1'h0 : dirty_2_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6104 = _GEN_11694 & _GEN_11689 ? 1'h0 : dirty_3_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6105 = _GEN_11694 & _GEN_441 ? 1'h0 : dirty_3_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6106 = _GEN_11697 & _GEN_11689 ? 1'h0 : dirty_4_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6107 = _GEN_11697 & _GEN_441 ? 1'h0 : dirty_4_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6108 = _GEN_11700 & _GEN_11689 ? 1'h0 : dirty_5_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6109 = _GEN_11700 & _GEN_441 ? 1'h0 : dirty_5_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6110 = _GEN_11703 & _GEN_11689 ? 1'h0 : dirty_6_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6111 = _GEN_11703 & _GEN_441 ? 1'h0 : dirty_6_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6112 = _GEN_11706 & _GEN_11689 ? 1'h0 : dirty_7_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6113 = _GEN_11706 & _GEN_441 ? 1'h0 : dirty_7_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6114 = _GEN_11709 & _GEN_11689 ? 1'h0 : dirty_8_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6115 = _GEN_11709 & _GEN_441 ? 1'h0 : dirty_8_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6116 = _GEN_11712 & _GEN_11689 ? 1'h0 : dirty_9_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6117 = _GEN_11712 & _GEN_441 ? 1'h0 : dirty_9_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6118 = _GEN_11715 & _GEN_11689 ? 1'h0 : dirty_10_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6119 = _GEN_11715 & _GEN_441 ? 1'h0 : dirty_10_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6120 = _GEN_11718 & _GEN_11689 ? 1'h0 : dirty_11_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6121 = _GEN_11718 & _GEN_441 ? 1'h0 : dirty_11_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6122 = _GEN_11721 & _GEN_11689 ? 1'h0 : dirty_12_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6123 = _GEN_11721 & _GEN_441 ? 1'h0 : dirty_12_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6124 = _GEN_11724 & _GEN_11689 ? 1'h0 : dirty_13_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6125 = _GEN_11724 & _GEN_441 ? 1'h0 : dirty_13_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6126 = _GEN_11727 & _GEN_11689 ? 1'h0 : dirty_14_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6127 = _GEN_11727 & _GEN_441 ? 1'h0 : dirty_14_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6128 = _GEN_11730 & _GEN_11689 ? 1'h0 : dirty_15_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6129 = _GEN_11730 & _GEN_441 ? 1'h0 : dirty_15_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6130 = _GEN_11733 & _GEN_11689 ? 1'h0 : dirty_16_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6131 = _GEN_11733 & _GEN_441 ? 1'h0 : dirty_16_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6132 = _GEN_11736 & _GEN_11689 ? 1'h0 : dirty_17_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6133 = _GEN_11736 & _GEN_441 ? 1'h0 : dirty_17_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6134 = _GEN_11739 & _GEN_11689 ? 1'h0 : dirty_18_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6135 = _GEN_11739 & _GEN_441 ? 1'h0 : dirty_18_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6136 = _GEN_11742 & _GEN_11689 ? 1'h0 : dirty_19_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6137 = _GEN_11742 & _GEN_441 ? 1'h0 : dirty_19_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6138 = _GEN_11745 & _GEN_11689 ? 1'h0 : dirty_20_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6139 = _GEN_11745 & _GEN_441 ? 1'h0 : dirty_20_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6140 = _GEN_11748 & _GEN_11689 ? 1'h0 : dirty_21_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6141 = _GEN_11748 & _GEN_441 ? 1'h0 : dirty_21_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6142 = _GEN_11751 & _GEN_11689 ? 1'h0 : dirty_22_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6143 = _GEN_11751 & _GEN_441 ? 1'h0 : dirty_22_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6144 = _GEN_11754 & _GEN_11689 ? 1'h0 : dirty_23_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6145 = _GEN_11754 & _GEN_441 ? 1'h0 : dirty_23_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6146 = _GEN_11757 & _GEN_11689 ? 1'h0 : dirty_24_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6147 = _GEN_11757 & _GEN_441 ? 1'h0 : dirty_24_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6148 = _GEN_11760 & _GEN_11689 ? 1'h0 : dirty_25_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6149 = _GEN_11760 & _GEN_441 ? 1'h0 : dirty_25_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6150 = _GEN_11763 & _GEN_11689 ? 1'h0 : dirty_26_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6151 = _GEN_11763 & _GEN_441 ? 1'h0 : dirty_26_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6152 = _GEN_11766 & _GEN_11689 ? 1'h0 : dirty_27_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6153 = _GEN_11766 & _GEN_441 ? 1'h0 : dirty_27_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6154 = _GEN_11769 & _GEN_11689 ? 1'h0 : dirty_28_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6155 = _GEN_11769 & _GEN_441 ? 1'h0 : dirty_28_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6156 = _GEN_11772 & _GEN_11689 ? 1'h0 : dirty_29_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6157 = _GEN_11772 & _GEN_441 ? 1'h0 : dirty_29_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6158 = _GEN_11775 & _GEN_11689 ? 1'h0 : dirty_30_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6159 = _GEN_11775 & _GEN_441 ? 1'h0 : dirty_30_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6160 = _GEN_11778 & _GEN_11689 ? 1'h0 : dirty_31_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6161 = _GEN_11778 & _GEN_441 ? 1'h0 : dirty_31_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6162 = _GEN_11781 & _GEN_11689 ? 1'h0 : dirty_32_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6163 = _GEN_11781 & _GEN_441 ? 1'h0 : dirty_32_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6164 = _GEN_11784 & _GEN_11689 ? 1'h0 : dirty_33_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6165 = _GEN_11784 & _GEN_441 ? 1'h0 : dirty_33_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6166 = _GEN_11787 & _GEN_11689 ? 1'h0 : dirty_34_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6167 = _GEN_11787 & _GEN_441 ? 1'h0 : dirty_34_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6168 = _GEN_11790 & _GEN_11689 ? 1'h0 : dirty_35_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6169 = _GEN_11790 & _GEN_441 ? 1'h0 : dirty_35_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6170 = _GEN_11793 & _GEN_11689 ? 1'h0 : dirty_36_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6171 = _GEN_11793 & _GEN_441 ? 1'h0 : dirty_36_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6172 = _GEN_11796 & _GEN_11689 ? 1'h0 : dirty_37_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6173 = _GEN_11796 & _GEN_441 ? 1'h0 : dirty_37_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6174 = _GEN_11799 & _GEN_11689 ? 1'h0 : dirty_38_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6175 = _GEN_11799 & _GEN_441 ? 1'h0 : dirty_38_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6176 = _GEN_11802 & _GEN_11689 ? 1'h0 : dirty_39_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6177 = _GEN_11802 & _GEN_441 ? 1'h0 : dirty_39_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6178 = _GEN_11805 & _GEN_11689 ? 1'h0 : dirty_40_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6179 = _GEN_11805 & _GEN_441 ? 1'h0 : dirty_40_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6180 = _GEN_11808 & _GEN_11689 ? 1'h0 : dirty_41_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6181 = _GEN_11808 & _GEN_441 ? 1'h0 : dirty_41_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6182 = _GEN_11811 & _GEN_11689 ? 1'h0 : dirty_42_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6183 = _GEN_11811 & _GEN_441 ? 1'h0 : dirty_42_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6184 = _GEN_11814 & _GEN_11689 ? 1'h0 : dirty_43_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6185 = _GEN_11814 & _GEN_441 ? 1'h0 : dirty_43_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6186 = _GEN_11817 & _GEN_11689 ? 1'h0 : dirty_44_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6187 = _GEN_11817 & _GEN_441 ? 1'h0 : dirty_44_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6188 = _GEN_11820 & _GEN_11689 ? 1'h0 : dirty_45_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6189 = _GEN_11820 & _GEN_441 ? 1'h0 : dirty_45_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6190 = _GEN_11823 & _GEN_11689 ? 1'h0 : dirty_46_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6191 = _GEN_11823 & _GEN_441 ? 1'h0 : dirty_46_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6192 = _GEN_11826 & _GEN_11689 ? 1'h0 : dirty_47_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6193 = _GEN_11826 & _GEN_441 ? 1'h0 : dirty_47_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6194 = _GEN_11829 & _GEN_11689 ? 1'h0 : dirty_48_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6195 = _GEN_11829 & _GEN_441 ? 1'h0 : dirty_48_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6196 = _GEN_11832 & _GEN_11689 ? 1'h0 : dirty_49_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6197 = _GEN_11832 & _GEN_441 ? 1'h0 : dirty_49_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6198 = _GEN_11835 & _GEN_11689 ? 1'h0 : dirty_50_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6199 = _GEN_11835 & _GEN_441 ? 1'h0 : dirty_50_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6200 = _GEN_11838 & _GEN_11689 ? 1'h0 : dirty_51_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6201 = _GEN_11838 & _GEN_441 ? 1'h0 : dirty_51_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6202 = _GEN_11841 & _GEN_11689 ? 1'h0 : dirty_52_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6203 = _GEN_11841 & _GEN_441 ? 1'h0 : dirty_52_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6204 = _GEN_11844 & _GEN_11689 ? 1'h0 : dirty_53_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6205 = _GEN_11844 & _GEN_441 ? 1'h0 : dirty_53_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6206 = _GEN_11847 & _GEN_11689 ? 1'h0 : dirty_54_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6207 = _GEN_11847 & _GEN_441 ? 1'h0 : dirty_54_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6208 = _GEN_11850 & _GEN_11689 ? 1'h0 : dirty_55_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6209 = _GEN_11850 & _GEN_441 ? 1'h0 : dirty_55_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6210 = _GEN_11853 & _GEN_11689 ? 1'h0 : dirty_56_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6211 = _GEN_11853 & _GEN_441 ? 1'h0 : dirty_56_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6212 = _GEN_11856 & _GEN_11689 ? 1'h0 : dirty_57_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6213 = _GEN_11856 & _GEN_441 ? 1'h0 : dirty_57_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6214 = _GEN_11859 & _GEN_11689 ? 1'h0 : dirty_58_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6215 = _GEN_11859 & _GEN_441 ? 1'h0 : dirty_58_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6216 = _GEN_11862 & _GEN_11689 ? 1'h0 : dirty_59_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6217 = _GEN_11862 & _GEN_441 ? 1'h0 : dirty_59_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6218 = _GEN_11865 & _GEN_11689 ? 1'h0 : dirty_60_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6219 = _GEN_11865 & _GEN_441 ? 1'h0 : dirty_60_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6220 = _GEN_11868 & _GEN_11689 ? 1'h0 : dirty_61_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6221 = _GEN_11868 & _GEN_441 ? 1'h0 : dirty_61_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6222 = _GEN_11871 & _GEN_11689 ? 1'h0 : dirty_62_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6223 = _GEN_11871 & _GEN_441 ? 1'h0 : dirty_62_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6224 = _GEN_11874 & _GEN_11689 ? 1'h0 : dirty_63_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6225 = _GEN_11874 & _GEN_441 ? 1'h0 : dirty_63_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6226 = _GEN_11878 & _GEN_11689 ? 1'h0 : dirty_64_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6227 = _GEN_11878 & _GEN_441 ? 1'h0 : dirty_64_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6228 = _GEN_11883 & _GEN_11689 ? 1'h0 : dirty_65_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6229 = _GEN_11883 & _GEN_441 ? 1'h0 : dirty_65_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6230 = _GEN_11888 & _GEN_11689 ? 1'h0 : dirty_66_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6231 = _GEN_11888 & _GEN_441 ? 1'h0 : dirty_66_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6232 = _GEN_11893 & _GEN_11689 ? 1'h0 : dirty_67_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6233 = _GEN_11893 & _GEN_441 ? 1'h0 : dirty_67_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6234 = _GEN_11898 & _GEN_11689 ? 1'h0 : dirty_68_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6235 = _GEN_11898 & _GEN_441 ? 1'h0 : dirty_68_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6236 = _GEN_11903 & _GEN_11689 ? 1'h0 : dirty_69_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6237 = _GEN_11903 & _GEN_441 ? 1'h0 : dirty_69_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6238 = _GEN_11908 & _GEN_11689 ? 1'h0 : dirty_70_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6239 = _GEN_11908 & _GEN_441 ? 1'h0 : dirty_70_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6240 = _GEN_11913 & _GEN_11689 ? 1'h0 : dirty_71_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6241 = _GEN_11913 & _GEN_441 ? 1'h0 : dirty_71_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6242 = _GEN_11918 & _GEN_11689 ? 1'h0 : dirty_72_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6243 = _GEN_11918 & _GEN_441 ? 1'h0 : dirty_72_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6244 = _GEN_11923 & _GEN_11689 ? 1'h0 : dirty_73_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6245 = _GEN_11923 & _GEN_441 ? 1'h0 : dirty_73_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6246 = _GEN_11928 & _GEN_11689 ? 1'h0 : dirty_74_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6247 = _GEN_11928 & _GEN_441 ? 1'h0 : dirty_74_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6248 = _GEN_11933 & _GEN_11689 ? 1'h0 : dirty_75_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6249 = _GEN_11933 & _GEN_441 ? 1'h0 : dirty_75_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6250 = _GEN_11938 & _GEN_11689 ? 1'h0 : dirty_76_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6251 = _GEN_11938 & _GEN_441 ? 1'h0 : dirty_76_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6252 = _GEN_11943 & _GEN_11689 ? 1'h0 : dirty_77_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6253 = _GEN_11943 & _GEN_441 ? 1'h0 : dirty_77_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6254 = _GEN_11948 & _GEN_11689 ? 1'h0 : dirty_78_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6255 = _GEN_11948 & _GEN_441 ? 1'h0 : dirty_78_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6256 = _GEN_11953 & _GEN_11689 ? 1'h0 : dirty_79_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6257 = _GEN_11953 & _GEN_441 ? 1'h0 : dirty_79_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6258 = _GEN_11958 & _GEN_11689 ? 1'h0 : dirty_80_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6259 = _GEN_11958 & _GEN_441 ? 1'h0 : dirty_80_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6260 = _GEN_11963 & _GEN_11689 ? 1'h0 : dirty_81_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6261 = _GEN_11963 & _GEN_441 ? 1'h0 : dirty_81_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6262 = _GEN_11968 & _GEN_11689 ? 1'h0 : dirty_82_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6263 = _GEN_11968 & _GEN_441 ? 1'h0 : dirty_82_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6264 = _GEN_11973 & _GEN_11689 ? 1'h0 : dirty_83_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6265 = _GEN_11973 & _GEN_441 ? 1'h0 : dirty_83_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6266 = _GEN_11978 & _GEN_11689 ? 1'h0 : dirty_84_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6267 = _GEN_11978 & _GEN_441 ? 1'h0 : dirty_84_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6268 = _GEN_11983 & _GEN_11689 ? 1'h0 : dirty_85_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6269 = _GEN_11983 & _GEN_441 ? 1'h0 : dirty_85_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6270 = _GEN_11988 & _GEN_11689 ? 1'h0 : dirty_86_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6271 = _GEN_11988 & _GEN_441 ? 1'h0 : dirty_86_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6272 = _GEN_11993 & _GEN_11689 ? 1'h0 : dirty_87_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6273 = _GEN_11993 & _GEN_441 ? 1'h0 : dirty_87_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6274 = _GEN_11998 & _GEN_11689 ? 1'h0 : dirty_88_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6275 = _GEN_11998 & _GEN_441 ? 1'h0 : dirty_88_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6276 = _GEN_12003 & _GEN_11689 ? 1'h0 : dirty_89_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6277 = _GEN_12003 & _GEN_441 ? 1'h0 : dirty_89_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6278 = _GEN_12008 & _GEN_11689 ? 1'h0 : dirty_90_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6279 = _GEN_12008 & _GEN_441 ? 1'h0 : dirty_90_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6280 = _GEN_12013 & _GEN_11689 ? 1'h0 : dirty_91_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6281 = _GEN_12013 & _GEN_441 ? 1'h0 : dirty_91_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6282 = _GEN_12018 & _GEN_11689 ? 1'h0 : dirty_92_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6283 = _GEN_12018 & _GEN_441 ? 1'h0 : dirty_92_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6284 = _GEN_12023 & _GEN_11689 ? 1'h0 : dirty_93_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6285 = _GEN_12023 & _GEN_441 ? 1'h0 : dirty_93_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6286 = _GEN_12028 & _GEN_11689 ? 1'h0 : dirty_94_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6287 = _GEN_12028 & _GEN_441 ? 1'h0 : dirty_94_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6288 = _GEN_12033 & _GEN_11689 ? 1'h0 : dirty_95_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6289 = _GEN_12033 & _GEN_441 ? 1'h0 : dirty_95_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6290 = _GEN_12038 & _GEN_11689 ? 1'h0 : dirty_96_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6291 = _GEN_12038 & _GEN_441 ? 1'h0 : dirty_96_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6292 = _GEN_12043 & _GEN_11689 ? 1'h0 : dirty_97_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6293 = _GEN_12043 & _GEN_441 ? 1'h0 : dirty_97_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6294 = _GEN_12048 & _GEN_11689 ? 1'h0 : dirty_98_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6295 = _GEN_12048 & _GEN_441 ? 1'h0 : dirty_98_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6296 = _GEN_12053 & _GEN_11689 ? 1'h0 : dirty_99_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6297 = _GEN_12053 & _GEN_441 ? 1'h0 : dirty_99_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6298 = _GEN_12058 & _GEN_11689 ? 1'h0 : dirty_100_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6299 = _GEN_12058 & _GEN_441 ? 1'h0 : dirty_100_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6300 = _GEN_12063 & _GEN_11689 ? 1'h0 : dirty_101_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6301 = _GEN_12063 & _GEN_441 ? 1'h0 : dirty_101_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6302 = _GEN_12068 & _GEN_11689 ? 1'h0 : dirty_102_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6303 = _GEN_12068 & _GEN_441 ? 1'h0 : dirty_102_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6304 = _GEN_12073 & _GEN_11689 ? 1'h0 : dirty_103_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6305 = _GEN_12073 & _GEN_441 ? 1'h0 : dirty_103_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6306 = _GEN_12078 & _GEN_11689 ? 1'h0 : dirty_104_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6307 = _GEN_12078 & _GEN_441 ? 1'h0 : dirty_104_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6308 = _GEN_12083 & _GEN_11689 ? 1'h0 : dirty_105_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6309 = _GEN_12083 & _GEN_441 ? 1'h0 : dirty_105_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6310 = _GEN_12088 & _GEN_11689 ? 1'h0 : dirty_106_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6311 = _GEN_12088 & _GEN_441 ? 1'h0 : dirty_106_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6312 = _GEN_12093 & _GEN_11689 ? 1'h0 : dirty_107_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6313 = _GEN_12093 & _GEN_441 ? 1'h0 : dirty_107_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6314 = _GEN_12098 & _GEN_11689 ? 1'h0 : dirty_108_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6315 = _GEN_12098 & _GEN_441 ? 1'h0 : dirty_108_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6316 = _GEN_12103 & _GEN_11689 ? 1'h0 : dirty_109_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6317 = _GEN_12103 & _GEN_441 ? 1'h0 : dirty_109_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6318 = _GEN_12108 & _GEN_11689 ? 1'h0 : dirty_110_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6319 = _GEN_12108 & _GEN_441 ? 1'h0 : dirty_110_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6320 = _GEN_12113 & _GEN_11689 ? 1'h0 : dirty_111_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6321 = _GEN_12113 & _GEN_441 ? 1'h0 : dirty_111_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6322 = _GEN_12118 & _GEN_11689 ? 1'h0 : dirty_112_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6323 = _GEN_12118 & _GEN_441 ? 1'h0 : dirty_112_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6324 = _GEN_12123 & _GEN_11689 ? 1'h0 : dirty_113_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6325 = _GEN_12123 & _GEN_441 ? 1'h0 : dirty_113_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6326 = _GEN_12128 & _GEN_11689 ? 1'h0 : dirty_114_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6327 = _GEN_12128 & _GEN_441 ? 1'h0 : dirty_114_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6328 = _GEN_12133 & _GEN_11689 ? 1'h0 : dirty_115_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6329 = _GEN_12133 & _GEN_441 ? 1'h0 : dirty_115_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6330 = _GEN_12138 & _GEN_11689 ? 1'h0 : dirty_116_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6331 = _GEN_12138 & _GEN_441 ? 1'h0 : dirty_116_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6332 = _GEN_12143 & _GEN_11689 ? 1'h0 : dirty_117_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6333 = _GEN_12143 & _GEN_441 ? 1'h0 : dirty_117_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6334 = _GEN_12148 & _GEN_11689 ? 1'h0 : dirty_118_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6335 = _GEN_12148 & _GEN_441 ? 1'h0 : dirty_118_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6336 = _GEN_12153 & _GEN_11689 ? 1'h0 : dirty_119_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6337 = _GEN_12153 & _GEN_441 ? 1'h0 : dirty_119_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6338 = _GEN_12158 & _GEN_11689 ? 1'h0 : dirty_120_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6339 = _GEN_12158 & _GEN_441 ? 1'h0 : dirty_120_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6340 = _GEN_12163 & _GEN_11689 ? 1'h0 : dirty_121_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6341 = _GEN_12163 & _GEN_441 ? 1'h0 : dirty_121_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6342 = _GEN_12168 & _GEN_11689 ? 1'h0 : dirty_122_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6343 = _GEN_12168 & _GEN_441 ? 1'h0 : dirty_122_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6344 = _GEN_12173 & _GEN_11689 ? 1'h0 : dirty_123_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6345 = _GEN_12173 & _GEN_441 ? 1'h0 : dirty_123_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6346 = _GEN_12178 & _GEN_11689 ? 1'h0 : dirty_124_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6347 = _GEN_12178 & _GEN_441 ? 1'h0 : dirty_124_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6348 = _GEN_12183 & _GEN_11689 ? 1'h0 : dirty_125_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6349 = _GEN_12183 & _GEN_441 ? 1'h0 : dirty_125_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6350 = _GEN_12188 & _GEN_11689 ? 1'h0 : dirty_126_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6351 = _GEN_12188 & _GEN_441 ? 1'h0 : dirty_126_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6352 = _GEN_12193 & _GEN_11689 ? 1'h0 : dirty_127_0; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6353 = _GEN_12193 & _GEN_441 ? 1'h0 : dirty_127_1; // @[DCache.scala 456:{54,54} 69:22]
  wire  _GEN_6354 = io_axi_b_valid ? _GEN_6098 : dirty_0_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6355 = io_axi_b_valid ? _GEN_6099 : dirty_0_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6356 = io_axi_b_valid ? _GEN_6100 : dirty_1_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6357 = io_axi_b_valid ? _GEN_6101 : dirty_1_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6358 = io_axi_b_valid ? _GEN_6102 : dirty_2_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6359 = io_axi_b_valid ? _GEN_6103 : dirty_2_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6360 = io_axi_b_valid ? _GEN_6104 : dirty_3_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6361 = io_axi_b_valid ? _GEN_6105 : dirty_3_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6362 = io_axi_b_valid ? _GEN_6106 : dirty_4_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6363 = io_axi_b_valid ? _GEN_6107 : dirty_4_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6364 = io_axi_b_valid ? _GEN_6108 : dirty_5_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6365 = io_axi_b_valid ? _GEN_6109 : dirty_5_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6366 = io_axi_b_valid ? _GEN_6110 : dirty_6_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6367 = io_axi_b_valid ? _GEN_6111 : dirty_6_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6368 = io_axi_b_valid ? _GEN_6112 : dirty_7_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6369 = io_axi_b_valid ? _GEN_6113 : dirty_7_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6370 = io_axi_b_valid ? _GEN_6114 : dirty_8_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6371 = io_axi_b_valid ? _GEN_6115 : dirty_8_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6372 = io_axi_b_valid ? _GEN_6116 : dirty_9_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6373 = io_axi_b_valid ? _GEN_6117 : dirty_9_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6374 = io_axi_b_valid ? _GEN_6118 : dirty_10_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6375 = io_axi_b_valid ? _GEN_6119 : dirty_10_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6376 = io_axi_b_valid ? _GEN_6120 : dirty_11_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6377 = io_axi_b_valid ? _GEN_6121 : dirty_11_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6378 = io_axi_b_valid ? _GEN_6122 : dirty_12_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6379 = io_axi_b_valid ? _GEN_6123 : dirty_12_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6380 = io_axi_b_valid ? _GEN_6124 : dirty_13_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6381 = io_axi_b_valid ? _GEN_6125 : dirty_13_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6382 = io_axi_b_valid ? _GEN_6126 : dirty_14_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6383 = io_axi_b_valid ? _GEN_6127 : dirty_14_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6384 = io_axi_b_valid ? _GEN_6128 : dirty_15_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6385 = io_axi_b_valid ? _GEN_6129 : dirty_15_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6386 = io_axi_b_valid ? _GEN_6130 : dirty_16_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6387 = io_axi_b_valid ? _GEN_6131 : dirty_16_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6388 = io_axi_b_valid ? _GEN_6132 : dirty_17_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6389 = io_axi_b_valid ? _GEN_6133 : dirty_17_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6390 = io_axi_b_valid ? _GEN_6134 : dirty_18_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6391 = io_axi_b_valid ? _GEN_6135 : dirty_18_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6392 = io_axi_b_valid ? _GEN_6136 : dirty_19_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6393 = io_axi_b_valid ? _GEN_6137 : dirty_19_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6394 = io_axi_b_valid ? _GEN_6138 : dirty_20_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6395 = io_axi_b_valid ? _GEN_6139 : dirty_20_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6396 = io_axi_b_valid ? _GEN_6140 : dirty_21_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6397 = io_axi_b_valid ? _GEN_6141 : dirty_21_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6398 = io_axi_b_valid ? _GEN_6142 : dirty_22_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6399 = io_axi_b_valid ? _GEN_6143 : dirty_22_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6400 = io_axi_b_valid ? _GEN_6144 : dirty_23_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6401 = io_axi_b_valid ? _GEN_6145 : dirty_23_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6402 = io_axi_b_valid ? _GEN_6146 : dirty_24_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6403 = io_axi_b_valid ? _GEN_6147 : dirty_24_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6404 = io_axi_b_valid ? _GEN_6148 : dirty_25_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6405 = io_axi_b_valid ? _GEN_6149 : dirty_25_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6406 = io_axi_b_valid ? _GEN_6150 : dirty_26_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6407 = io_axi_b_valid ? _GEN_6151 : dirty_26_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6408 = io_axi_b_valid ? _GEN_6152 : dirty_27_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6409 = io_axi_b_valid ? _GEN_6153 : dirty_27_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6410 = io_axi_b_valid ? _GEN_6154 : dirty_28_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6411 = io_axi_b_valid ? _GEN_6155 : dirty_28_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6412 = io_axi_b_valid ? _GEN_6156 : dirty_29_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6413 = io_axi_b_valid ? _GEN_6157 : dirty_29_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6414 = io_axi_b_valid ? _GEN_6158 : dirty_30_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6415 = io_axi_b_valid ? _GEN_6159 : dirty_30_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6416 = io_axi_b_valid ? _GEN_6160 : dirty_31_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6417 = io_axi_b_valid ? _GEN_6161 : dirty_31_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6418 = io_axi_b_valid ? _GEN_6162 : dirty_32_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6419 = io_axi_b_valid ? _GEN_6163 : dirty_32_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6420 = io_axi_b_valid ? _GEN_6164 : dirty_33_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6421 = io_axi_b_valid ? _GEN_6165 : dirty_33_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6422 = io_axi_b_valid ? _GEN_6166 : dirty_34_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6423 = io_axi_b_valid ? _GEN_6167 : dirty_34_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6424 = io_axi_b_valid ? _GEN_6168 : dirty_35_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6425 = io_axi_b_valid ? _GEN_6169 : dirty_35_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6426 = io_axi_b_valid ? _GEN_6170 : dirty_36_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6427 = io_axi_b_valid ? _GEN_6171 : dirty_36_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6428 = io_axi_b_valid ? _GEN_6172 : dirty_37_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6429 = io_axi_b_valid ? _GEN_6173 : dirty_37_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6430 = io_axi_b_valid ? _GEN_6174 : dirty_38_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6431 = io_axi_b_valid ? _GEN_6175 : dirty_38_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6432 = io_axi_b_valid ? _GEN_6176 : dirty_39_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6433 = io_axi_b_valid ? _GEN_6177 : dirty_39_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6434 = io_axi_b_valid ? _GEN_6178 : dirty_40_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6435 = io_axi_b_valid ? _GEN_6179 : dirty_40_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6436 = io_axi_b_valid ? _GEN_6180 : dirty_41_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6437 = io_axi_b_valid ? _GEN_6181 : dirty_41_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6438 = io_axi_b_valid ? _GEN_6182 : dirty_42_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6439 = io_axi_b_valid ? _GEN_6183 : dirty_42_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6440 = io_axi_b_valid ? _GEN_6184 : dirty_43_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6441 = io_axi_b_valid ? _GEN_6185 : dirty_43_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6442 = io_axi_b_valid ? _GEN_6186 : dirty_44_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6443 = io_axi_b_valid ? _GEN_6187 : dirty_44_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6444 = io_axi_b_valid ? _GEN_6188 : dirty_45_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6445 = io_axi_b_valid ? _GEN_6189 : dirty_45_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6446 = io_axi_b_valid ? _GEN_6190 : dirty_46_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6447 = io_axi_b_valid ? _GEN_6191 : dirty_46_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6448 = io_axi_b_valid ? _GEN_6192 : dirty_47_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6449 = io_axi_b_valid ? _GEN_6193 : dirty_47_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6450 = io_axi_b_valid ? _GEN_6194 : dirty_48_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6451 = io_axi_b_valid ? _GEN_6195 : dirty_48_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6452 = io_axi_b_valid ? _GEN_6196 : dirty_49_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6453 = io_axi_b_valid ? _GEN_6197 : dirty_49_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6454 = io_axi_b_valid ? _GEN_6198 : dirty_50_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6455 = io_axi_b_valid ? _GEN_6199 : dirty_50_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6456 = io_axi_b_valid ? _GEN_6200 : dirty_51_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6457 = io_axi_b_valid ? _GEN_6201 : dirty_51_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6458 = io_axi_b_valid ? _GEN_6202 : dirty_52_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6459 = io_axi_b_valid ? _GEN_6203 : dirty_52_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6460 = io_axi_b_valid ? _GEN_6204 : dirty_53_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6461 = io_axi_b_valid ? _GEN_6205 : dirty_53_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6462 = io_axi_b_valid ? _GEN_6206 : dirty_54_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6463 = io_axi_b_valid ? _GEN_6207 : dirty_54_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6464 = io_axi_b_valid ? _GEN_6208 : dirty_55_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6465 = io_axi_b_valid ? _GEN_6209 : dirty_55_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6466 = io_axi_b_valid ? _GEN_6210 : dirty_56_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6467 = io_axi_b_valid ? _GEN_6211 : dirty_56_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6468 = io_axi_b_valid ? _GEN_6212 : dirty_57_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6469 = io_axi_b_valid ? _GEN_6213 : dirty_57_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6470 = io_axi_b_valid ? _GEN_6214 : dirty_58_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6471 = io_axi_b_valid ? _GEN_6215 : dirty_58_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6472 = io_axi_b_valid ? _GEN_6216 : dirty_59_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6473 = io_axi_b_valid ? _GEN_6217 : dirty_59_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6474 = io_axi_b_valid ? _GEN_6218 : dirty_60_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6475 = io_axi_b_valid ? _GEN_6219 : dirty_60_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6476 = io_axi_b_valid ? _GEN_6220 : dirty_61_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6477 = io_axi_b_valid ? _GEN_6221 : dirty_61_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6478 = io_axi_b_valid ? _GEN_6222 : dirty_62_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6479 = io_axi_b_valid ? _GEN_6223 : dirty_62_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6480 = io_axi_b_valid ? _GEN_6224 : dirty_63_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6481 = io_axi_b_valid ? _GEN_6225 : dirty_63_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6482 = io_axi_b_valid ? _GEN_6226 : dirty_64_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6483 = io_axi_b_valid ? _GEN_6227 : dirty_64_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6484 = io_axi_b_valid ? _GEN_6228 : dirty_65_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6485 = io_axi_b_valid ? _GEN_6229 : dirty_65_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6486 = io_axi_b_valid ? _GEN_6230 : dirty_66_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6487 = io_axi_b_valid ? _GEN_6231 : dirty_66_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6488 = io_axi_b_valid ? _GEN_6232 : dirty_67_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6489 = io_axi_b_valid ? _GEN_6233 : dirty_67_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6490 = io_axi_b_valid ? _GEN_6234 : dirty_68_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6491 = io_axi_b_valid ? _GEN_6235 : dirty_68_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6492 = io_axi_b_valid ? _GEN_6236 : dirty_69_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6493 = io_axi_b_valid ? _GEN_6237 : dirty_69_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6494 = io_axi_b_valid ? _GEN_6238 : dirty_70_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6495 = io_axi_b_valid ? _GEN_6239 : dirty_70_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6496 = io_axi_b_valid ? _GEN_6240 : dirty_71_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6497 = io_axi_b_valid ? _GEN_6241 : dirty_71_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6498 = io_axi_b_valid ? _GEN_6242 : dirty_72_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6499 = io_axi_b_valid ? _GEN_6243 : dirty_72_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6500 = io_axi_b_valid ? _GEN_6244 : dirty_73_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6501 = io_axi_b_valid ? _GEN_6245 : dirty_73_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6502 = io_axi_b_valid ? _GEN_6246 : dirty_74_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6503 = io_axi_b_valid ? _GEN_6247 : dirty_74_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6504 = io_axi_b_valid ? _GEN_6248 : dirty_75_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6505 = io_axi_b_valid ? _GEN_6249 : dirty_75_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6506 = io_axi_b_valid ? _GEN_6250 : dirty_76_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6507 = io_axi_b_valid ? _GEN_6251 : dirty_76_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6508 = io_axi_b_valid ? _GEN_6252 : dirty_77_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6509 = io_axi_b_valid ? _GEN_6253 : dirty_77_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6510 = io_axi_b_valid ? _GEN_6254 : dirty_78_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6511 = io_axi_b_valid ? _GEN_6255 : dirty_78_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6512 = io_axi_b_valid ? _GEN_6256 : dirty_79_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6513 = io_axi_b_valid ? _GEN_6257 : dirty_79_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6514 = io_axi_b_valid ? _GEN_6258 : dirty_80_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6515 = io_axi_b_valid ? _GEN_6259 : dirty_80_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6516 = io_axi_b_valid ? _GEN_6260 : dirty_81_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6517 = io_axi_b_valid ? _GEN_6261 : dirty_81_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6518 = io_axi_b_valid ? _GEN_6262 : dirty_82_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6519 = io_axi_b_valid ? _GEN_6263 : dirty_82_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6520 = io_axi_b_valid ? _GEN_6264 : dirty_83_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6521 = io_axi_b_valid ? _GEN_6265 : dirty_83_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6522 = io_axi_b_valid ? _GEN_6266 : dirty_84_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6523 = io_axi_b_valid ? _GEN_6267 : dirty_84_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6524 = io_axi_b_valid ? _GEN_6268 : dirty_85_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6525 = io_axi_b_valid ? _GEN_6269 : dirty_85_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6526 = io_axi_b_valid ? _GEN_6270 : dirty_86_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6527 = io_axi_b_valid ? _GEN_6271 : dirty_86_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6528 = io_axi_b_valid ? _GEN_6272 : dirty_87_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6529 = io_axi_b_valid ? _GEN_6273 : dirty_87_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6530 = io_axi_b_valid ? _GEN_6274 : dirty_88_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6531 = io_axi_b_valid ? _GEN_6275 : dirty_88_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6532 = io_axi_b_valid ? _GEN_6276 : dirty_89_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6533 = io_axi_b_valid ? _GEN_6277 : dirty_89_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6534 = io_axi_b_valid ? _GEN_6278 : dirty_90_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6535 = io_axi_b_valid ? _GEN_6279 : dirty_90_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6536 = io_axi_b_valid ? _GEN_6280 : dirty_91_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6537 = io_axi_b_valid ? _GEN_6281 : dirty_91_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6538 = io_axi_b_valid ? _GEN_6282 : dirty_92_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6539 = io_axi_b_valid ? _GEN_6283 : dirty_92_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6540 = io_axi_b_valid ? _GEN_6284 : dirty_93_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6541 = io_axi_b_valid ? _GEN_6285 : dirty_93_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6542 = io_axi_b_valid ? _GEN_6286 : dirty_94_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6543 = io_axi_b_valid ? _GEN_6287 : dirty_94_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6544 = io_axi_b_valid ? _GEN_6288 : dirty_95_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6545 = io_axi_b_valid ? _GEN_6289 : dirty_95_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6546 = io_axi_b_valid ? _GEN_6290 : dirty_96_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6547 = io_axi_b_valid ? _GEN_6291 : dirty_96_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6548 = io_axi_b_valid ? _GEN_6292 : dirty_97_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6549 = io_axi_b_valid ? _GEN_6293 : dirty_97_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6550 = io_axi_b_valid ? _GEN_6294 : dirty_98_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6551 = io_axi_b_valid ? _GEN_6295 : dirty_98_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6552 = io_axi_b_valid ? _GEN_6296 : dirty_99_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6553 = io_axi_b_valid ? _GEN_6297 : dirty_99_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6554 = io_axi_b_valid ? _GEN_6298 : dirty_100_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6555 = io_axi_b_valid ? _GEN_6299 : dirty_100_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6556 = io_axi_b_valid ? _GEN_6300 : dirty_101_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6557 = io_axi_b_valid ? _GEN_6301 : dirty_101_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6558 = io_axi_b_valid ? _GEN_6302 : dirty_102_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6559 = io_axi_b_valid ? _GEN_6303 : dirty_102_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6560 = io_axi_b_valid ? _GEN_6304 : dirty_103_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6561 = io_axi_b_valid ? _GEN_6305 : dirty_103_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6562 = io_axi_b_valid ? _GEN_6306 : dirty_104_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6563 = io_axi_b_valid ? _GEN_6307 : dirty_104_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6564 = io_axi_b_valid ? _GEN_6308 : dirty_105_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6565 = io_axi_b_valid ? _GEN_6309 : dirty_105_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6566 = io_axi_b_valid ? _GEN_6310 : dirty_106_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6567 = io_axi_b_valid ? _GEN_6311 : dirty_106_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6568 = io_axi_b_valid ? _GEN_6312 : dirty_107_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6569 = io_axi_b_valid ? _GEN_6313 : dirty_107_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6570 = io_axi_b_valid ? _GEN_6314 : dirty_108_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6571 = io_axi_b_valid ? _GEN_6315 : dirty_108_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6572 = io_axi_b_valid ? _GEN_6316 : dirty_109_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6573 = io_axi_b_valid ? _GEN_6317 : dirty_109_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6574 = io_axi_b_valid ? _GEN_6318 : dirty_110_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6575 = io_axi_b_valid ? _GEN_6319 : dirty_110_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6576 = io_axi_b_valid ? _GEN_6320 : dirty_111_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6577 = io_axi_b_valid ? _GEN_6321 : dirty_111_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6578 = io_axi_b_valid ? _GEN_6322 : dirty_112_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6579 = io_axi_b_valid ? _GEN_6323 : dirty_112_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6580 = io_axi_b_valid ? _GEN_6324 : dirty_113_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6581 = io_axi_b_valid ? _GEN_6325 : dirty_113_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6582 = io_axi_b_valid ? _GEN_6326 : dirty_114_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6583 = io_axi_b_valid ? _GEN_6327 : dirty_114_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6584 = io_axi_b_valid ? _GEN_6328 : dirty_115_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6585 = io_axi_b_valid ? _GEN_6329 : dirty_115_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6586 = io_axi_b_valid ? _GEN_6330 : dirty_116_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6587 = io_axi_b_valid ? _GEN_6331 : dirty_116_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6588 = io_axi_b_valid ? _GEN_6332 : dirty_117_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6589 = io_axi_b_valid ? _GEN_6333 : dirty_117_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6590 = io_axi_b_valid ? _GEN_6334 : dirty_118_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6591 = io_axi_b_valid ? _GEN_6335 : dirty_118_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6592 = io_axi_b_valid ? _GEN_6336 : dirty_119_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6593 = io_axi_b_valid ? _GEN_6337 : dirty_119_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6594 = io_axi_b_valid ? _GEN_6338 : dirty_120_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6595 = io_axi_b_valid ? _GEN_6339 : dirty_120_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6596 = io_axi_b_valid ? _GEN_6340 : dirty_121_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6597 = io_axi_b_valid ? _GEN_6341 : dirty_121_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6598 = io_axi_b_valid ? _GEN_6342 : dirty_122_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6599 = io_axi_b_valid ? _GEN_6343 : dirty_122_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6600 = io_axi_b_valid ? _GEN_6344 : dirty_123_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6601 = io_axi_b_valid ? _GEN_6345 : dirty_123_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6602 = io_axi_b_valid ? _GEN_6346 : dirty_124_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6603 = io_axi_b_valid ? _GEN_6347 : dirty_124_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6604 = io_axi_b_valid ? _GEN_6348 : dirty_125_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6605 = io_axi_b_valid ? _GEN_6349 : dirty_125_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6606 = io_axi_b_valid ? _GEN_6350 : dirty_126_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6607 = io_axi_b_valid ? _GEN_6351 : dirty_126_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6608 = io_axi_b_valid ? _GEN_6352 : dirty_127_0; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6609 = io_axi_b_valid ? _GEN_6353 : dirty_127_1; // @[DCache.scala 455:34 69:22]
  wire  _GEN_6610 = io_axi_b_valid ? 1'h0 : replace_writeback; // @[DCache.scala 455:34 101:40 457:54]
  wire [9:0] _GEN_6611 = replace_writeback ? _GEN_5176 : bram_replace_addr; // @[DCache.scala 420:35 90:40]
  wire [9:0] _GEN_6612 = replace_writeback ? bram_replace_addr : bram_read_ready_addr; // @[DCache.scala 420:35 424:55 91:40]
  wire [31:0] _GEN_6613 = replace_writeback ? _GEN_6039 : bram_r_buffer_0; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6614 = replace_writeback ? _GEN_6040 : bram_r_buffer_1; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6615 = replace_writeback ? _GEN_6041 : bram_r_buffer_2; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6616 = replace_writeback ? _GEN_6042 : bram_r_buffer_3; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6617 = replace_writeback ? _GEN_6043 : bram_r_buffer_4; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6618 = replace_writeback ? _GEN_6044 : bram_r_buffer_5; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6619 = replace_writeback ? _GEN_6045 : bram_r_buffer_6; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6620 = replace_writeback ? _GEN_6046 : bram_r_buffer_7; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6621 = replace_writeback ? _GEN_6047 : bram_r_buffer_8; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6622 = replace_writeback ? _GEN_6048 : bram_r_buffer_9; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6623 = replace_writeback ? _GEN_6049 : bram_r_buffer_10; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6624 = replace_writeback ? _GEN_6050 : bram_r_buffer_11; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6625 = replace_writeback ? _GEN_6051 : bram_r_buffer_12; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6626 = replace_writeback ? _GEN_6052 : bram_r_buffer_13; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6627 = replace_writeback ? _GEN_6053 : bram_r_buffer_14; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6628 = replace_writeback ? _GEN_6054 : bram_r_buffer_15; // @[DCache.scala 420:35 94:40]
  wire [31:0] _GEN_6629 = replace_writeback ? _GEN_6061 : _GEN_281; // @[DCache.scala 420:35]
  wire [7:0] _GEN_6630 = replace_writeback ? _GEN_5200 : _GEN_285; // @[DCache.scala 420:35]
  wire [2:0] _GEN_6631 = replace_writeback ? _GEN_5201 : _GEN_282; // @[DCache.scala 420:35]
  wire  _GEN_6632 = replace_writeback ? _GEN_5208 : _GEN_276; // @[DCache.scala 420:35]
  wire [31:0] _GEN_6633 = replace_writeback ? _GEN_6095 : _GEN_283; // @[DCache.scala 420:35]
  wire [3:0] _GEN_6634 = replace_writeback ? _GEN_5204 : _GEN_284; // @[DCache.scala 420:35]
  wire  _GEN_6635 = replace_writeback ? _GEN_5235 : _GEN_278; // @[DCache.scala 420:35]
  wire  _GEN_6636 = replace_writeback ? _GEN_5232 : _GEN_277; // @[DCache.scala 420:35]
  wire  _GEN_6637 = replace_writeback ? _GEN_5207 : aw_handshake; // @[DCache.scala 420:35 100:40]
  wire [3:0] _GEN_6638 = replace_writeback ? _GEN_5234 : axi_wcnt; // @[DCache.scala 420:35 89:40]
  wire  _GEN_6639 = replace_writeback ? _GEN_6354 : dirty_0_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6640 = replace_writeback ? _GEN_6355 : dirty_0_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6641 = replace_writeback ? _GEN_6356 : dirty_1_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6642 = replace_writeback ? _GEN_6357 : dirty_1_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6643 = replace_writeback ? _GEN_6358 : dirty_2_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6644 = replace_writeback ? _GEN_6359 : dirty_2_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6645 = replace_writeback ? _GEN_6360 : dirty_3_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6646 = replace_writeback ? _GEN_6361 : dirty_3_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6647 = replace_writeback ? _GEN_6362 : dirty_4_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6648 = replace_writeback ? _GEN_6363 : dirty_4_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6649 = replace_writeback ? _GEN_6364 : dirty_5_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6650 = replace_writeback ? _GEN_6365 : dirty_5_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6651 = replace_writeback ? _GEN_6366 : dirty_6_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6652 = replace_writeback ? _GEN_6367 : dirty_6_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6653 = replace_writeback ? _GEN_6368 : dirty_7_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6654 = replace_writeback ? _GEN_6369 : dirty_7_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6655 = replace_writeback ? _GEN_6370 : dirty_8_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6656 = replace_writeback ? _GEN_6371 : dirty_8_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6657 = replace_writeback ? _GEN_6372 : dirty_9_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6658 = replace_writeback ? _GEN_6373 : dirty_9_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6659 = replace_writeback ? _GEN_6374 : dirty_10_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6660 = replace_writeback ? _GEN_6375 : dirty_10_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6661 = replace_writeback ? _GEN_6376 : dirty_11_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6662 = replace_writeback ? _GEN_6377 : dirty_11_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6663 = replace_writeback ? _GEN_6378 : dirty_12_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6664 = replace_writeback ? _GEN_6379 : dirty_12_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6665 = replace_writeback ? _GEN_6380 : dirty_13_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6666 = replace_writeback ? _GEN_6381 : dirty_13_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6667 = replace_writeback ? _GEN_6382 : dirty_14_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6668 = replace_writeback ? _GEN_6383 : dirty_14_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6669 = replace_writeback ? _GEN_6384 : dirty_15_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6670 = replace_writeback ? _GEN_6385 : dirty_15_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6671 = replace_writeback ? _GEN_6386 : dirty_16_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6672 = replace_writeback ? _GEN_6387 : dirty_16_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6673 = replace_writeback ? _GEN_6388 : dirty_17_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6674 = replace_writeback ? _GEN_6389 : dirty_17_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6675 = replace_writeback ? _GEN_6390 : dirty_18_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6676 = replace_writeback ? _GEN_6391 : dirty_18_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6677 = replace_writeback ? _GEN_6392 : dirty_19_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6678 = replace_writeback ? _GEN_6393 : dirty_19_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6679 = replace_writeback ? _GEN_6394 : dirty_20_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6680 = replace_writeback ? _GEN_6395 : dirty_20_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6681 = replace_writeback ? _GEN_6396 : dirty_21_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6682 = replace_writeback ? _GEN_6397 : dirty_21_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6683 = replace_writeback ? _GEN_6398 : dirty_22_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6684 = replace_writeback ? _GEN_6399 : dirty_22_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6685 = replace_writeback ? _GEN_6400 : dirty_23_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6686 = replace_writeback ? _GEN_6401 : dirty_23_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6687 = replace_writeback ? _GEN_6402 : dirty_24_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6688 = replace_writeback ? _GEN_6403 : dirty_24_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6689 = replace_writeback ? _GEN_6404 : dirty_25_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6690 = replace_writeback ? _GEN_6405 : dirty_25_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6691 = replace_writeback ? _GEN_6406 : dirty_26_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6692 = replace_writeback ? _GEN_6407 : dirty_26_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6693 = replace_writeback ? _GEN_6408 : dirty_27_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6694 = replace_writeback ? _GEN_6409 : dirty_27_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6695 = replace_writeback ? _GEN_6410 : dirty_28_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6696 = replace_writeback ? _GEN_6411 : dirty_28_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6697 = replace_writeback ? _GEN_6412 : dirty_29_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6698 = replace_writeback ? _GEN_6413 : dirty_29_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6699 = replace_writeback ? _GEN_6414 : dirty_30_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6700 = replace_writeback ? _GEN_6415 : dirty_30_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6701 = replace_writeback ? _GEN_6416 : dirty_31_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6702 = replace_writeback ? _GEN_6417 : dirty_31_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6703 = replace_writeback ? _GEN_6418 : dirty_32_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6704 = replace_writeback ? _GEN_6419 : dirty_32_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6705 = replace_writeback ? _GEN_6420 : dirty_33_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6706 = replace_writeback ? _GEN_6421 : dirty_33_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6707 = replace_writeback ? _GEN_6422 : dirty_34_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6708 = replace_writeback ? _GEN_6423 : dirty_34_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6709 = replace_writeback ? _GEN_6424 : dirty_35_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6710 = replace_writeback ? _GEN_6425 : dirty_35_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6711 = replace_writeback ? _GEN_6426 : dirty_36_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6712 = replace_writeback ? _GEN_6427 : dirty_36_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6713 = replace_writeback ? _GEN_6428 : dirty_37_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6714 = replace_writeback ? _GEN_6429 : dirty_37_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6715 = replace_writeback ? _GEN_6430 : dirty_38_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6716 = replace_writeback ? _GEN_6431 : dirty_38_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6717 = replace_writeback ? _GEN_6432 : dirty_39_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6718 = replace_writeback ? _GEN_6433 : dirty_39_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6719 = replace_writeback ? _GEN_6434 : dirty_40_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6720 = replace_writeback ? _GEN_6435 : dirty_40_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6721 = replace_writeback ? _GEN_6436 : dirty_41_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6722 = replace_writeback ? _GEN_6437 : dirty_41_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6723 = replace_writeback ? _GEN_6438 : dirty_42_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6724 = replace_writeback ? _GEN_6439 : dirty_42_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6725 = replace_writeback ? _GEN_6440 : dirty_43_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6726 = replace_writeback ? _GEN_6441 : dirty_43_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6727 = replace_writeback ? _GEN_6442 : dirty_44_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6728 = replace_writeback ? _GEN_6443 : dirty_44_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6729 = replace_writeback ? _GEN_6444 : dirty_45_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6730 = replace_writeback ? _GEN_6445 : dirty_45_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6731 = replace_writeback ? _GEN_6446 : dirty_46_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6732 = replace_writeback ? _GEN_6447 : dirty_46_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6733 = replace_writeback ? _GEN_6448 : dirty_47_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6734 = replace_writeback ? _GEN_6449 : dirty_47_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6735 = replace_writeback ? _GEN_6450 : dirty_48_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6736 = replace_writeback ? _GEN_6451 : dirty_48_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6737 = replace_writeback ? _GEN_6452 : dirty_49_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6738 = replace_writeback ? _GEN_6453 : dirty_49_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6739 = replace_writeback ? _GEN_6454 : dirty_50_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6740 = replace_writeback ? _GEN_6455 : dirty_50_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6741 = replace_writeback ? _GEN_6456 : dirty_51_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6742 = replace_writeback ? _GEN_6457 : dirty_51_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6743 = replace_writeback ? _GEN_6458 : dirty_52_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6744 = replace_writeback ? _GEN_6459 : dirty_52_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6745 = replace_writeback ? _GEN_6460 : dirty_53_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6746 = replace_writeback ? _GEN_6461 : dirty_53_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6747 = replace_writeback ? _GEN_6462 : dirty_54_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6748 = replace_writeback ? _GEN_6463 : dirty_54_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6749 = replace_writeback ? _GEN_6464 : dirty_55_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6750 = replace_writeback ? _GEN_6465 : dirty_55_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6751 = replace_writeback ? _GEN_6466 : dirty_56_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6752 = replace_writeback ? _GEN_6467 : dirty_56_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6753 = replace_writeback ? _GEN_6468 : dirty_57_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6754 = replace_writeback ? _GEN_6469 : dirty_57_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6755 = replace_writeback ? _GEN_6470 : dirty_58_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6756 = replace_writeback ? _GEN_6471 : dirty_58_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6757 = replace_writeback ? _GEN_6472 : dirty_59_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6758 = replace_writeback ? _GEN_6473 : dirty_59_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6759 = replace_writeback ? _GEN_6474 : dirty_60_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6760 = replace_writeback ? _GEN_6475 : dirty_60_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6761 = replace_writeback ? _GEN_6476 : dirty_61_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6762 = replace_writeback ? _GEN_6477 : dirty_61_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6763 = replace_writeback ? _GEN_6478 : dirty_62_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6764 = replace_writeback ? _GEN_6479 : dirty_62_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6765 = replace_writeback ? _GEN_6480 : dirty_63_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6766 = replace_writeback ? _GEN_6481 : dirty_63_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6767 = replace_writeback ? _GEN_6482 : dirty_64_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6768 = replace_writeback ? _GEN_6483 : dirty_64_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6769 = replace_writeback ? _GEN_6484 : dirty_65_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6770 = replace_writeback ? _GEN_6485 : dirty_65_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6771 = replace_writeback ? _GEN_6486 : dirty_66_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6772 = replace_writeback ? _GEN_6487 : dirty_66_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6773 = replace_writeback ? _GEN_6488 : dirty_67_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6774 = replace_writeback ? _GEN_6489 : dirty_67_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6775 = replace_writeback ? _GEN_6490 : dirty_68_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6776 = replace_writeback ? _GEN_6491 : dirty_68_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6777 = replace_writeback ? _GEN_6492 : dirty_69_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6778 = replace_writeback ? _GEN_6493 : dirty_69_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6779 = replace_writeback ? _GEN_6494 : dirty_70_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6780 = replace_writeback ? _GEN_6495 : dirty_70_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6781 = replace_writeback ? _GEN_6496 : dirty_71_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6782 = replace_writeback ? _GEN_6497 : dirty_71_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6783 = replace_writeback ? _GEN_6498 : dirty_72_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6784 = replace_writeback ? _GEN_6499 : dirty_72_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6785 = replace_writeback ? _GEN_6500 : dirty_73_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6786 = replace_writeback ? _GEN_6501 : dirty_73_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6787 = replace_writeback ? _GEN_6502 : dirty_74_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6788 = replace_writeback ? _GEN_6503 : dirty_74_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6789 = replace_writeback ? _GEN_6504 : dirty_75_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6790 = replace_writeback ? _GEN_6505 : dirty_75_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6791 = replace_writeback ? _GEN_6506 : dirty_76_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6792 = replace_writeback ? _GEN_6507 : dirty_76_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6793 = replace_writeback ? _GEN_6508 : dirty_77_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6794 = replace_writeback ? _GEN_6509 : dirty_77_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6795 = replace_writeback ? _GEN_6510 : dirty_78_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6796 = replace_writeback ? _GEN_6511 : dirty_78_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6797 = replace_writeback ? _GEN_6512 : dirty_79_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6798 = replace_writeback ? _GEN_6513 : dirty_79_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6799 = replace_writeback ? _GEN_6514 : dirty_80_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6800 = replace_writeback ? _GEN_6515 : dirty_80_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6801 = replace_writeback ? _GEN_6516 : dirty_81_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6802 = replace_writeback ? _GEN_6517 : dirty_81_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6803 = replace_writeback ? _GEN_6518 : dirty_82_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6804 = replace_writeback ? _GEN_6519 : dirty_82_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6805 = replace_writeback ? _GEN_6520 : dirty_83_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6806 = replace_writeback ? _GEN_6521 : dirty_83_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6807 = replace_writeback ? _GEN_6522 : dirty_84_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6808 = replace_writeback ? _GEN_6523 : dirty_84_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6809 = replace_writeback ? _GEN_6524 : dirty_85_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6810 = replace_writeback ? _GEN_6525 : dirty_85_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6811 = replace_writeback ? _GEN_6526 : dirty_86_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6812 = replace_writeback ? _GEN_6527 : dirty_86_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6813 = replace_writeback ? _GEN_6528 : dirty_87_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6814 = replace_writeback ? _GEN_6529 : dirty_87_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6815 = replace_writeback ? _GEN_6530 : dirty_88_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6816 = replace_writeback ? _GEN_6531 : dirty_88_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6817 = replace_writeback ? _GEN_6532 : dirty_89_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6818 = replace_writeback ? _GEN_6533 : dirty_89_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6819 = replace_writeback ? _GEN_6534 : dirty_90_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6820 = replace_writeback ? _GEN_6535 : dirty_90_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6821 = replace_writeback ? _GEN_6536 : dirty_91_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6822 = replace_writeback ? _GEN_6537 : dirty_91_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6823 = replace_writeback ? _GEN_6538 : dirty_92_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6824 = replace_writeback ? _GEN_6539 : dirty_92_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6825 = replace_writeback ? _GEN_6540 : dirty_93_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6826 = replace_writeback ? _GEN_6541 : dirty_93_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6827 = replace_writeback ? _GEN_6542 : dirty_94_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6828 = replace_writeback ? _GEN_6543 : dirty_94_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6829 = replace_writeback ? _GEN_6544 : dirty_95_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6830 = replace_writeback ? _GEN_6545 : dirty_95_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6831 = replace_writeback ? _GEN_6546 : dirty_96_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6832 = replace_writeback ? _GEN_6547 : dirty_96_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6833 = replace_writeback ? _GEN_6548 : dirty_97_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6834 = replace_writeback ? _GEN_6549 : dirty_97_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6835 = replace_writeback ? _GEN_6550 : dirty_98_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6836 = replace_writeback ? _GEN_6551 : dirty_98_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6837 = replace_writeback ? _GEN_6552 : dirty_99_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6838 = replace_writeback ? _GEN_6553 : dirty_99_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6839 = replace_writeback ? _GEN_6554 : dirty_100_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6840 = replace_writeback ? _GEN_6555 : dirty_100_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6841 = replace_writeback ? _GEN_6556 : dirty_101_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6842 = replace_writeback ? _GEN_6557 : dirty_101_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6843 = replace_writeback ? _GEN_6558 : dirty_102_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6844 = replace_writeback ? _GEN_6559 : dirty_102_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6845 = replace_writeback ? _GEN_6560 : dirty_103_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6846 = replace_writeback ? _GEN_6561 : dirty_103_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6847 = replace_writeback ? _GEN_6562 : dirty_104_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6848 = replace_writeback ? _GEN_6563 : dirty_104_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6849 = replace_writeback ? _GEN_6564 : dirty_105_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6850 = replace_writeback ? _GEN_6565 : dirty_105_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6851 = replace_writeback ? _GEN_6566 : dirty_106_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6852 = replace_writeback ? _GEN_6567 : dirty_106_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6853 = replace_writeback ? _GEN_6568 : dirty_107_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6854 = replace_writeback ? _GEN_6569 : dirty_107_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6855 = replace_writeback ? _GEN_6570 : dirty_108_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6856 = replace_writeback ? _GEN_6571 : dirty_108_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6857 = replace_writeback ? _GEN_6572 : dirty_109_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6858 = replace_writeback ? _GEN_6573 : dirty_109_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6859 = replace_writeback ? _GEN_6574 : dirty_110_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6860 = replace_writeback ? _GEN_6575 : dirty_110_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6861 = replace_writeback ? _GEN_6576 : dirty_111_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6862 = replace_writeback ? _GEN_6577 : dirty_111_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6863 = replace_writeback ? _GEN_6578 : dirty_112_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6864 = replace_writeback ? _GEN_6579 : dirty_112_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6865 = replace_writeback ? _GEN_6580 : dirty_113_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6866 = replace_writeback ? _GEN_6581 : dirty_113_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6867 = replace_writeback ? _GEN_6582 : dirty_114_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6868 = replace_writeback ? _GEN_6583 : dirty_114_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6869 = replace_writeback ? _GEN_6584 : dirty_115_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6870 = replace_writeback ? _GEN_6585 : dirty_115_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6871 = replace_writeback ? _GEN_6586 : dirty_116_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6872 = replace_writeback ? _GEN_6587 : dirty_116_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6873 = replace_writeback ? _GEN_6588 : dirty_117_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6874 = replace_writeback ? _GEN_6589 : dirty_117_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6875 = replace_writeback ? _GEN_6590 : dirty_118_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6876 = replace_writeback ? _GEN_6591 : dirty_118_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6877 = replace_writeback ? _GEN_6592 : dirty_119_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6878 = replace_writeback ? _GEN_6593 : dirty_119_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6879 = replace_writeback ? _GEN_6594 : dirty_120_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6880 = replace_writeback ? _GEN_6595 : dirty_120_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6881 = replace_writeback ? _GEN_6596 : dirty_121_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6882 = replace_writeback ? _GEN_6597 : dirty_121_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6883 = replace_writeback ? _GEN_6598 : dirty_122_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6884 = replace_writeback ? _GEN_6599 : dirty_122_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6885 = replace_writeback ? _GEN_6600 : dirty_123_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6886 = replace_writeback ? _GEN_6601 : dirty_123_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6887 = replace_writeback ? _GEN_6602 : dirty_124_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6888 = replace_writeback ? _GEN_6603 : dirty_124_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6889 = replace_writeback ? _GEN_6604 : dirty_125_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6890 = replace_writeback ? _GEN_6605 : dirty_125_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6891 = replace_writeback ? _GEN_6606 : dirty_126_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6892 = replace_writeback ? _GEN_6607 : dirty_126_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6893 = replace_writeback ? _GEN_6608 : dirty_127_0; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6894 = replace_writeback ? _GEN_6609 : dirty_127_1; // @[DCache.scala 420:35 69:22]
  wire  _GEN_6895 = replace_writeback ? _GEN_6610 : replace_writeback; // @[DCache.scala 420:35 101:40]
  wire [31:0] _ar_addr_T_5 = {M_mem_pa[31:6],6'h0}; // @[Cat.scala 33:92]
  wire [3:0] _GEN_6896 = ~_GEN_441 ? 4'hf : bram_replace_wea_0; // @[DCache.scala 468:{49,49} 73:33]
  wire [3:0] _GEN_6897 = _GEN_441 ? 4'hf : bram_replace_wea_1; // @[DCache.scala 468:{49,49} 73:33]
  wire  _GEN_6898 = _GEN_11689 | tag_wstrb_0; // @[DCache.scala 469:{49,49} 72:33]
  wire  _GEN_6899 = _GEN_441 | tag_wstrb_1; // @[DCache.scala 469:{49,49} 72:33]
  wire [31:0] _GEN_6900 = ~ar_handshake ? _ar_addr_T_5 : ar_addr; // @[DCache.scala 199:24 461:31 462:49]
  wire [7:0] _GEN_6901 = ~ar_handshake ? 8'hf : ar_len; // @[DCache.scala 199:24 461:31 463:49]
  wire [2:0] _GEN_6902 = ~ar_handshake ? 3'h2 : ar_size; // @[DCache.scala 199:24 461:31 464:49]
  wire  _GEN_6903 = ~ar_handshake | arvalid; // @[DCache.scala 200:24 461:31 465:49]
  wire  _GEN_6904 = ~ar_handshake | rready; // @[DCache.scala 203:23 461:31 466:49]
  wire  _GEN_6905 = ~ar_handshake | ar_handshake; // @[DCache.scala 461:31 467:49 99:40]
  wire [3:0] _GEN_6906 = ~ar_handshake ? _GEN_6896 : bram_replace_wea_0; // @[DCache.scala 461:31 73:33]
  wire [3:0] _GEN_6907 = ~ar_handshake ? _GEN_6897 : bram_replace_wea_1; // @[DCache.scala 461:31 73:33]
  wire  _GEN_6908 = ~ar_handshake ? _GEN_6898 : tag_wstrb_0; // @[DCache.scala 461:31 72:33]
  wire  _GEN_6909 = ~ar_handshake ? _GEN_6899 : tag_wstrb_1; // @[DCache.scala 461:31 72:33]
  wire [19:0] _GEN_6910 = ~ar_handshake ? M_mem_pa[31:12] : tag_wdata; // @[DCache.scala 461:31 470:49 77:26]
  wire  _T_57 = io_axi_ar_ready & io_axi_ar_valid; // @[Decoupled.scala 52:35]
  wire  _GEN_6911 = ~_GEN_441 ? 1'h0 : _GEN_6908; // @[DCache.scala 473:{42,42}]
  wire  _GEN_6912 = _GEN_441 ? 1'h0 : _GEN_6909; // @[DCache.scala 473:{42,42}]
  wire  _GEN_6913 = _T_57 ? _GEN_6911 : _GEN_6908; // @[DCache.scala 472:32]
  wire  _GEN_6914 = _T_57 ? _GEN_6912 : _GEN_6909; // @[DCache.scala 472:32]
  wire  _GEN_6915 = _T_57 ? 1'h0 : _GEN_6903; // @[DCache.scala 472:32 474:42]
  wire  _T_58 = io_axi_r_ready & io_axi_r_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _GEN_6916 = ~_GEN_441 ? 4'h0 : _GEN_6906; // @[DCache.scala 479:{51,51}]
  wire [3:0] _GEN_6917 = _GEN_441 ? 4'h0 : _GEN_6907; // @[DCache.scala 479:{51,51}]
  wire [9:0] _bram_replace_write_addr_T_2 = bram_replace_write_addr + 10'h1; // @[DCache.scala 481:66]
  wire  _GEN_6918 = io_axi_r_bits_last ? 1'h0 : _GEN_6904; // @[DCache.scala 477:38 478:51]
  wire [3:0] _GEN_6919 = io_axi_r_bits_last ? _GEN_6916 : _GEN_6906; // @[DCache.scala 477:38]
  wire [3:0] _GEN_6920 = io_axi_r_bits_last ? _GEN_6917 : _GEN_6907; // @[DCache.scala 477:38]
  wire [9:0] _GEN_6921 = io_axi_r_bits_last ? bram_replace_write_addr : _bram_replace_write_addr_T_2; // @[DCache.scala 477:38 481:39 92:40]
  wire  _GEN_6922 = _T_58 ? _GEN_6918 : _GEN_6904; // @[DCache.scala 476:31]
  wire [3:0] _GEN_6923 = _T_58 ? _GEN_6919 : _GEN_6906; // @[DCache.scala 476:31]
  wire [3:0] _GEN_6924 = _T_58 ? _GEN_6920 : _GEN_6907; // @[DCache.scala 476:31]
  wire [9:0] _GEN_6925 = _T_58 ? _GEN_6921 : bram_replace_write_addr; // @[DCache.scala 476:31 92:40]
  wire  _T_66 = (~replace_writeback | io_axi_b_valid) & (ar_handshake & io_axi_r_valid & io_axi_r_bits_last |
    ar_handshake & ~rready); // @[DCache.scala 485:54]
  wire  _GEN_6926 = _GEN_11687 & _GEN_11689 | valid_0_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6927 = _GEN_11687 & _GEN_441 | valid_0_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6928 = _GEN_11688 & _GEN_11689 | valid_1_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6929 = _GEN_11688 & _GEN_441 | valid_1_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6930 = _GEN_11691 & _GEN_11689 | valid_2_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6931 = _GEN_11691 & _GEN_441 | valid_2_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6932 = _GEN_11694 & _GEN_11689 | valid_3_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6933 = _GEN_11694 & _GEN_441 | valid_3_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6934 = _GEN_11697 & _GEN_11689 | valid_4_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6935 = _GEN_11697 & _GEN_441 | valid_4_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6936 = _GEN_11700 & _GEN_11689 | valid_5_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6937 = _GEN_11700 & _GEN_441 | valid_5_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6938 = _GEN_11703 & _GEN_11689 | valid_6_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6939 = _GEN_11703 & _GEN_441 | valid_6_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6940 = _GEN_11706 & _GEN_11689 | valid_7_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6941 = _GEN_11706 & _GEN_441 | valid_7_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6942 = _GEN_11709 & _GEN_11689 | valid_8_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6943 = _GEN_11709 & _GEN_441 | valid_8_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6944 = _GEN_11712 & _GEN_11689 | valid_9_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6945 = _GEN_11712 & _GEN_441 | valid_9_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6946 = _GEN_11715 & _GEN_11689 | valid_10_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6947 = _GEN_11715 & _GEN_441 | valid_10_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6948 = _GEN_11718 & _GEN_11689 | valid_11_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6949 = _GEN_11718 & _GEN_441 | valid_11_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6950 = _GEN_11721 & _GEN_11689 | valid_12_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6951 = _GEN_11721 & _GEN_441 | valid_12_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6952 = _GEN_11724 & _GEN_11689 | valid_13_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6953 = _GEN_11724 & _GEN_441 | valid_13_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6954 = _GEN_11727 & _GEN_11689 | valid_14_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6955 = _GEN_11727 & _GEN_441 | valid_14_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6956 = _GEN_11730 & _GEN_11689 | valid_15_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6957 = _GEN_11730 & _GEN_441 | valid_15_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6958 = _GEN_11733 & _GEN_11689 | valid_16_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6959 = _GEN_11733 & _GEN_441 | valid_16_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6960 = _GEN_11736 & _GEN_11689 | valid_17_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6961 = _GEN_11736 & _GEN_441 | valid_17_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6962 = _GEN_11739 & _GEN_11689 | valid_18_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6963 = _GEN_11739 & _GEN_441 | valid_18_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6964 = _GEN_11742 & _GEN_11689 | valid_19_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6965 = _GEN_11742 & _GEN_441 | valid_19_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6966 = _GEN_11745 & _GEN_11689 | valid_20_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6967 = _GEN_11745 & _GEN_441 | valid_20_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6968 = _GEN_11748 & _GEN_11689 | valid_21_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6969 = _GEN_11748 & _GEN_441 | valid_21_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6970 = _GEN_11751 & _GEN_11689 | valid_22_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6971 = _GEN_11751 & _GEN_441 | valid_22_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6972 = _GEN_11754 & _GEN_11689 | valid_23_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6973 = _GEN_11754 & _GEN_441 | valid_23_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6974 = _GEN_11757 & _GEN_11689 | valid_24_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6975 = _GEN_11757 & _GEN_441 | valid_24_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6976 = _GEN_11760 & _GEN_11689 | valid_25_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6977 = _GEN_11760 & _GEN_441 | valid_25_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6978 = _GEN_11763 & _GEN_11689 | valid_26_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6979 = _GEN_11763 & _GEN_441 | valid_26_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6980 = _GEN_11766 & _GEN_11689 | valid_27_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6981 = _GEN_11766 & _GEN_441 | valid_27_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6982 = _GEN_11769 & _GEN_11689 | valid_28_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6983 = _GEN_11769 & _GEN_441 | valid_28_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6984 = _GEN_11772 & _GEN_11689 | valid_29_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6985 = _GEN_11772 & _GEN_441 | valid_29_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6986 = _GEN_11775 & _GEN_11689 | valid_30_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6987 = _GEN_11775 & _GEN_441 | valid_30_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6988 = _GEN_11778 & _GEN_11689 | valid_31_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6989 = _GEN_11778 & _GEN_441 | valid_31_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6990 = _GEN_11781 & _GEN_11689 | valid_32_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6991 = _GEN_11781 & _GEN_441 | valid_32_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6992 = _GEN_11784 & _GEN_11689 | valid_33_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6993 = _GEN_11784 & _GEN_441 | valid_33_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6994 = _GEN_11787 & _GEN_11689 | valid_34_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6995 = _GEN_11787 & _GEN_441 | valid_34_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6996 = _GEN_11790 & _GEN_11689 | valid_35_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6997 = _GEN_11790 & _GEN_441 | valid_35_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6998 = _GEN_11793 & _GEN_11689 | valid_36_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_6999 = _GEN_11793 & _GEN_441 | valid_36_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7000 = _GEN_11796 & _GEN_11689 | valid_37_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7001 = _GEN_11796 & _GEN_441 | valid_37_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7002 = _GEN_11799 & _GEN_11689 | valid_38_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7003 = _GEN_11799 & _GEN_441 | valid_38_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7004 = _GEN_11802 & _GEN_11689 | valid_39_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7005 = _GEN_11802 & _GEN_441 | valid_39_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7006 = _GEN_11805 & _GEN_11689 | valid_40_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7007 = _GEN_11805 & _GEN_441 | valid_40_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7008 = _GEN_11808 & _GEN_11689 | valid_41_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7009 = _GEN_11808 & _GEN_441 | valid_41_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7010 = _GEN_11811 & _GEN_11689 | valid_42_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7011 = _GEN_11811 & _GEN_441 | valid_42_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7012 = _GEN_11814 & _GEN_11689 | valid_43_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7013 = _GEN_11814 & _GEN_441 | valid_43_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7014 = _GEN_11817 & _GEN_11689 | valid_44_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7015 = _GEN_11817 & _GEN_441 | valid_44_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7016 = _GEN_11820 & _GEN_11689 | valid_45_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7017 = _GEN_11820 & _GEN_441 | valid_45_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7018 = _GEN_11823 & _GEN_11689 | valid_46_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7019 = _GEN_11823 & _GEN_441 | valid_46_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7020 = _GEN_11826 & _GEN_11689 | valid_47_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7021 = _GEN_11826 & _GEN_441 | valid_47_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7022 = _GEN_11829 & _GEN_11689 | valid_48_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7023 = _GEN_11829 & _GEN_441 | valid_48_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7024 = _GEN_11832 & _GEN_11689 | valid_49_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7025 = _GEN_11832 & _GEN_441 | valid_49_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7026 = _GEN_11835 & _GEN_11689 | valid_50_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7027 = _GEN_11835 & _GEN_441 | valid_50_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7028 = _GEN_11838 & _GEN_11689 | valid_51_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7029 = _GEN_11838 & _GEN_441 | valid_51_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7030 = _GEN_11841 & _GEN_11689 | valid_52_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7031 = _GEN_11841 & _GEN_441 | valid_52_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7032 = _GEN_11844 & _GEN_11689 | valid_53_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7033 = _GEN_11844 & _GEN_441 | valid_53_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7034 = _GEN_11847 & _GEN_11689 | valid_54_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7035 = _GEN_11847 & _GEN_441 | valid_54_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7036 = _GEN_11850 & _GEN_11689 | valid_55_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7037 = _GEN_11850 & _GEN_441 | valid_55_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7038 = _GEN_11853 & _GEN_11689 | valid_56_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7039 = _GEN_11853 & _GEN_441 | valid_56_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7040 = _GEN_11856 & _GEN_11689 | valid_57_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7041 = _GEN_11856 & _GEN_441 | valid_57_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7042 = _GEN_11859 & _GEN_11689 | valid_58_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7043 = _GEN_11859 & _GEN_441 | valid_58_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7044 = _GEN_11862 & _GEN_11689 | valid_59_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7045 = _GEN_11862 & _GEN_441 | valid_59_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7046 = _GEN_11865 & _GEN_11689 | valid_60_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7047 = _GEN_11865 & _GEN_441 | valid_60_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7048 = _GEN_11868 & _GEN_11689 | valid_61_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7049 = _GEN_11868 & _GEN_441 | valid_61_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7050 = _GEN_11871 & _GEN_11689 | valid_62_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7051 = _GEN_11871 & _GEN_441 | valid_62_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7052 = _GEN_11874 & _GEN_11689 | valid_63_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7053 = _GEN_11874 & _GEN_441 | valid_63_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7054 = _GEN_11878 & _GEN_11689 | valid_64_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7055 = _GEN_11878 & _GEN_441 | valid_64_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7056 = _GEN_11883 & _GEN_11689 | valid_65_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7057 = _GEN_11883 & _GEN_441 | valid_65_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7058 = _GEN_11888 & _GEN_11689 | valid_66_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7059 = _GEN_11888 & _GEN_441 | valid_66_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7060 = _GEN_11893 & _GEN_11689 | valid_67_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7061 = _GEN_11893 & _GEN_441 | valid_67_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7062 = _GEN_11898 & _GEN_11689 | valid_68_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7063 = _GEN_11898 & _GEN_441 | valid_68_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7064 = _GEN_11903 & _GEN_11689 | valid_69_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7065 = _GEN_11903 & _GEN_441 | valid_69_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7066 = _GEN_11908 & _GEN_11689 | valid_70_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7067 = _GEN_11908 & _GEN_441 | valid_70_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7068 = _GEN_11913 & _GEN_11689 | valid_71_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7069 = _GEN_11913 & _GEN_441 | valid_71_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7070 = _GEN_11918 & _GEN_11689 | valid_72_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7071 = _GEN_11918 & _GEN_441 | valid_72_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7072 = _GEN_11923 & _GEN_11689 | valid_73_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7073 = _GEN_11923 & _GEN_441 | valid_73_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7074 = _GEN_11928 & _GEN_11689 | valid_74_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7075 = _GEN_11928 & _GEN_441 | valid_74_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7076 = _GEN_11933 & _GEN_11689 | valid_75_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7077 = _GEN_11933 & _GEN_441 | valid_75_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7078 = _GEN_11938 & _GEN_11689 | valid_76_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7079 = _GEN_11938 & _GEN_441 | valid_76_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7080 = _GEN_11943 & _GEN_11689 | valid_77_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7081 = _GEN_11943 & _GEN_441 | valid_77_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7082 = _GEN_11948 & _GEN_11689 | valid_78_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7083 = _GEN_11948 & _GEN_441 | valid_78_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7084 = _GEN_11953 & _GEN_11689 | valid_79_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7085 = _GEN_11953 & _GEN_441 | valid_79_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7086 = _GEN_11958 & _GEN_11689 | valid_80_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7087 = _GEN_11958 & _GEN_441 | valid_80_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7088 = _GEN_11963 & _GEN_11689 | valid_81_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7089 = _GEN_11963 & _GEN_441 | valid_81_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7090 = _GEN_11968 & _GEN_11689 | valid_82_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7091 = _GEN_11968 & _GEN_441 | valid_82_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7092 = _GEN_11973 & _GEN_11689 | valid_83_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7093 = _GEN_11973 & _GEN_441 | valid_83_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7094 = _GEN_11978 & _GEN_11689 | valid_84_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7095 = _GEN_11978 & _GEN_441 | valid_84_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7096 = _GEN_11983 & _GEN_11689 | valid_85_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7097 = _GEN_11983 & _GEN_441 | valid_85_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7098 = _GEN_11988 & _GEN_11689 | valid_86_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7099 = _GEN_11988 & _GEN_441 | valid_86_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7100 = _GEN_11993 & _GEN_11689 | valid_87_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7101 = _GEN_11993 & _GEN_441 | valid_87_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7102 = _GEN_11998 & _GEN_11689 | valid_88_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7103 = _GEN_11998 & _GEN_441 | valid_88_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7104 = _GEN_12003 & _GEN_11689 | valid_89_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7105 = _GEN_12003 & _GEN_441 | valid_89_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7106 = _GEN_12008 & _GEN_11689 | valid_90_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7107 = _GEN_12008 & _GEN_441 | valid_90_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7108 = _GEN_12013 & _GEN_11689 | valid_91_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7109 = _GEN_12013 & _GEN_441 | valid_91_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7110 = _GEN_12018 & _GEN_11689 | valid_92_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7111 = _GEN_12018 & _GEN_441 | valid_92_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7112 = _GEN_12023 & _GEN_11689 | valid_93_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7113 = _GEN_12023 & _GEN_441 | valid_93_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7114 = _GEN_12028 & _GEN_11689 | valid_94_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7115 = _GEN_12028 & _GEN_441 | valid_94_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7116 = _GEN_12033 & _GEN_11689 | valid_95_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7117 = _GEN_12033 & _GEN_441 | valid_95_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7118 = _GEN_12038 & _GEN_11689 | valid_96_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7119 = _GEN_12038 & _GEN_441 | valid_96_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7120 = _GEN_12043 & _GEN_11689 | valid_97_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7121 = _GEN_12043 & _GEN_441 | valid_97_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7122 = _GEN_12048 & _GEN_11689 | valid_98_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7123 = _GEN_12048 & _GEN_441 | valid_98_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7124 = _GEN_12053 & _GEN_11689 | valid_99_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7125 = _GEN_12053 & _GEN_441 | valid_99_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7126 = _GEN_12058 & _GEN_11689 | valid_100_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7127 = _GEN_12058 & _GEN_441 | valid_100_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7128 = _GEN_12063 & _GEN_11689 | valid_101_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7129 = _GEN_12063 & _GEN_441 | valid_101_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7130 = _GEN_12068 & _GEN_11689 | valid_102_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7131 = _GEN_12068 & _GEN_441 | valid_102_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7132 = _GEN_12073 & _GEN_11689 | valid_103_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7133 = _GEN_12073 & _GEN_441 | valid_103_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7134 = _GEN_12078 & _GEN_11689 | valid_104_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7135 = _GEN_12078 & _GEN_441 | valid_104_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7136 = _GEN_12083 & _GEN_11689 | valid_105_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7137 = _GEN_12083 & _GEN_441 | valid_105_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7138 = _GEN_12088 & _GEN_11689 | valid_106_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7139 = _GEN_12088 & _GEN_441 | valid_106_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7140 = _GEN_12093 & _GEN_11689 | valid_107_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7141 = _GEN_12093 & _GEN_441 | valid_107_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7142 = _GEN_12098 & _GEN_11689 | valid_108_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7143 = _GEN_12098 & _GEN_441 | valid_108_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7144 = _GEN_12103 & _GEN_11689 | valid_109_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7145 = _GEN_12103 & _GEN_441 | valid_109_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7146 = _GEN_12108 & _GEN_11689 | valid_110_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7147 = _GEN_12108 & _GEN_441 | valid_110_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7148 = _GEN_12113 & _GEN_11689 | valid_111_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7149 = _GEN_12113 & _GEN_441 | valid_111_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7150 = _GEN_12118 & _GEN_11689 | valid_112_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7151 = _GEN_12118 & _GEN_441 | valid_112_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7152 = _GEN_12123 & _GEN_11689 | valid_113_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7153 = _GEN_12123 & _GEN_441 | valid_113_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7154 = _GEN_12128 & _GEN_11689 | valid_114_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7155 = _GEN_12128 & _GEN_441 | valid_114_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7156 = _GEN_12133 & _GEN_11689 | valid_115_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7157 = _GEN_12133 & _GEN_441 | valid_115_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7158 = _GEN_12138 & _GEN_11689 | valid_116_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7159 = _GEN_12138 & _GEN_441 | valid_116_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7160 = _GEN_12143 & _GEN_11689 | valid_117_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7161 = _GEN_12143 & _GEN_441 | valid_117_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7162 = _GEN_12148 & _GEN_11689 | valid_118_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7163 = _GEN_12148 & _GEN_441 | valid_118_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7164 = _GEN_12153 & _GEN_11689 | valid_119_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7165 = _GEN_12153 & _GEN_441 | valid_119_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7166 = _GEN_12158 & _GEN_11689 | valid_120_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7167 = _GEN_12158 & _GEN_441 | valid_120_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7168 = _GEN_12163 & _GEN_11689 | valid_121_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7169 = _GEN_12163 & _GEN_441 | valid_121_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7170 = _GEN_12168 & _GEN_11689 | valid_122_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7171 = _GEN_12168 & _GEN_441 | valid_122_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7172 = _GEN_12173 & _GEN_11689 | valid_123_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7173 = _GEN_12173 & _GEN_441 | valid_123_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7174 = _GEN_12178 & _GEN_11689 | valid_124_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7175 = _GEN_12178 & _GEN_441 | valid_124_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7176 = _GEN_12183 & _GEN_11689 | valid_125_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7177 = _GEN_12183 & _GEN_441 | valid_125_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7178 = _GEN_12188 & _GEN_11689 | valid_126_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7179 = _GEN_12188 & _GEN_441 | valid_126_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7180 = _GEN_12193 & _GEN_11689 | valid_127_0; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7181 = _GEN_12193 & _GEN_441 | valid_127_1; // @[DCache.scala 488:{52,52} 68:22]
  wire  _GEN_7182 = _T_66 ? 1'h0 : bram_use_replace_addr; // @[DCache.scala 486:13 487:52 95:40]
  wire  _GEN_7183 = _T_66 ? _GEN_6926 : valid_0_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7184 = _T_66 ? _GEN_6927 : valid_0_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7185 = _T_66 ? _GEN_6928 : valid_1_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7186 = _T_66 ? _GEN_6929 : valid_1_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7187 = _T_66 ? _GEN_6930 : valid_2_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7188 = _T_66 ? _GEN_6931 : valid_2_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7189 = _T_66 ? _GEN_6932 : valid_3_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7190 = _T_66 ? _GEN_6933 : valid_3_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7191 = _T_66 ? _GEN_6934 : valid_4_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7192 = _T_66 ? _GEN_6935 : valid_4_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7193 = _T_66 ? _GEN_6936 : valid_5_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7194 = _T_66 ? _GEN_6937 : valid_5_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7195 = _T_66 ? _GEN_6938 : valid_6_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7196 = _T_66 ? _GEN_6939 : valid_6_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7197 = _T_66 ? _GEN_6940 : valid_7_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7198 = _T_66 ? _GEN_6941 : valid_7_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7199 = _T_66 ? _GEN_6942 : valid_8_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7200 = _T_66 ? _GEN_6943 : valid_8_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7201 = _T_66 ? _GEN_6944 : valid_9_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7202 = _T_66 ? _GEN_6945 : valid_9_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7203 = _T_66 ? _GEN_6946 : valid_10_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7204 = _T_66 ? _GEN_6947 : valid_10_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7205 = _T_66 ? _GEN_6948 : valid_11_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7206 = _T_66 ? _GEN_6949 : valid_11_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7207 = _T_66 ? _GEN_6950 : valid_12_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7208 = _T_66 ? _GEN_6951 : valid_12_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7209 = _T_66 ? _GEN_6952 : valid_13_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7210 = _T_66 ? _GEN_6953 : valid_13_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7211 = _T_66 ? _GEN_6954 : valid_14_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7212 = _T_66 ? _GEN_6955 : valid_14_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7213 = _T_66 ? _GEN_6956 : valid_15_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7214 = _T_66 ? _GEN_6957 : valid_15_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7215 = _T_66 ? _GEN_6958 : valid_16_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7216 = _T_66 ? _GEN_6959 : valid_16_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7217 = _T_66 ? _GEN_6960 : valid_17_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7218 = _T_66 ? _GEN_6961 : valid_17_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7219 = _T_66 ? _GEN_6962 : valid_18_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7220 = _T_66 ? _GEN_6963 : valid_18_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7221 = _T_66 ? _GEN_6964 : valid_19_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7222 = _T_66 ? _GEN_6965 : valid_19_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7223 = _T_66 ? _GEN_6966 : valid_20_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7224 = _T_66 ? _GEN_6967 : valid_20_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7225 = _T_66 ? _GEN_6968 : valid_21_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7226 = _T_66 ? _GEN_6969 : valid_21_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7227 = _T_66 ? _GEN_6970 : valid_22_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7228 = _T_66 ? _GEN_6971 : valid_22_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7229 = _T_66 ? _GEN_6972 : valid_23_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7230 = _T_66 ? _GEN_6973 : valid_23_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7231 = _T_66 ? _GEN_6974 : valid_24_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7232 = _T_66 ? _GEN_6975 : valid_24_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7233 = _T_66 ? _GEN_6976 : valid_25_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7234 = _T_66 ? _GEN_6977 : valid_25_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7235 = _T_66 ? _GEN_6978 : valid_26_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7236 = _T_66 ? _GEN_6979 : valid_26_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7237 = _T_66 ? _GEN_6980 : valid_27_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7238 = _T_66 ? _GEN_6981 : valid_27_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7239 = _T_66 ? _GEN_6982 : valid_28_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7240 = _T_66 ? _GEN_6983 : valid_28_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7241 = _T_66 ? _GEN_6984 : valid_29_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7242 = _T_66 ? _GEN_6985 : valid_29_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7243 = _T_66 ? _GEN_6986 : valid_30_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7244 = _T_66 ? _GEN_6987 : valid_30_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7245 = _T_66 ? _GEN_6988 : valid_31_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7246 = _T_66 ? _GEN_6989 : valid_31_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7247 = _T_66 ? _GEN_6990 : valid_32_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7248 = _T_66 ? _GEN_6991 : valid_32_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7249 = _T_66 ? _GEN_6992 : valid_33_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7250 = _T_66 ? _GEN_6993 : valid_33_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7251 = _T_66 ? _GEN_6994 : valid_34_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7252 = _T_66 ? _GEN_6995 : valid_34_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7253 = _T_66 ? _GEN_6996 : valid_35_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7254 = _T_66 ? _GEN_6997 : valid_35_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7255 = _T_66 ? _GEN_6998 : valid_36_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7256 = _T_66 ? _GEN_6999 : valid_36_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7257 = _T_66 ? _GEN_7000 : valid_37_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7258 = _T_66 ? _GEN_7001 : valid_37_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7259 = _T_66 ? _GEN_7002 : valid_38_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7260 = _T_66 ? _GEN_7003 : valid_38_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7261 = _T_66 ? _GEN_7004 : valid_39_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7262 = _T_66 ? _GEN_7005 : valid_39_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7263 = _T_66 ? _GEN_7006 : valid_40_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7264 = _T_66 ? _GEN_7007 : valid_40_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7265 = _T_66 ? _GEN_7008 : valid_41_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7266 = _T_66 ? _GEN_7009 : valid_41_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7267 = _T_66 ? _GEN_7010 : valid_42_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7268 = _T_66 ? _GEN_7011 : valid_42_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7269 = _T_66 ? _GEN_7012 : valid_43_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7270 = _T_66 ? _GEN_7013 : valid_43_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7271 = _T_66 ? _GEN_7014 : valid_44_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7272 = _T_66 ? _GEN_7015 : valid_44_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7273 = _T_66 ? _GEN_7016 : valid_45_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7274 = _T_66 ? _GEN_7017 : valid_45_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7275 = _T_66 ? _GEN_7018 : valid_46_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7276 = _T_66 ? _GEN_7019 : valid_46_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7277 = _T_66 ? _GEN_7020 : valid_47_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7278 = _T_66 ? _GEN_7021 : valid_47_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7279 = _T_66 ? _GEN_7022 : valid_48_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7280 = _T_66 ? _GEN_7023 : valid_48_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7281 = _T_66 ? _GEN_7024 : valid_49_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7282 = _T_66 ? _GEN_7025 : valid_49_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7283 = _T_66 ? _GEN_7026 : valid_50_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7284 = _T_66 ? _GEN_7027 : valid_50_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7285 = _T_66 ? _GEN_7028 : valid_51_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7286 = _T_66 ? _GEN_7029 : valid_51_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7287 = _T_66 ? _GEN_7030 : valid_52_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7288 = _T_66 ? _GEN_7031 : valid_52_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7289 = _T_66 ? _GEN_7032 : valid_53_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7290 = _T_66 ? _GEN_7033 : valid_53_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7291 = _T_66 ? _GEN_7034 : valid_54_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7292 = _T_66 ? _GEN_7035 : valid_54_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7293 = _T_66 ? _GEN_7036 : valid_55_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7294 = _T_66 ? _GEN_7037 : valid_55_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7295 = _T_66 ? _GEN_7038 : valid_56_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7296 = _T_66 ? _GEN_7039 : valid_56_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7297 = _T_66 ? _GEN_7040 : valid_57_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7298 = _T_66 ? _GEN_7041 : valid_57_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7299 = _T_66 ? _GEN_7042 : valid_58_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7300 = _T_66 ? _GEN_7043 : valid_58_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7301 = _T_66 ? _GEN_7044 : valid_59_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7302 = _T_66 ? _GEN_7045 : valid_59_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7303 = _T_66 ? _GEN_7046 : valid_60_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7304 = _T_66 ? _GEN_7047 : valid_60_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7305 = _T_66 ? _GEN_7048 : valid_61_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7306 = _T_66 ? _GEN_7049 : valid_61_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7307 = _T_66 ? _GEN_7050 : valid_62_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7308 = _T_66 ? _GEN_7051 : valid_62_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7309 = _T_66 ? _GEN_7052 : valid_63_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7310 = _T_66 ? _GEN_7053 : valid_63_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7311 = _T_66 ? _GEN_7054 : valid_64_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7312 = _T_66 ? _GEN_7055 : valid_64_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7313 = _T_66 ? _GEN_7056 : valid_65_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7314 = _T_66 ? _GEN_7057 : valid_65_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7315 = _T_66 ? _GEN_7058 : valid_66_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7316 = _T_66 ? _GEN_7059 : valid_66_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7317 = _T_66 ? _GEN_7060 : valid_67_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7318 = _T_66 ? _GEN_7061 : valid_67_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7319 = _T_66 ? _GEN_7062 : valid_68_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7320 = _T_66 ? _GEN_7063 : valid_68_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7321 = _T_66 ? _GEN_7064 : valid_69_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7322 = _T_66 ? _GEN_7065 : valid_69_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7323 = _T_66 ? _GEN_7066 : valid_70_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7324 = _T_66 ? _GEN_7067 : valid_70_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7325 = _T_66 ? _GEN_7068 : valid_71_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7326 = _T_66 ? _GEN_7069 : valid_71_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7327 = _T_66 ? _GEN_7070 : valid_72_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7328 = _T_66 ? _GEN_7071 : valid_72_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7329 = _T_66 ? _GEN_7072 : valid_73_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7330 = _T_66 ? _GEN_7073 : valid_73_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7331 = _T_66 ? _GEN_7074 : valid_74_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7332 = _T_66 ? _GEN_7075 : valid_74_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7333 = _T_66 ? _GEN_7076 : valid_75_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7334 = _T_66 ? _GEN_7077 : valid_75_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7335 = _T_66 ? _GEN_7078 : valid_76_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7336 = _T_66 ? _GEN_7079 : valid_76_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7337 = _T_66 ? _GEN_7080 : valid_77_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7338 = _T_66 ? _GEN_7081 : valid_77_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7339 = _T_66 ? _GEN_7082 : valid_78_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7340 = _T_66 ? _GEN_7083 : valid_78_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7341 = _T_66 ? _GEN_7084 : valid_79_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7342 = _T_66 ? _GEN_7085 : valid_79_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7343 = _T_66 ? _GEN_7086 : valid_80_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7344 = _T_66 ? _GEN_7087 : valid_80_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7345 = _T_66 ? _GEN_7088 : valid_81_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7346 = _T_66 ? _GEN_7089 : valid_81_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7347 = _T_66 ? _GEN_7090 : valid_82_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7348 = _T_66 ? _GEN_7091 : valid_82_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7349 = _T_66 ? _GEN_7092 : valid_83_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7350 = _T_66 ? _GEN_7093 : valid_83_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7351 = _T_66 ? _GEN_7094 : valid_84_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7352 = _T_66 ? _GEN_7095 : valid_84_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7353 = _T_66 ? _GEN_7096 : valid_85_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7354 = _T_66 ? _GEN_7097 : valid_85_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7355 = _T_66 ? _GEN_7098 : valid_86_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7356 = _T_66 ? _GEN_7099 : valid_86_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7357 = _T_66 ? _GEN_7100 : valid_87_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7358 = _T_66 ? _GEN_7101 : valid_87_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7359 = _T_66 ? _GEN_7102 : valid_88_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7360 = _T_66 ? _GEN_7103 : valid_88_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7361 = _T_66 ? _GEN_7104 : valid_89_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7362 = _T_66 ? _GEN_7105 : valid_89_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7363 = _T_66 ? _GEN_7106 : valid_90_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7364 = _T_66 ? _GEN_7107 : valid_90_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7365 = _T_66 ? _GEN_7108 : valid_91_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7366 = _T_66 ? _GEN_7109 : valid_91_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7367 = _T_66 ? _GEN_7110 : valid_92_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7368 = _T_66 ? _GEN_7111 : valid_92_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7369 = _T_66 ? _GEN_7112 : valid_93_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7370 = _T_66 ? _GEN_7113 : valid_93_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7371 = _T_66 ? _GEN_7114 : valid_94_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7372 = _T_66 ? _GEN_7115 : valid_94_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7373 = _T_66 ? _GEN_7116 : valid_95_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7374 = _T_66 ? _GEN_7117 : valid_95_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7375 = _T_66 ? _GEN_7118 : valid_96_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7376 = _T_66 ? _GEN_7119 : valid_96_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7377 = _T_66 ? _GEN_7120 : valid_97_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7378 = _T_66 ? _GEN_7121 : valid_97_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7379 = _T_66 ? _GEN_7122 : valid_98_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7380 = _T_66 ? _GEN_7123 : valid_98_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7381 = _T_66 ? _GEN_7124 : valid_99_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7382 = _T_66 ? _GEN_7125 : valid_99_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7383 = _T_66 ? _GEN_7126 : valid_100_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7384 = _T_66 ? _GEN_7127 : valid_100_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7385 = _T_66 ? _GEN_7128 : valid_101_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7386 = _T_66 ? _GEN_7129 : valid_101_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7387 = _T_66 ? _GEN_7130 : valid_102_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7388 = _T_66 ? _GEN_7131 : valid_102_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7389 = _T_66 ? _GEN_7132 : valid_103_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7390 = _T_66 ? _GEN_7133 : valid_103_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7391 = _T_66 ? _GEN_7134 : valid_104_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7392 = _T_66 ? _GEN_7135 : valid_104_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7393 = _T_66 ? _GEN_7136 : valid_105_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7394 = _T_66 ? _GEN_7137 : valid_105_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7395 = _T_66 ? _GEN_7138 : valid_106_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7396 = _T_66 ? _GEN_7139 : valid_106_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7397 = _T_66 ? _GEN_7140 : valid_107_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7398 = _T_66 ? _GEN_7141 : valid_107_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7399 = _T_66 ? _GEN_7142 : valid_108_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7400 = _T_66 ? _GEN_7143 : valid_108_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7401 = _T_66 ? _GEN_7144 : valid_109_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7402 = _T_66 ? _GEN_7145 : valid_109_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7403 = _T_66 ? _GEN_7146 : valid_110_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7404 = _T_66 ? _GEN_7147 : valid_110_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7405 = _T_66 ? _GEN_7148 : valid_111_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7406 = _T_66 ? _GEN_7149 : valid_111_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7407 = _T_66 ? _GEN_7150 : valid_112_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7408 = _T_66 ? _GEN_7151 : valid_112_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7409 = _T_66 ? _GEN_7152 : valid_113_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7410 = _T_66 ? _GEN_7153 : valid_113_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7411 = _T_66 ? _GEN_7154 : valid_114_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7412 = _T_66 ? _GEN_7155 : valid_114_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7413 = _T_66 ? _GEN_7156 : valid_115_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7414 = _T_66 ? _GEN_7157 : valid_115_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7415 = _T_66 ? _GEN_7158 : valid_116_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7416 = _T_66 ? _GEN_7159 : valid_116_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7417 = _T_66 ? _GEN_7160 : valid_117_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7418 = _T_66 ? _GEN_7161 : valid_117_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7419 = _T_66 ? _GEN_7162 : valid_118_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7420 = _T_66 ? _GEN_7163 : valid_118_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7421 = _T_66 ? _GEN_7164 : valid_119_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7422 = _T_66 ? _GEN_7165 : valid_119_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7423 = _T_66 ? _GEN_7166 : valid_120_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7424 = _T_66 ? _GEN_7167 : valid_120_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7425 = _T_66 ? _GEN_7168 : valid_121_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7426 = _T_66 ? _GEN_7169 : valid_121_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7427 = _T_66 ? _GEN_7170 : valid_122_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7428 = _T_66 ? _GEN_7171 : valid_122_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7429 = _T_66 ? _GEN_7172 : valid_123_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7430 = _T_66 ? _GEN_7173 : valid_123_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7431 = _T_66 ? _GEN_7174 : valid_124_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7432 = _T_66 ? _GEN_7175 : valid_124_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7433 = _T_66 ? _GEN_7176 : valid_125_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7434 = _T_66 ? _GEN_7177 : valid_125_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7435 = _T_66 ? _GEN_7178 : valid_126_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7436 = _T_66 ? _GEN_7179 : valid_126_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7437 = _T_66 ? _GEN_7180 : valid_127_0; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7438 = _T_66 ? _GEN_7181 : valid_127_1; // @[DCache.scala 486:13 68:22]
  wire  _GEN_7439 = ~bram_use_replace_addr ? 1'h0 : replace_working; // @[DCache.scala 490:40 491:29 98:40]
  wire [2:0] _GEN_7440 = ~bram_use_replace_addr ? 3'h0 : state; // @[DCache.scala 490:40 492:29 65:96]
  wire [9:0] _GEN_7441 = replace_working ? _GEN_6611 : _bram_replace_addr_T_4; // @[DCache.scala 419:31 498:29]
  wire [9:0] _GEN_7442 = replace_working ? _GEN_6612 : bram_read_ready_addr; // @[DCache.scala 419:31 91:40]
  wire [31:0] _GEN_7443 = replace_working ? _GEN_6613 : bram_r_buffer_0; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7444 = replace_working ? _GEN_6614 : bram_r_buffer_1; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7445 = replace_working ? _GEN_6615 : bram_r_buffer_2; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7446 = replace_working ? _GEN_6616 : bram_r_buffer_3; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7447 = replace_working ? _GEN_6617 : bram_r_buffer_4; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7448 = replace_working ? _GEN_6618 : bram_r_buffer_5; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7449 = replace_working ? _GEN_6619 : bram_r_buffer_6; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7450 = replace_working ? _GEN_6620 : bram_r_buffer_7; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7451 = replace_working ? _GEN_6621 : bram_r_buffer_8; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7452 = replace_working ? _GEN_6622 : bram_r_buffer_9; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7453 = replace_working ? _GEN_6623 : bram_r_buffer_10; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7454 = replace_working ? _GEN_6624 : bram_r_buffer_11; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7455 = replace_working ? _GEN_6625 : bram_r_buffer_12; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7456 = replace_working ? _GEN_6626 : bram_r_buffer_13; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7457 = replace_working ? _GEN_6627 : bram_r_buffer_14; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7458 = replace_working ? _GEN_6628 : bram_r_buffer_15; // @[DCache.scala 419:31 94:40]
  wire [31:0] _GEN_7459 = replace_working ? _GEN_6629 : _GEN_281; // @[DCache.scala 419:31]
  wire [7:0] _GEN_7460 = replace_working ? _GEN_6630 : _GEN_285; // @[DCache.scala 419:31]
  wire [2:0] _GEN_7461 = replace_working ? _GEN_6631 : _GEN_282; // @[DCache.scala 419:31]
  wire  _GEN_7462 = replace_working ? _GEN_6632 : _GEN_276; // @[DCache.scala 419:31]
  wire [31:0] _GEN_7463 = replace_working ? _GEN_6633 : _GEN_283; // @[DCache.scala 419:31]
  wire [3:0] _GEN_7464 = replace_working ? _GEN_6634 : _GEN_284; // @[DCache.scala 419:31]
  wire  _GEN_7465 = replace_working ? _GEN_6635 : _GEN_278; // @[DCache.scala 419:31]
  wire  _GEN_7466 = replace_working ? _GEN_6636 : _GEN_277; // @[DCache.scala 419:31]
  wire  _GEN_7467 = replace_working & _GEN_6637; // @[DCache.scala 419:31 496:29]
  wire [3:0] _GEN_7468 = replace_working ? _GEN_6638 : axi_wcnt; // @[DCache.scala 419:31 89:40]
  wire  _GEN_7469 = replace_working ? _GEN_6639 : dirty_0_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7470 = replace_working ? _GEN_6640 : dirty_0_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7471 = replace_working ? _GEN_6641 : dirty_1_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7472 = replace_working ? _GEN_6642 : dirty_1_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7473 = replace_working ? _GEN_6643 : dirty_2_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7474 = replace_working ? _GEN_6644 : dirty_2_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7475 = replace_working ? _GEN_6645 : dirty_3_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7476 = replace_working ? _GEN_6646 : dirty_3_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7477 = replace_working ? _GEN_6647 : dirty_4_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7478 = replace_working ? _GEN_6648 : dirty_4_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7479 = replace_working ? _GEN_6649 : dirty_5_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7480 = replace_working ? _GEN_6650 : dirty_5_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7481 = replace_working ? _GEN_6651 : dirty_6_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7482 = replace_working ? _GEN_6652 : dirty_6_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7483 = replace_working ? _GEN_6653 : dirty_7_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7484 = replace_working ? _GEN_6654 : dirty_7_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7485 = replace_working ? _GEN_6655 : dirty_8_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7486 = replace_working ? _GEN_6656 : dirty_8_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7487 = replace_working ? _GEN_6657 : dirty_9_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7488 = replace_working ? _GEN_6658 : dirty_9_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7489 = replace_working ? _GEN_6659 : dirty_10_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7490 = replace_working ? _GEN_6660 : dirty_10_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7491 = replace_working ? _GEN_6661 : dirty_11_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7492 = replace_working ? _GEN_6662 : dirty_11_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7493 = replace_working ? _GEN_6663 : dirty_12_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7494 = replace_working ? _GEN_6664 : dirty_12_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7495 = replace_working ? _GEN_6665 : dirty_13_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7496 = replace_working ? _GEN_6666 : dirty_13_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7497 = replace_working ? _GEN_6667 : dirty_14_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7498 = replace_working ? _GEN_6668 : dirty_14_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7499 = replace_working ? _GEN_6669 : dirty_15_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7500 = replace_working ? _GEN_6670 : dirty_15_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7501 = replace_working ? _GEN_6671 : dirty_16_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7502 = replace_working ? _GEN_6672 : dirty_16_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7503 = replace_working ? _GEN_6673 : dirty_17_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7504 = replace_working ? _GEN_6674 : dirty_17_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7505 = replace_working ? _GEN_6675 : dirty_18_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7506 = replace_working ? _GEN_6676 : dirty_18_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7507 = replace_working ? _GEN_6677 : dirty_19_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7508 = replace_working ? _GEN_6678 : dirty_19_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7509 = replace_working ? _GEN_6679 : dirty_20_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7510 = replace_working ? _GEN_6680 : dirty_20_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7511 = replace_working ? _GEN_6681 : dirty_21_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7512 = replace_working ? _GEN_6682 : dirty_21_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7513 = replace_working ? _GEN_6683 : dirty_22_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7514 = replace_working ? _GEN_6684 : dirty_22_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7515 = replace_working ? _GEN_6685 : dirty_23_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7516 = replace_working ? _GEN_6686 : dirty_23_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7517 = replace_working ? _GEN_6687 : dirty_24_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7518 = replace_working ? _GEN_6688 : dirty_24_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7519 = replace_working ? _GEN_6689 : dirty_25_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7520 = replace_working ? _GEN_6690 : dirty_25_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7521 = replace_working ? _GEN_6691 : dirty_26_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7522 = replace_working ? _GEN_6692 : dirty_26_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7523 = replace_working ? _GEN_6693 : dirty_27_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7524 = replace_working ? _GEN_6694 : dirty_27_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7525 = replace_working ? _GEN_6695 : dirty_28_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7526 = replace_working ? _GEN_6696 : dirty_28_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7527 = replace_working ? _GEN_6697 : dirty_29_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7528 = replace_working ? _GEN_6698 : dirty_29_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7529 = replace_working ? _GEN_6699 : dirty_30_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7530 = replace_working ? _GEN_6700 : dirty_30_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7531 = replace_working ? _GEN_6701 : dirty_31_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7532 = replace_working ? _GEN_6702 : dirty_31_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7533 = replace_working ? _GEN_6703 : dirty_32_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7534 = replace_working ? _GEN_6704 : dirty_32_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7535 = replace_working ? _GEN_6705 : dirty_33_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7536 = replace_working ? _GEN_6706 : dirty_33_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7537 = replace_working ? _GEN_6707 : dirty_34_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7538 = replace_working ? _GEN_6708 : dirty_34_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7539 = replace_working ? _GEN_6709 : dirty_35_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7540 = replace_working ? _GEN_6710 : dirty_35_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7541 = replace_working ? _GEN_6711 : dirty_36_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7542 = replace_working ? _GEN_6712 : dirty_36_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7543 = replace_working ? _GEN_6713 : dirty_37_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7544 = replace_working ? _GEN_6714 : dirty_37_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7545 = replace_working ? _GEN_6715 : dirty_38_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7546 = replace_working ? _GEN_6716 : dirty_38_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7547 = replace_working ? _GEN_6717 : dirty_39_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7548 = replace_working ? _GEN_6718 : dirty_39_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7549 = replace_working ? _GEN_6719 : dirty_40_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7550 = replace_working ? _GEN_6720 : dirty_40_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7551 = replace_working ? _GEN_6721 : dirty_41_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7552 = replace_working ? _GEN_6722 : dirty_41_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7553 = replace_working ? _GEN_6723 : dirty_42_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7554 = replace_working ? _GEN_6724 : dirty_42_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7555 = replace_working ? _GEN_6725 : dirty_43_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7556 = replace_working ? _GEN_6726 : dirty_43_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7557 = replace_working ? _GEN_6727 : dirty_44_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7558 = replace_working ? _GEN_6728 : dirty_44_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7559 = replace_working ? _GEN_6729 : dirty_45_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7560 = replace_working ? _GEN_6730 : dirty_45_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7561 = replace_working ? _GEN_6731 : dirty_46_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7562 = replace_working ? _GEN_6732 : dirty_46_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7563 = replace_working ? _GEN_6733 : dirty_47_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7564 = replace_working ? _GEN_6734 : dirty_47_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7565 = replace_working ? _GEN_6735 : dirty_48_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7566 = replace_working ? _GEN_6736 : dirty_48_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7567 = replace_working ? _GEN_6737 : dirty_49_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7568 = replace_working ? _GEN_6738 : dirty_49_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7569 = replace_working ? _GEN_6739 : dirty_50_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7570 = replace_working ? _GEN_6740 : dirty_50_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7571 = replace_working ? _GEN_6741 : dirty_51_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7572 = replace_working ? _GEN_6742 : dirty_51_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7573 = replace_working ? _GEN_6743 : dirty_52_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7574 = replace_working ? _GEN_6744 : dirty_52_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7575 = replace_working ? _GEN_6745 : dirty_53_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7576 = replace_working ? _GEN_6746 : dirty_53_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7577 = replace_working ? _GEN_6747 : dirty_54_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7578 = replace_working ? _GEN_6748 : dirty_54_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7579 = replace_working ? _GEN_6749 : dirty_55_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7580 = replace_working ? _GEN_6750 : dirty_55_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7581 = replace_working ? _GEN_6751 : dirty_56_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7582 = replace_working ? _GEN_6752 : dirty_56_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7583 = replace_working ? _GEN_6753 : dirty_57_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7584 = replace_working ? _GEN_6754 : dirty_57_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7585 = replace_working ? _GEN_6755 : dirty_58_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7586 = replace_working ? _GEN_6756 : dirty_58_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7587 = replace_working ? _GEN_6757 : dirty_59_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7588 = replace_working ? _GEN_6758 : dirty_59_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7589 = replace_working ? _GEN_6759 : dirty_60_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7590 = replace_working ? _GEN_6760 : dirty_60_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7591 = replace_working ? _GEN_6761 : dirty_61_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7592 = replace_working ? _GEN_6762 : dirty_61_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7593 = replace_working ? _GEN_6763 : dirty_62_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7594 = replace_working ? _GEN_6764 : dirty_62_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7595 = replace_working ? _GEN_6765 : dirty_63_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7596 = replace_working ? _GEN_6766 : dirty_63_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7597 = replace_working ? _GEN_6767 : dirty_64_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7598 = replace_working ? _GEN_6768 : dirty_64_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7599 = replace_working ? _GEN_6769 : dirty_65_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7600 = replace_working ? _GEN_6770 : dirty_65_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7601 = replace_working ? _GEN_6771 : dirty_66_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7602 = replace_working ? _GEN_6772 : dirty_66_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7603 = replace_working ? _GEN_6773 : dirty_67_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7604 = replace_working ? _GEN_6774 : dirty_67_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7605 = replace_working ? _GEN_6775 : dirty_68_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7606 = replace_working ? _GEN_6776 : dirty_68_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7607 = replace_working ? _GEN_6777 : dirty_69_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7608 = replace_working ? _GEN_6778 : dirty_69_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7609 = replace_working ? _GEN_6779 : dirty_70_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7610 = replace_working ? _GEN_6780 : dirty_70_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7611 = replace_working ? _GEN_6781 : dirty_71_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7612 = replace_working ? _GEN_6782 : dirty_71_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7613 = replace_working ? _GEN_6783 : dirty_72_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7614 = replace_working ? _GEN_6784 : dirty_72_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7615 = replace_working ? _GEN_6785 : dirty_73_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7616 = replace_working ? _GEN_6786 : dirty_73_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7617 = replace_working ? _GEN_6787 : dirty_74_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7618 = replace_working ? _GEN_6788 : dirty_74_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7619 = replace_working ? _GEN_6789 : dirty_75_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7620 = replace_working ? _GEN_6790 : dirty_75_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7621 = replace_working ? _GEN_6791 : dirty_76_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7622 = replace_working ? _GEN_6792 : dirty_76_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7623 = replace_working ? _GEN_6793 : dirty_77_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7624 = replace_working ? _GEN_6794 : dirty_77_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7625 = replace_working ? _GEN_6795 : dirty_78_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7626 = replace_working ? _GEN_6796 : dirty_78_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7627 = replace_working ? _GEN_6797 : dirty_79_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7628 = replace_working ? _GEN_6798 : dirty_79_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7629 = replace_working ? _GEN_6799 : dirty_80_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7630 = replace_working ? _GEN_6800 : dirty_80_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7631 = replace_working ? _GEN_6801 : dirty_81_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7632 = replace_working ? _GEN_6802 : dirty_81_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7633 = replace_working ? _GEN_6803 : dirty_82_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7634 = replace_working ? _GEN_6804 : dirty_82_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7635 = replace_working ? _GEN_6805 : dirty_83_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7636 = replace_working ? _GEN_6806 : dirty_83_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7637 = replace_working ? _GEN_6807 : dirty_84_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7638 = replace_working ? _GEN_6808 : dirty_84_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7639 = replace_working ? _GEN_6809 : dirty_85_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7640 = replace_working ? _GEN_6810 : dirty_85_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7641 = replace_working ? _GEN_6811 : dirty_86_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7642 = replace_working ? _GEN_6812 : dirty_86_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7643 = replace_working ? _GEN_6813 : dirty_87_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7644 = replace_working ? _GEN_6814 : dirty_87_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7645 = replace_working ? _GEN_6815 : dirty_88_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7646 = replace_working ? _GEN_6816 : dirty_88_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7647 = replace_working ? _GEN_6817 : dirty_89_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7648 = replace_working ? _GEN_6818 : dirty_89_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7649 = replace_working ? _GEN_6819 : dirty_90_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7650 = replace_working ? _GEN_6820 : dirty_90_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7651 = replace_working ? _GEN_6821 : dirty_91_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7652 = replace_working ? _GEN_6822 : dirty_91_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7653 = replace_working ? _GEN_6823 : dirty_92_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7654 = replace_working ? _GEN_6824 : dirty_92_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7655 = replace_working ? _GEN_6825 : dirty_93_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7656 = replace_working ? _GEN_6826 : dirty_93_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7657 = replace_working ? _GEN_6827 : dirty_94_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7658 = replace_working ? _GEN_6828 : dirty_94_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7659 = replace_working ? _GEN_6829 : dirty_95_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7660 = replace_working ? _GEN_6830 : dirty_95_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7661 = replace_working ? _GEN_6831 : dirty_96_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7662 = replace_working ? _GEN_6832 : dirty_96_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7663 = replace_working ? _GEN_6833 : dirty_97_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7664 = replace_working ? _GEN_6834 : dirty_97_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7665 = replace_working ? _GEN_6835 : dirty_98_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7666 = replace_working ? _GEN_6836 : dirty_98_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7667 = replace_working ? _GEN_6837 : dirty_99_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7668 = replace_working ? _GEN_6838 : dirty_99_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7669 = replace_working ? _GEN_6839 : dirty_100_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7670 = replace_working ? _GEN_6840 : dirty_100_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7671 = replace_working ? _GEN_6841 : dirty_101_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7672 = replace_working ? _GEN_6842 : dirty_101_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7673 = replace_working ? _GEN_6843 : dirty_102_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7674 = replace_working ? _GEN_6844 : dirty_102_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7675 = replace_working ? _GEN_6845 : dirty_103_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7676 = replace_working ? _GEN_6846 : dirty_103_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7677 = replace_working ? _GEN_6847 : dirty_104_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7678 = replace_working ? _GEN_6848 : dirty_104_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7679 = replace_working ? _GEN_6849 : dirty_105_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7680 = replace_working ? _GEN_6850 : dirty_105_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7681 = replace_working ? _GEN_6851 : dirty_106_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7682 = replace_working ? _GEN_6852 : dirty_106_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7683 = replace_working ? _GEN_6853 : dirty_107_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7684 = replace_working ? _GEN_6854 : dirty_107_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7685 = replace_working ? _GEN_6855 : dirty_108_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7686 = replace_working ? _GEN_6856 : dirty_108_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7687 = replace_working ? _GEN_6857 : dirty_109_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7688 = replace_working ? _GEN_6858 : dirty_109_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7689 = replace_working ? _GEN_6859 : dirty_110_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7690 = replace_working ? _GEN_6860 : dirty_110_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7691 = replace_working ? _GEN_6861 : dirty_111_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7692 = replace_working ? _GEN_6862 : dirty_111_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7693 = replace_working ? _GEN_6863 : dirty_112_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7694 = replace_working ? _GEN_6864 : dirty_112_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7695 = replace_working ? _GEN_6865 : dirty_113_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7696 = replace_working ? _GEN_6866 : dirty_113_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7697 = replace_working ? _GEN_6867 : dirty_114_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7698 = replace_working ? _GEN_6868 : dirty_114_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7699 = replace_working ? _GEN_6869 : dirty_115_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7700 = replace_working ? _GEN_6870 : dirty_115_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7701 = replace_working ? _GEN_6871 : dirty_116_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7702 = replace_working ? _GEN_6872 : dirty_116_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7703 = replace_working ? _GEN_6873 : dirty_117_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7704 = replace_working ? _GEN_6874 : dirty_117_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7705 = replace_working ? _GEN_6875 : dirty_118_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7706 = replace_working ? _GEN_6876 : dirty_118_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7707 = replace_working ? _GEN_6877 : dirty_119_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7708 = replace_working ? _GEN_6878 : dirty_119_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7709 = replace_working ? _GEN_6879 : dirty_120_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7710 = replace_working ? _GEN_6880 : dirty_120_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7711 = replace_working ? _GEN_6881 : dirty_121_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7712 = replace_working ? _GEN_6882 : dirty_121_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7713 = replace_working ? _GEN_6883 : dirty_122_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7714 = replace_working ? _GEN_6884 : dirty_122_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7715 = replace_working ? _GEN_6885 : dirty_123_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7716 = replace_working ? _GEN_6886 : dirty_123_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7717 = replace_working ? _GEN_6887 : dirty_124_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7718 = replace_working ? _GEN_6888 : dirty_124_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7719 = replace_working ? _GEN_6889 : dirty_125_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7720 = replace_working ? _GEN_6890 : dirty_125_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7721 = replace_working ? _GEN_6891 : dirty_126_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7722 = replace_working ? _GEN_6892 : dirty_126_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7723 = replace_working ? _GEN_6893 : dirty_127_0; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7724 = replace_working ? _GEN_6894 : dirty_127_1; // @[DCache.scala 419:31 69:22]
  wire  _GEN_7725 = replace_working ? _GEN_6895 : replace_writeback; // @[DCache.scala 419:31 101:40]
  wire [31:0] _GEN_7726 = replace_working ? _GEN_6900 : ar_addr; // @[DCache.scala 199:24 419:31]
  wire [7:0] _GEN_7727 = replace_working ? _GEN_6901 : ar_len; // @[DCache.scala 199:24 419:31]
  wire [2:0] _GEN_7728 = replace_working ? _GEN_6902 : ar_size; // @[DCache.scala 199:24 419:31]
  wire  _GEN_7729 = replace_working ? _GEN_6915 : arvalid; // @[DCache.scala 200:24 419:31]
  wire  _GEN_7730 = replace_working ? _GEN_6922 : rready; // @[DCache.scala 203:23 419:31]
  wire  _GEN_7731 = replace_working & _GEN_6905; // @[DCache.scala 419:31 495:29]
  wire [3:0] _GEN_7732 = replace_working ? _GEN_6923 : bram_replace_wea_0; // @[DCache.scala 419:31 73:33]
  wire [3:0] _GEN_7733 = replace_working ? _GEN_6924 : bram_replace_wea_1; // @[DCache.scala 419:31 73:33]
  wire  _GEN_7734 = replace_working ? _GEN_6913 : tag_wstrb_0; // @[DCache.scala 419:31 72:33]
  wire  _GEN_7735 = replace_working ? _GEN_6914 : tag_wstrb_1; // @[DCache.scala 419:31 72:33]
  wire [19:0] _GEN_7736 = replace_working ? _GEN_6910 : tag_wdata; // @[DCache.scala 419:31 77:26]
  wire [9:0] _GEN_7737 = replace_working ? _GEN_6925 : bram_replace_write_addr; // @[DCache.scala 419:31 92:40]
  wire  _GEN_7738 = replace_working ? _GEN_7182 : bram_use_replace_addr; // @[DCache.scala 419:31 95:40]
  wire  _GEN_7739 = replace_working ? _GEN_7183 : valid_0_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7740 = replace_working ? _GEN_7184 : valid_0_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7741 = replace_working ? _GEN_7185 : valid_1_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7742 = replace_working ? _GEN_7186 : valid_1_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7743 = replace_working ? _GEN_7187 : valid_2_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7744 = replace_working ? _GEN_7188 : valid_2_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7745 = replace_working ? _GEN_7189 : valid_3_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7746 = replace_working ? _GEN_7190 : valid_3_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7747 = replace_working ? _GEN_7191 : valid_4_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7748 = replace_working ? _GEN_7192 : valid_4_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7749 = replace_working ? _GEN_7193 : valid_5_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7750 = replace_working ? _GEN_7194 : valid_5_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7751 = replace_working ? _GEN_7195 : valid_6_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7752 = replace_working ? _GEN_7196 : valid_6_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7753 = replace_working ? _GEN_7197 : valid_7_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7754 = replace_working ? _GEN_7198 : valid_7_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7755 = replace_working ? _GEN_7199 : valid_8_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7756 = replace_working ? _GEN_7200 : valid_8_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7757 = replace_working ? _GEN_7201 : valid_9_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7758 = replace_working ? _GEN_7202 : valid_9_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7759 = replace_working ? _GEN_7203 : valid_10_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7760 = replace_working ? _GEN_7204 : valid_10_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7761 = replace_working ? _GEN_7205 : valid_11_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7762 = replace_working ? _GEN_7206 : valid_11_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7763 = replace_working ? _GEN_7207 : valid_12_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7764 = replace_working ? _GEN_7208 : valid_12_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7765 = replace_working ? _GEN_7209 : valid_13_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7766 = replace_working ? _GEN_7210 : valid_13_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7767 = replace_working ? _GEN_7211 : valid_14_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7768 = replace_working ? _GEN_7212 : valid_14_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7769 = replace_working ? _GEN_7213 : valid_15_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7770 = replace_working ? _GEN_7214 : valid_15_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7771 = replace_working ? _GEN_7215 : valid_16_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7772 = replace_working ? _GEN_7216 : valid_16_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7773 = replace_working ? _GEN_7217 : valid_17_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7774 = replace_working ? _GEN_7218 : valid_17_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7775 = replace_working ? _GEN_7219 : valid_18_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7776 = replace_working ? _GEN_7220 : valid_18_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7777 = replace_working ? _GEN_7221 : valid_19_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7778 = replace_working ? _GEN_7222 : valid_19_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7779 = replace_working ? _GEN_7223 : valid_20_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7780 = replace_working ? _GEN_7224 : valid_20_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7781 = replace_working ? _GEN_7225 : valid_21_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7782 = replace_working ? _GEN_7226 : valid_21_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7783 = replace_working ? _GEN_7227 : valid_22_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7784 = replace_working ? _GEN_7228 : valid_22_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7785 = replace_working ? _GEN_7229 : valid_23_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7786 = replace_working ? _GEN_7230 : valid_23_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7787 = replace_working ? _GEN_7231 : valid_24_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7788 = replace_working ? _GEN_7232 : valid_24_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7789 = replace_working ? _GEN_7233 : valid_25_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7790 = replace_working ? _GEN_7234 : valid_25_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7791 = replace_working ? _GEN_7235 : valid_26_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7792 = replace_working ? _GEN_7236 : valid_26_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7793 = replace_working ? _GEN_7237 : valid_27_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7794 = replace_working ? _GEN_7238 : valid_27_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7795 = replace_working ? _GEN_7239 : valid_28_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7796 = replace_working ? _GEN_7240 : valid_28_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7797 = replace_working ? _GEN_7241 : valid_29_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7798 = replace_working ? _GEN_7242 : valid_29_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7799 = replace_working ? _GEN_7243 : valid_30_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7800 = replace_working ? _GEN_7244 : valid_30_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7801 = replace_working ? _GEN_7245 : valid_31_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7802 = replace_working ? _GEN_7246 : valid_31_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7803 = replace_working ? _GEN_7247 : valid_32_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7804 = replace_working ? _GEN_7248 : valid_32_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7805 = replace_working ? _GEN_7249 : valid_33_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7806 = replace_working ? _GEN_7250 : valid_33_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7807 = replace_working ? _GEN_7251 : valid_34_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7808 = replace_working ? _GEN_7252 : valid_34_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7809 = replace_working ? _GEN_7253 : valid_35_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7810 = replace_working ? _GEN_7254 : valid_35_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7811 = replace_working ? _GEN_7255 : valid_36_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7812 = replace_working ? _GEN_7256 : valid_36_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7813 = replace_working ? _GEN_7257 : valid_37_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7814 = replace_working ? _GEN_7258 : valid_37_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7815 = replace_working ? _GEN_7259 : valid_38_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7816 = replace_working ? _GEN_7260 : valid_38_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7817 = replace_working ? _GEN_7261 : valid_39_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7818 = replace_working ? _GEN_7262 : valid_39_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7819 = replace_working ? _GEN_7263 : valid_40_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7820 = replace_working ? _GEN_7264 : valid_40_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7821 = replace_working ? _GEN_7265 : valid_41_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7822 = replace_working ? _GEN_7266 : valid_41_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7823 = replace_working ? _GEN_7267 : valid_42_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7824 = replace_working ? _GEN_7268 : valid_42_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7825 = replace_working ? _GEN_7269 : valid_43_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7826 = replace_working ? _GEN_7270 : valid_43_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7827 = replace_working ? _GEN_7271 : valid_44_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7828 = replace_working ? _GEN_7272 : valid_44_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7829 = replace_working ? _GEN_7273 : valid_45_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7830 = replace_working ? _GEN_7274 : valid_45_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7831 = replace_working ? _GEN_7275 : valid_46_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7832 = replace_working ? _GEN_7276 : valid_46_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7833 = replace_working ? _GEN_7277 : valid_47_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7834 = replace_working ? _GEN_7278 : valid_47_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7835 = replace_working ? _GEN_7279 : valid_48_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7836 = replace_working ? _GEN_7280 : valid_48_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7837 = replace_working ? _GEN_7281 : valid_49_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7838 = replace_working ? _GEN_7282 : valid_49_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7839 = replace_working ? _GEN_7283 : valid_50_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7840 = replace_working ? _GEN_7284 : valid_50_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7841 = replace_working ? _GEN_7285 : valid_51_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7842 = replace_working ? _GEN_7286 : valid_51_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7843 = replace_working ? _GEN_7287 : valid_52_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7844 = replace_working ? _GEN_7288 : valid_52_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7845 = replace_working ? _GEN_7289 : valid_53_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7846 = replace_working ? _GEN_7290 : valid_53_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7847 = replace_working ? _GEN_7291 : valid_54_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7848 = replace_working ? _GEN_7292 : valid_54_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7849 = replace_working ? _GEN_7293 : valid_55_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7850 = replace_working ? _GEN_7294 : valid_55_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7851 = replace_working ? _GEN_7295 : valid_56_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7852 = replace_working ? _GEN_7296 : valid_56_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7853 = replace_working ? _GEN_7297 : valid_57_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7854 = replace_working ? _GEN_7298 : valid_57_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7855 = replace_working ? _GEN_7299 : valid_58_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7856 = replace_working ? _GEN_7300 : valid_58_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7857 = replace_working ? _GEN_7301 : valid_59_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7858 = replace_working ? _GEN_7302 : valid_59_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7859 = replace_working ? _GEN_7303 : valid_60_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7860 = replace_working ? _GEN_7304 : valid_60_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7861 = replace_working ? _GEN_7305 : valid_61_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7862 = replace_working ? _GEN_7306 : valid_61_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7863 = replace_working ? _GEN_7307 : valid_62_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7864 = replace_working ? _GEN_7308 : valid_62_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7865 = replace_working ? _GEN_7309 : valid_63_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7866 = replace_working ? _GEN_7310 : valid_63_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7867 = replace_working ? _GEN_7311 : valid_64_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7868 = replace_working ? _GEN_7312 : valid_64_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7869 = replace_working ? _GEN_7313 : valid_65_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7870 = replace_working ? _GEN_7314 : valid_65_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7871 = replace_working ? _GEN_7315 : valid_66_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7872 = replace_working ? _GEN_7316 : valid_66_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7873 = replace_working ? _GEN_7317 : valid_67_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7874 = replace_working ? _GEN_7318 : valid_67_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7875 = replace_working ? _GEN_7319 : valid_68_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7876 = replace_working ? _GEN_7320 : valid_68_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7877 = replace_working ? _GEN_7321 : valid_69_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7878 = replace_working ? _GEN_7322 : valid_69_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7879 = replace_working ? _GEN_7323 : valid_70_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7880 = replace_working ? _GEN_7324 : valid_70_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7881 = replace_working ? _GEN_7325 : valid_71_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7882 = replace_working ? _GEN_7326 : valid_71_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7883 = replace_working ? _GEN_7327 : valid_72_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7884 = replace_working ? _GEN_7328 : valid_72_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7885 = replace_working ? _GEN_7329 : valid_73_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7886 = replace_working ? _GEN_7330 : valid_73_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7887 = replace_working ? _GEN_7331 : valid_74_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7888 = replace_working ? _GEN_7332 : valid_74_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7889 = replace_working ? _GEN_7333 : valid_75_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7890 = replace_working ? _GEN_7334 : valid_75_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7891 = replace_working ? _GEN_7335 : valid_76_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7892 = replace_working ? _GEN_7336 : valid_76_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7893 = replace_working ? _GEN_7337 : valid_77_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7894 = replace_working ? _GEN_7338 : valid_77_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7895 = replace_working ? _GEN_7339 : valid_78_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7896 = replace_working ? _GEN_7340 : valid_78_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7897 = replace_working ? _GEN_7341 : valid_79_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7898 = replace_working ? _GEN_7342 : valid_79_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7899 = replace_working ? _GEN_7343 : valid_80_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7900 = replace_working ? _GEN_7344 : valid_80_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7901 = replace_working ? _GEN_7345 : valid_81_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7902 = replace_working ? _GEN_7346 : valid_81_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7903 = replace_working ? _GEN_7347 : valid_82_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7904 = replace_working ? _GEN_7348 : valid_82_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7905 = replace_working ? _GEN_7349 : valid_83_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7906 = replace_working ? _GEN_7350 : valid_83_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7907 = replace_working ? _GEN_7351 : valid_84_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7908 = replace_working ? _GEN_7352 : valid_84_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7909 = replace_working ? _GEN_7353 : valid_85_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7910 = replace_working ? _GEN_7354 : valid_85_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7911 = replace_working ? _GEN_7355 : valid_86_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7912 = replace_working ? _GEN_7356 : valid_86_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7913 = replace_working ? _GEN_7357 : valid_87_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7914 = replace_working ? _GEN_7358 : valid_87_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7915 = replace_working ? _GEN_7359 : valid_88_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7916 = replace_working ? _GEN_7360 : valid_88_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7917 = replace_working ? _GEN_7361 : valid_89_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7918 = replace_working ? _GEN_7362 : valid_89_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7919 = replace_working ? _GEN_7363 : valid_90_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7920 = replace_working ? _GEN_7364 : valid_90_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7921 = replace_working ? _GEN_7365 : valid_91_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7922 = replace_working ? _GEN_7366 : valid_91_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7923 = replace_working ? _GEN_7367 : valid_92_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7924 = replace_working ? _GEN_7368 : valid_92_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7925 = replace_working ? _GEN_7369 : valid_93_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7926 = replace_working ? _GEN_7370 : valid_93_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7927 = replace_working ? _GEN_7371 : valid_94_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7928 = replace_working ? _GEN_7372 : valid_94_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7929 = replace_working ? _GEN_7373 : valid_95_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7930 = replace_working ? _GEN_7374 : valid_95_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7931 = replace_working ? _GEN_7375 : valid_96_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7932 = replace_working ? _GEN_7376 : valid_96_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7933 = replace_working ? _GEN_7377 : valid_97_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7934 = replace_working ? _GEN_7378 : valid_97_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7935 = replace_working ? _GEN_7379 : valid_98_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7936 = replace_working ? _GEN_7380 : valid_98_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7937 = replace_working ? _GEN_7381 : valid_99_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7938 = replace_working ? _GEN_7382 : valid_99_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7939 = replace_working ? _GEN_7383 : valid_100_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7940 = replace_working ? _GEN_7384 : valid_100_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7941 = replace_working ? _GEN_7385 : valid_101_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7942 = replace_working ? _GEN_7386 : valid_101_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7943 = replace_working ? _GEN_7387 : valid_102_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7944 = replace_working ? _GEN_7388 : valid_102_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7945 = replace_working ? _GEN_7389 : valid_103_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7946 = replace_working ? _GEN_7390 : valid_103_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7947 = replace_working ? _GEN_7391 : valid_104_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7948 = replace_working ? _GEN_7392 : valid_104_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7949 = replace_working ? _GEN_7393 : valid_105_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7950 = replace_working ? _GEN_7394 : valid_105_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7951 = replace_working ? _GEN_7395 : valid_106_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7952 = replace_working ? _GEN_7396 : valid_106_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7953 = replace_working ? _GEN_7397 : valid_107_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7954 = replace_working ? _GEN_7398 : valid_107_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7955 = replace_working ? _GEN_7399 : valid_108_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7956 = replace_working ? _GEN_7400 : valid_108_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7957 = replace_working ? _GEN_7401 : valid_109_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7958 = replace_working ? _GEN_7402 : valid_109_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7959 = replace_working ? _GEN_7403 : valid_110_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7960 = replace_working ? _GEN_7404 : valid_110_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7961 = replace_working ? _GEN_7405 : valid_111_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7962 = replace_working ? _GEN_7406 : valid_111_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7963 = replace_working ? _GEN_7407 : valid_112_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7964 = replace_working ? _GEN_7408 : valid_112_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7965 = replace_working ? _GEN_7409 : valid_113_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7966 = replace_working ? _GEN_7410 : valid_113_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7967 = replace_working ? _GEN_7411 : valid_114_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7968 = replace_working ? _GEN_7412 : valid_114_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7969 = replace_working ? _GEN_7413 : valid_115_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7970 = replace_working ? _GEN_7414 : valid_115_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7971 = replace_working ? _GEN_7415 : valid_116_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7972 = replace_working ? _GEN_7416 : valid_116_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7973 = replace_working ? _GEN_7417 : valid_117_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7974 = replace_working ? _GEN_7418 : valid_117_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7975 = replace_working ? _GEN_7419 : valid_118_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7976 = replace_working ? _GEN_7420 : valid_118_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7977 = replace_working ? _GEN_7421 : valid_119_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7978 = replace_working ? _GEN_7422 : valid_119_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7979 = replace_working ? _GEN_7423 : valid_120_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7980 = replace_working ? _GEN_7424 : valid_120_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7981 = replace_working ? _GEN_7425 : valid_121_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7982 = replace_working ? _GEN_7426 : valid_121_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7983 = replace_working ? _GEN_7427 : valid_122_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7984 = replace_working ? _GEN_7428 : valid_122_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7985 = replace_working ? _GEN_7429 : valid_123_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7986 = replace_working ? _GEN_7430 : valid_123_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7987 = replace_working ? _GEN_7431 : valid_124_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7988 = replace_working ? _GEN_7432 : valid_124_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7989 = replace_working ? _GEN_7433 : valid_125_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7990 = replace_working ? _GEN_7434 : valid_125_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7991 = replace_working ? _GEN_7435 : valid_126_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7992 = replace_working ? _GEN_7436 : valid_126_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7993 = replace_working ? _GEN_7437 : valid_127_0; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7994 = replace_working ? _GEN_7438 : valid_127_1; // @[DCache.scala 419:31 68:22]
  wire  _GEN_7995 = replace_working ? _GEN_7439 : 1'h1; // @[DCache.scala 419:31 497:29]
  wire [2:0] _GEN_7996 = replace_working ? _GEN_7440 : state; // @[DCache.scala 419:31 65:96]
  wire [9:0] _GEN_7997 = _T_12 ? _GEN_7441 : bram_replace_addr; // @[DCache.scala 418:67 90:40]
  wire [9:0] _GEN_7998 = _T_12 ? _GEN_7442 : bram_read_ready_addr; // @[DCache.scala 418:67 91:40]
  wire [31:0] _GEN_7999 = _T_12 ? _GEN_7443 : bram_r_buffer_0; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8000 = _T_12 ? _GEN_7444 : bram_r_buffer_1; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8001 = _T_12 ? _GEN_7445 : bram_r_buffer_2; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8002 = _T_12 ? _GEN_7446 : bram_r_buffer_3; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8003 = _T_12 ? _GEN_7447 : bram_r_buffer_4; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8004 = _T_12 ? _GEN_7448 : bram_r_buffer_5; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8005 = _T_12 ? _GEN_7449 : bram_r_buffer_6; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8006 = _T_12 ? _GEN_7450 : bram_r_buffer_7; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8007 = _T_12 ? _GEN_7451 : bram_r_buffer_8; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8008 = _T_12 ? _GEN_7452 : bram_r_buffer_9; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8009 = _T_12 ? _GEN_7453 : bram_r_buffer_10; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8010 = _T_12 ? _GEN_7454 : bram_r_buffer_11; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8011 = _T_12 ? _GEN_7455 : bram_r_buffer_12; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8012 = _T_12 ? _GEN_7456 : bram_r_buffer_13; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8013 = _T_12 ? _GEN_7457 : bram_r_buffer_14; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8014 = _T_12 ? _GEN_7458 : bram_r_buffer_15; // @[DCache.scala 418:67 94:40]
  wire [31:0] _GEN_8015 = _T_12 ? _GEN_7459 : _GEN_281; // @[DCache.scala 418:67]
  wire [7:0] _GEN_8016 = _T_12 ? _GEN_7460 : _GEN_285; // @[DCache.scala 418:67]
  wire [2:0] _GEN_8017 = _T_12 ? _GEN_7461 : _GEN_282; // @[DCache.scala 418:67]
  wire  _GEN_8018 = _T_12 ? _GEN_7462 : _GEN_276; // @[DCache.scala 418:67]
  wire [31:0] _GEN_8019 = _T_12 ? _GEN_7463 : _GEN_283; // @[DCache.scala 418:67]
  wire [3:0] _GEN_8020 = _T_12 ? _GEN_7464 : _GEN_284; // @[DCache.scala 418:67]
  wire  _GEN_8021 = _T_12 ? _GEN_7465 : _GEN_278; // @[DCache.scala 418:67]
  wire  _GEN_8022 = _T_12 ? _GEN_7466 : _GEN_277; // @[DCache.scala 418:67]
  wire  _GEN_8023 = _T_12 ? _GEN_7467 : aw_handshake; // @[DCache.scala 100:40 418:67]
  wire [3:0] _GEN_8024 = _T_12 ? _GEN_7468 : axi_wcnt; // @[DCache.scala 418:67 89:40]
  wire  _GEN_8025 = _T_12 ? _GEN_7469 : dirty_0_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8026 = _T_12 ? _GEN_7470 : dirty_0_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8027 = _T_12 ? _GEN_7471 : dirty_1_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8028 = _T_12 ? _GEN_7472 : dirty_1_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8029 = _T_12 ? _GEN_7473 : dirty_2_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8030 = _T_12 ? _GEN_7474 : dirty_2_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8031 = _T_12 ? _GEN_7475 : dirty_3_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8032 = _T_12 ? _GEN_7476 : dirty_3_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8033 = _T_12 ? _GEN_7477 : dirty_4_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8034 = _T_12 ? _GEN_7478 : dirty_4_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8035 = _T_12 ? _GEN_7479 : dirty_5_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8036 = _T_12 ? _GEN_7480 : dirty_5_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8037 = _T_12 ? _GEN_7481 : dirty_6_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8038 = _T_12 ? _GEN_7482 : dirty_6_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8039 = _T_12 ? _GEN_7483 : dirty_7_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8040 = _T_12 ? _GEN_7484 : dirty_7_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8041 = _T_12 ? _GEN_7485 : dirty_8_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8042 = _T_12 ? _GEN_7486 : dirty_8_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8043 = _T_12 ? _GEN_7487 : dirty_9_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8044 = _T_12 ? _GEN_7488 : dirty_9_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8045 = _T_12 ? _GEN_7489 : dirty_10_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8046 = _T_12 ? _GEN_7490 : dirty_10_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8047 = _T_12 ? _GEN_7491 : dirty_11_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8048 = _T_12 ? _GEN_7492 : dirty_11_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8049 = _T_12 ? _GEN_7493 : dirty_12_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8050 = _T_12 ? _GEN_7494 : dirty_12_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8051 = _T_12 ? _GEN_7495 : dirty_13_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8052 = _T_12 ? _GEN_7496 : dirty_13_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8053 = _T_12 ? _GEN_7497 : dirty_14_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8054 = _T_12 ? _GEN_7498 : dirty_14_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8055 = _T_12 ? _GEN_7499 : dirty_15_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8056 = _T_12 ? _GEN_7500 : dirty_15_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8057 = _T_12 ? _GEN_7501 : dirty_16_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8058 = _T_12 ? _GEN_7502 : dirty_16_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8059 = _T_12 ? _GEN_7503 : dirty_17_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8060 = _T_12 ? _GEN_7504 : dirty_17_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8061 = _T_12 ? _GEN_7505 : dirty_18_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8062 = _T_12 ? _GEN_7506 : dirty_18_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8063 = _T_12 ? _GEN_7507 : dirty_19_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8064 = _T_12 ? _GEN_7508 : dirty_19_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8065 = _T_12 ? _GEN_7509 : dirty_20_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8066 = _T_12 ? _GEN_7510 : dirty_20_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8067 = _T_12 ? _GEN_7511 : dirty_21_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8068 = _T_12 ? _GEN_7512 : dirty_21_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8069 = _T_12 ? _GEN_7513 : dirty_22_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8070 = _T_12 ? _GEN_7514 : dirty_22_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8071 = _T_12 ? _GEN_7515 : dirty_23_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8072 = _T_12 ? _GEN_7516 : dirty_23_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8073 = _T_12 ? _GEN_7517 : dirty_24_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8074 = _T_12 ? _GEN_7518 : dirty_24_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8075 = _T_12 ? _GEN_7519 : dirty_25_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8076 = _T_12 ? _GEN_7520 : dirty_25_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8077 = _T_12 ? _GEN_7521 : dirty_26_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8078 = _T_12 ? _GEN_7522 : dirty_26_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8079 = _T_12 ? _GEN_7523 : dirty_27_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8080 = _T_12 ? _GEN_7524 : dirty_27_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8081 = _T_12 ? _GEN_7525 : dirty_28_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8082 = _T_12 ? _GEN_7526 : dirty_28_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8083 = _T_12 ? _GEN_7527 : dirty_29_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8084 = _T_12 ? _GEN_7528 : dirty_29_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8085 = _T_12 ? _GEN_7529 : dirty_30_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8086 = _T_12 ? _GEN_7530 : dirty_30_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8087 = _T_12 ? _GEN_7531 : dirty_31_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8088 = _T_12 ? _GEN_7532 : dirty_31_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8089 = _T_12 ? _GEN_7533 : dirty_32_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8090 = _T_12 ? _GEN_7534 : dirty_32_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8091 = _T_12 ? _GEN_7535 : dirty_33_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8092 = _T_12 ? _GEN_7536 : dirty_33_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8093 = _T_12 ? _GEN_7537 : dirty_34_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8094 = _T_12 ? _GEN_7538 : dirty_34_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8095 = _T_12 ? _GEN_7539 : dirty_35_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8096 = _T_12 ? _GEN_7540 : dirty_35_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8097 = _T_12 ? _GEN_7541 : dirty_36_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8098 = _T_12 ? _GEN_7542 : dirty_36_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8099 = _T_12 ? _GEN_7543 : dirty_37_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8100 = _T_12 ? _GEN_7544 : dirty_37_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8101 = _T_12 ? _GEN_7545 : dirty_38_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8102 = _T_12 ? _GEN_7546 : dirty_38_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8103 = _T_12 ? _GEN_7547 : dirty_39_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8104 = _T_12 ? _GEN_7548 : dirty_39_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8105 = _T_12 ? _GEN_7549 : dirty_40_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8106 = _T_12 ? _GEN_7550 : dirty_40_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8107 = _T_12 ? _GEN_7551 : dirty_41_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8108 = _T_12 ? _GEN_7552 : dirty_41_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8109 = _T_12 ? _GEN_7553 : dirty_42_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8110 = _T_12 ? _GEN_7554 : dirty_42_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8111 = _T_12 ? _GEN_7555 : dirty_43_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8112 = _T_12 ? _GEN_7556 : dirty_43_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8113 = _T_12 ? _GEN_7557 : dirty_44_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8114 = _T_12 ? _GEN_7558 : dirty_44_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8115 = _T_12 ? _GEN_7559 : dirty_45_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8116 = _T_12 ? _GEN_7560 : dirty_45_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8117 = _T_12 ? _GEN_7561 : dirty_46_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8118 = _T_12 ? _GEN_7562 : dirty_46_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8119 = _T_12 ? _GEN_7563 : dirty_47_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8120 = _T_12 ? _GEN_7564 : dirty_47_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8121 = _T_12 ? _GEN_7565 : dirty_48_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8122 = _T_12 ? _GEN_7566 : dirty_48_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8123 = _T_12 ? _GEN_7567 : dirty_49_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8124 = _T_12 ? _GEN_7568 : dirty_49_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8125 = _T_12 ? _GEN_7569 : dirty_50_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8126 = _T_12 ? _GEN_7570 : dirty_50_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8127 = _T_12 ? _GEN_7571 : dirty_51_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8128 = _T_12 ? _GEN_7572 : dirty_51_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8129 = _T_12 ? _GEN_7573 : dirty_52_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8130 = _T_12 ? _GEN_7574 : dirty_52_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8131 = _T_12 ? _GEN_7575 : dirty_53_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8132 = _T_12 ? _GEN_7576 : dirty_53_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8133 = _T_12 ? _GEN_7577 : dirty_54_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8134 = _T_12 ? _GEN_7578 : dirty_54_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8135 = _T_12 ? _GEN_7579 : dirty_55_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8136 = _T_12 ? _GEN_7580 : dirty_55_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8137 = _T_12 ? _GEN_7581 : dirty_56_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8138 = _T_12 ? _GEN_7582 : dirty_56_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8139 = _T_12 ? _GEN_7583 : dirty_57_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8140 = _T_12 ? _GEN_7584 : dirty_57_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8141 = _T_12 ? _GEN_7585 : dirty_58_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8142 = _T_12 ? _GEN_7586 : dirty_58_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8143 = _T_12 ? _GEN_7587 : dirty_59_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8144 = _T_12 ? _GEN_7588 : dirty_59_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8145 = _T_12 ? _GEN_7589 : dirty_60_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8146 = _T_12 ? _GEN_7590 : dirty_60_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8147 = _T_12 ? _GEN_7591 : dirty_61_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8148 = _T_12 ? _GEN_7592 : dirty_61_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8149 = _T_12 ? _GEN_7593 : dirty_62_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8150 = _T_12 ? _GEN_7594 : dirty_62_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8151 = _T_12 ? _GEN_7595 : dirty_63_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8152 = _T_12 ? _GEN_7596 : dirty_63_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8153 = _T_12 ? _GEN_7597 : dirty_64_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8154 = _T_12 ? _GEN_7598 : dirty_64_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8155 = _T_12 ? _GEN_7599 : dirty_65_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8156 = _T_12 ? _GEN_7600 : dirty_65_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8157 = _T_12 ? _GEN_7601 : dirty_66_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8158 = _T_12 ? _GEN_7602 : dirty_66_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8159 = _T_12 ? _GEN_7603 : dirty_67_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8160 = _T_12 ? _GEN_7604 : dirty_67_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8161 = _T_12 ? _GEN_7605 : dirty_68_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8162 = _T_12 ? _GEN_7606 : dirty_68_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8163 = _T_12 ? _GEN_7607 : dirty_69_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8164 = _T_12 ? _GEN_7608 : dirty_69_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8165 = _T_12 ? _GEN_7609 : dirty_70_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8166 = _T_12 ? _GEN_7610 : dirty_70_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8167 = _T_12 ? _GEN_7611 : dirty_71_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8168 = _T_12 ? _GEN_7612 : dirty_71_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8169 = _T_12 ? _GEN_7613 : dirty_72_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8170 = _T_12 ? _GEN_7614 : dirty_72_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8171 = _T_12 ? _GEN_7615 : dirty_73_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8172 = _T_12 ? _GEN_7616 : dirty_73_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8173 = _T_12 ? _GEN_7617 : dirty_74_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8174 = _T_12 ? _GEN_7618 : dirty_74_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8175 = _T_12 ? _GEN_7619 : dirty_75_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8176 = _T_12 ? _GEN_7620 : dirty_75_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8177 = _T_12 ? _GEN_7621 : dirty_76_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8178 = _T_12 ? _GEN_7622 : dirty_76_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8179 = _T_12 ? _GEN_7623 : dirty_77_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8180 = _T_12 ? _GEN_7624 : dirty_77_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8181 = _T_12 ? _GEN_7625 : dirty_78_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8182 = _T_12 ? _GEN_7626 : dirty_78_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8183 = _T_12 ? _GEN_7627 : dirty_79_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8184 = _T_12 ? _GEN_7628 : dirty_79_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8185 = _T_12 ? _GEN_7629 : dirty_80_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8186 = _T_12 ? _GEN_7630 : dirty_80_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8187 = _T_12 ? _GEN_7631 : dirty_81_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8188 = _T_12 ? _GEN_7632 : dirty_81_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8189 = _T_12 ? _GEN_7633 : dirty_82_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8190 = _T_12 ? _GEN_7634 : dirty_82_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8191 = _T_12 ? _GEN_7635 : dirty_83_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8192 = _T_12 ? _GEN_7636 : dirty_83_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8193 = _T_12 ? _GEN_7637 : dirty_84_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8194 = _T_12 ? _GEN_7638 : dirty_84_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8195 = _T_12 ? _GEN_7639 : dirty_85_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8196 = _T_12 ? _GEN_7640 : dirty_85_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8197 = _T_12 ? _GEN_7641 : dirty_86_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8198 = _T_12 ? _GEN_7642 : dirty_86_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8199 = _T_12 ? _GEN_7643 : dirty_87_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8200 = _T_12 ? _GEN_7644 : dirty_87_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8201 = _T_12 ? _GEN_7645 : dirty_88_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8202 = _T_12 ? _GEN_7646 : dirty_88_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8203 = _T_12 ? _GEN_7647 : dirty_89_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8204 = _T_12 ? _GEN_7648 : dirty_89_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8205 = _T_12 ? _GEN_7649 : dirty_90_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8206 = _T_12 ? _GEN_7650 : dirty_90_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8207 = _T_12 ? _GEN_7651 : dirty_91_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8208 = _T_12 ? _GEN_7652 : dirty_91_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8209 = _T_12 ? _GEN_7653 : dirty_92_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8210 = _T_12 ? _GEN_7654 : dirty_92_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8211 = _T_12 ? _GEN_7655 : dirty_93_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8212 = _T_12 ? _GEN_7656 : dirty_93_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8213 = _T_12 ? _GEN_7657 : dirty_94_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8214 = _T_12 ? _GEN_7658 : dirty_94_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8215 = _T_12 ? _GEN_7659 : dirty_95_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8216 = _T_12 ? _GEN_7660 : dirty_95_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8217 = _T_12 ? _GEN_7661 : dirty_96_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8218 = _T_12 ? _GEN_7662 : dirty_96_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8219 = _T_12 ? _GEN_7663 : dirty_97_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8220 = _T_12 ? _GEN_7664 : dirty_97_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8221 = _T_12 ? _GEN_7665 : dirty_98_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8222 = _T_12 ? _GEN_7666 : dirty_98_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8223 = _T_12 ? _GEN_7667 : dirty_99_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8224 = _T_12 ? _GEN_7668 : dirty_99_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8225 = _T_12 ? _GEN_7669 : dirty_100_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8226 = _T_12 ? _GEN_7670 : dirty_100_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8227 = _T_12 ? _GEN_7671 : dirty_101_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8228 = _T_12 ? _GEN_7672 : dirty_101_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8229 = _T_12 ? _GEN_7673 : dirty_102_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8230 = _T_12 ? _GEN_7674 : dirty_102_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8231 = _T_12 ? _GEN_7675 : dirty_103_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8232 = _T_12 ? _GEN_7676 : dirty_103_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8233 = _T_12 ? _GEN_7677 : dirty_104_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8234 = _T_12 ? _GEN_7678 : dirty_104_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8235 = _T_12 ? _GEN_7679 : dirty_105_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8236 = _T_12 ? _GEN_7680 : dirty_105_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8237 = _T_12 ? _GEN_7681 : dirty_106_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8238 = _T_12 ? _GEN_7682 : dirty_106_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8239 = _T_12 ? _GEN_7683 : dirty_107_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8240 = _T_12 ? _GEN_7684 : dirty_107_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8241 = _T_12 ? _GEN_7685 : dirty_108_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8242 = _T_12 ? _GEN_7686 : dirty_108_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8243 = _T_12 ? _GEN_7687 : dirty_109_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8244 = _T_12 ? _GEN_7688 : dirty_109_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8245 = _T_12 ? _GEN_7689 : dirty_110_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8246 = _T_12 ? _GEN_7690 : dirty_110_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8247 = _T_12 ? _GEN_7691 : dirty_111_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8248 = _T_12 ? _GEN_7692 : dirty_111_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8249 = _T_12 ? _GEN_7693 : dirty_112_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8250 = _T_12 ? _GEN_7694 : dirty_112_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8251 = _T_12 ? _GEN_7695 : dirty_113_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8252 = _T_12 ? _GEN_7696 : dirty_113_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8253 = _T_12 ? _GEN_7697 : dirty_114_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8254 = _T_12 ? _GEN_7698 : dirty_114_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8255 = _T_12 ? _GEN_7699 : dirty_115_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8256 = _T_12 ? _GEN_7700 : dirty_115_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8257 = _T_12 ? _GEN_7701 : dirty_116_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8258 = _T_12 ? _GEN_7702 : dirty_116_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8259 = _T_12 ? _GEN_7703 : dirty_117_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8260 = _T_12 ? _GEN_7704 : dirty_117_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8261 = _T_12 ? _GEN_7705 : dirty_118_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8262 = _T_12 ? _GEN_7706 : dirty_118_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8263 = _T_12 ? _GEN_7707 : dirty_119_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8264 = _T_12 ? _GEN_7708 : dirty_119_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8265 = _T_12 ? _GEN_7709 : dirty_120_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8266 = _T_12 ? _GEN_7710 : dirty_120_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8267 = _T_12 ? _GEN_7711 : dirty_121_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8268 = _T_12 ? _GEN_7712 : dirty_121_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8269 = _T_12 ? _GEN_7713 : dirty_122_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8270 = _T_12 ? _GEN_7714 : dirty_122_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8271 = _T_12 ? _GEN_7715 : dirty_123_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8272 = _T_12 ? _GEN_7716 : dirty_123_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8273 = _T_12 ? _GEN_7717 : dirty_124_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8274 = _T_12 ? _GEN_7718 : dirty_124_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8275 = _T_12 ? _GEN_7719 : dirty_125_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8276 = _T_12 ? _GEN_7720 : dirty_125_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8277 = _T_12 ? _GEN_7721 : dirty_126_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8278 = _T_12 ? _GEN_7722 : dirty_126_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8279 = _T_12 ? _GEN_7723 : dirty_127_0; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8280 = _T_12 ? _GEN_7724 : dirty_127_1; // @[DCache.scala 418:67 69:22]
  wire  _GEN_8281 = _T_12 ? _GEN_7725 : replace_writeback; // @[DCache.scala 101:40 418:67]
  wire [31:0] _GEN_8282 = _T_12 ? _GEN_7726 : ar_addr; // @[DCache.scala 199:24 418:67]
  wire [7:0] _GEN_8283 = _T_12 ? _GEN_7727 : ar_len; // @[DCache.scala 199:24 418:67]
  wire [2:0] _GEN_8284 = _T_12 ? _GEN_7728 : ar_size; // @[DCache.scala 199:24 418:67]
  wire  _GEN_8285 = _T_12 ? _GEN_7729 : arvalid; // @[DCache.scala 200:24 418:67]
  wire  _GEN_8286 = _T_12 ? _GEN_7730 : rready; // @[DCache.scala 203:23 418:67]
  wire  _GEN_8287 = _T_12 ? _GEN_7731 : ar_handshake; // @[DCache.scala 418:67 99:40]
  wire [3:0] _GEN_8288 = _T_12 ? _GEN_7732 : bram_replace_wea_0; // @[DCache.scala 418:67 73:33]
  wire [3:0] _GEN_8289 = _T_12 ? _GEN_7733 : bram_replace_wea_1; // @[DCache.scala 418:67 73:33]
  wire  _GEN_8290 = _T_12 ? _GEN_7734 : tag_wstrb_0; // @[DCache.scala 418:67 72:33]
  wire  _GEN_8291 = _T_12 ? _GEN_7735 : tag_wstrb_1; // @[DCache.scala 418:67 72:33]
  wire [19:0] _GEN_8292 = _T_12 ? _GEN_7736 : tag_wdata; // @[DCache.scala 418:67 77:26]
  wire [9:0] _GEN_8293 = _T_12 ? _GEN_7737 : bram_replace_write_addr; // @[DCache.scala 418:67 92:40]
  wire  _GEN_8294 = _T_12 ? _GEN_7738 : bram_use_replace_addr; // @[DCache.scala 418:67 95:40]
  wire  _GEN_8295 = _T_12 ? _GEN_7739 : valid_0_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8296 = _T_12 ? _GEN_7740 : valid_0_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8297 = _T_12 ? _GEN_7741 : valid_1_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8298 = _T_12 ? _GEN_7742 : valid_1_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8299 = _T_12 ? _GEN_7743 : valid_2_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8300 = _T_12 ? _GEN_7744 : valid_2_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8301 = _T_12 ? _GEN_7745 : valid_3_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8302 = _T_12 ? _GEN_7746 : valid_3_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8303 = _T_12 ? _GEN_7747 : valid_4_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8304 = _T_12 ? _GEN_7748 : valid_4_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8305 = _T_12 ? _GEN_7749 : valid_5_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8306 = _T_12 ? _GEN_7750 : valid_5_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8307 = _T_12 ? _GEN_7751 : valid_6_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8308 = _T_12 ? _GEN_7752 : valid_6_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8309 = _T_12 ? _GEN_7753 : valid_7_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8310 = _T_12 ? _GEN_7754 : valid_7_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8311 = _T_12 ? _GEN_7755 : valid_8_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8312 = _T_12 ? _GEN_7756 : valid_8_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8313 = _T_12 ? _GEN_7757 : valid_9_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8314 = _T_12 ? _GEN_7758 : valid_9_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8315 = _T_12 ? _GEN_7759 : valid_10_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8316 = _T_12 ? _GEN_7760 : valid_10_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8317 = _T_12 ? _GEN_7761 : valid_11_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8318 = _T_12 ? _GEN_7762 : valid_11_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8319 = _T_12 ? _GEN_7763 : valid_12_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8320 = _T_12 ? _GEN_7764 : valid_12_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8321 = _T_12 ? _GEN_7765 : valid_13_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8322 = _T_12 ? _GEN_7766 : valid_13_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8323 = _T_12 ? _GEN_7767 : valid_14_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8324 = _T_12 ? _GEN_7768 : valid_14_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8325 = _T_12 ? _GEN_7769 : valid_15_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8326 = _T_12 ? _GEN_7770 : valid_15_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8327 = _T_12 ? _GEN_7771 : valid_16_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8328 = _T_12 ? _GEN_7772 : valid_16_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8329 = _T_12 ? _GEN_7773 : valid_17_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8330 = _T_12 ? _GEN_7774 : valid_17_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8331 = _T_12 ? _GEN_7775 : valid_18_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8332 = _T_12 ? _GEN_7776 : valid_18_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8333 = _T_12 ? _GEN_7777 : valid_19_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8334 = _T_12 ? _GEN_7778 : valid_19_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8335 = _T_12 ? _GEN_7779 : valid_20_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8336 = _T_12 ? _GEN_7780 : valid_20_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8337 = _T_12 ? _GEN_7781 : valid_21_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8338 = _T_12 ? _GEN_7782 : valid_21_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8339 = _T_12 ? _GEN_7783 : valid_22_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8340 = _T_12 ? _GEN_7784 : valid_22_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8341 = _T_12 ? _GEN_7785 : valid_23_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8342 = _T_12 ? _GEN_7786 : valid_23_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8343 = _T_12 ? _GEN_7787 : valid_24_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8344 = _T_12 ? _GEN_7788 : valid_24_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8345 = _T_12 ? _GEN_7789 : valid_25_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8346 = _T_12 ? _GEN_7790 : valid_25_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8347 = _T_12 ? _GEN_7791 : valid_26_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8348 = _T_12 ? _GEN_7792 : valid_26_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8349 = _T_12 ? _GEN_7793 : valid_27_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8350 = _T_12 ? _GEN_7794 : valid_27_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8351 = _T_12 ? _GEN_7795 : valid_28_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8352 = _T_12 ? _GEN_7796 : valid_28_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8353 = _T_12 ? _GEN_7797 : valid_29_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8354 = _T_12 ? _GEN_7798 : valid_29_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8355 = _T_12 ? _GEN_7799 : valid_30_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8356 = _T_12 ? _GEN_7800 : valid_30_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8357 = _T_12 ? _GEN_7801 : valid_31_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8358 = _T_12 ? _GEN_7802 : valid_31_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8359 = _T_12 ? _GEN_7803 : valid_32_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8360 = _T_12 ? _GEN_7804 : valid_32_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8361 = _T_12 ? _GEN_7805 : valid_33_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8362 = _T_12 ? _GEN_7806 : valid_33_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8363 = _T_12 ? _GEN_7807 : valid_34_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8364 = _T_12 ? _GEN_7808 : valid_34_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8365 = _T_12 ? _GEN_7809 : valid_35_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8366 = _T_12 ? _GEN_7810 : valid_35_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8367 = _T_12 ? _GEN_7811 : valid_36_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8368 = _T_12 ? _GEN_7812 : valid_36_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8369 = _T_12 ? _GEN_7813 : valid_37_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8370 = _T_12 ? _GEN_7814 : valid_37_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8371 = _T_12 ? _GEN_7815 : valid_38_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8372 = _T_12 ? _GEN_7816 : valid_38_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8373 = _T_12 ? _GEN_7817 : valid_39_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8374 = _T_12 ? _GEN_7818 : valid_39_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8375 = _T_12 ? _GEN_7819 : valid_40_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8376 = _T_12 ? _GEN_7820 : valid_40_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8377 = _T_12 ? _GEN_7821 : valid_41_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8378 = _T_12 ? _GEN_7822 : valid_41_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8379 = _T_12 ? _GEN_7823 : valid_42_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8380 = _T_12 ? _GEN_7824 : valid_42_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8381 = _T_12 ? _GEN_7825 : valid_43_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8382 = _T_12 ? _GEN_7826 : valid_43_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8383 = _T_12 ? _GEN_7827 : valid_44_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8384 = _T_12 ? _GEN_7828 : valid_44_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8385 = _T_12 ? _GEN_7829 : valid_45_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8386 = _T_12 ? _GEN_7830 : valid_45_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8387 = _T_12 ? _GEN_7831 : valid_46_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8388 = _T_12 ? _GEN_7832 : valid_46_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8389 = _T_12 ? _GEN_7833 : valid_47_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8390 = _T_12 ? _GEN_7834 : valid_47_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8391 = _T_12 ? _GEN_7835 : valid_48_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8392 = _T_12 ? _GEN_7836 : valid_48_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8393 = _T_12 ? _GEN_7837 : valid_49_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8394 = _T_12 ? _GEN_7838 : valid_49_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8395 = _T_12 ? _GEN_7839 : valid_50_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8396 = _T_12 ? _GEN_7840 : valid_50_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8397 = _T_12 ? _GEN_7841 : valid_51_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8398 = _T_12 ? _GEN_7842 : valid_51_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8399 = _T_12 ? _GEN_7843 : valid_52_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8400 = _T_12 ? _GEN_7844 : valid_52_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8401 = _T_12 ? _GEN_7845 : valid_53_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8402 = _T_12 ? _GEN_7846 : valid_53_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8403 = _T_12 ? _GEN_7847 : valid_54_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8404 = _T_12 ? _GEN_7848 : valid_54_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8405 = _T_12 ? _GEN_7849 : valid_55_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8406 = _T_12 ? _GEN_7850 : valid_55_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8407 = _T_12 ? _GEN_7851 : valid_56_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8408 = _T_12 ? _GEN_7852 : valid_56_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8409 = _T_12 ? _GEN_7853 : valid_57_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8410 = _T_12 ? _GEN_7854 : valid_57_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8411 = _T_12 ? _GEN_7855 : valid_58_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8412 = _T_12 ? _GEN_7856 : valid_58_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8413 = _T_12 ? _GEN_7857 : valid_59_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8414 = _T_12 ? _GEN_7858 : valid_59_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8415 = _T_12 ? _GEN_7859 : valid_60_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8416 = _T_12 ? _GEN_7860 : valid_60_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8417 = _T_12 ? _GEN_7861 : valid_61_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8418 = _T_12 ? _GEN_7862 : valid_61_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8419 = _T_12 ? _GEN_7863 : valid_62_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8420 = _T_12 ? _GEN_7864 : valid_62_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8421 = _T_12 ? _GEN_7865 : valid_63_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8422 = _T_12 ? _GEN_7866 : valid_63_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8423 = _T_12 ? _GEN_7867 : valid_64_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8424 = _T_12 ? _GEN_7868 : valid_64_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8425 = _T_12 ? _GEN_7869 : valid_65_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8426 = _T_12 ? _GEN_7870 : valid_65_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8427 = _T_12 ? _GEN_7871 : valid_66_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8428 = _T_12 ? _GEN_7872 : valid_66_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8429 = _T_12 ? _GEN_7873 : valid_67_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8430 = _T_12 ? _GEN_7874 : valid_67_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8431 = _T_12 ? _GEN_7875 : valid_68_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8432 = _T_12 ? _GEN_7876 : valid_68_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8433 = _T_12 ? _GEN_7877 : valid_69_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8434 = _T_12 ? _GEN_7878 : valid_69_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8435 = _T_12 ? _GEN_7879 : valid_70_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8436 = _T_12 ? _GEN_7880 : valid_70_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8437 = _T_12 ? _GEN_7881 : valid_71_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8438 = _T_12 ? _GEN_7882 : valid_71_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8439 = _T_12 ? _GEN_7883 : valid_72_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8440 = _T_12 ? _GEN_7884 : valid_72_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8441 = _T_12 ? _GEN_7885 : valid_73_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8442 = _T_12 ? _GEN_7886 : valid_73_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8443 = _T_12 ? _GEN_7887 : valid_74_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8444 = _T_12 ? _GEN_7888 : valid_74_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8445 = _T_12 ? _GEN_7889 : valid_75_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8446 = _T_12 ? _GEN_7890 : valid_75_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8447 = _T_12 ? _GEN_7891 : valid_76_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8448 = _T_12 ? _GEN_7892 : valid_76_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8449 = _T_12 ? _GEN_7893 : valid_77_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8450 = _T_12 ? _GEN_7894 : valid_77_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8451 = _T_12 ? _GEN_7895 : valid_78_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8452 = _T_12 ? _GEN_7896 : valid_78_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8453 = _T_12 ? _GEN_7897 : valid_79_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8454 = _T_12 ? _GEN_7898 : valid_79_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8455 = _T_12 ? _GEN_7899 : valid_80_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8456 = _T_12 ? _GEN_7900 : valid_80_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8457 = _T_12 ? _GEN_7901 : valid_81_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8458 = _T_12 ? _GEN_7902 : valid_81_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8459 = _T_12 ? _GEN_7903 : valid_82_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8460 = _T_12 ? _GEN_7904 : valid_82_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8461 = _T_12 ? _GEN_7905 : valid_83_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8462 = _T_12 ? _GEN_7906 : valid_83_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8463 = _T_12 ? _GEN_7907 : valid_84_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8464 = _T_12 ? _GEN_7908 : valid_84_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8465 = _T_12 ? _GEN_7909 : valid_85_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8466 = _T_12 ? _GEN_7910 : valid_85_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8467 = _T_12 ? _GEN_7911 : valid_86_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8468 = _T_12 ? _GEN_7912 : valid_86_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8469 = _T_12 ? _GEN_7913 : valid_87_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8470 = _T_12 ? _GEN_7914 : valid_87_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8471 = _T_12 ? _GEN_7915 : valid_88_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8472 = _T_12 ? _GEN_7916 : valid_88_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8473 = _T_12 ? _GEN_7917 : valid_89_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8474 = _T_12 ? _GEN_7918 : valid_89_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8475 = _T_12 ? _GEN_7919 : valid_90_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8476 = _T_12 ? _GEN_7920 : valid_90_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8477 = _T_12 ? _GEN_7921 : valid_91_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8478 = _T_12 ? _GEN_7922 : valid_91_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8479 = _T_12 ? _GEN_7923 : valid_92_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8480 = _T_12 ? _GEN_7924 : valid_92_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8481 = _T_12 ? _GEN_7925 : valid_93_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8482 = _T_12 ? _GEN_7926 : valid_93_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8483 = _T_12 ? _GEN_7927 : valid_94_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8484 = _T_12 ? _GEN_7928 : valid_94_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8485 = _T_12 ? _GEN_7929 : valid_95_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8486 = _T_12 ? _GEN_7930 : valid_95_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8487 = _T_12 ? _GEN_7931 : valid_96_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8488 = _T_12 ? _GEN_7932 : valid_96_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8489 = _T_12 ? _GEN_7933 : valid_97_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8490 = _T_12 ? _GEN_7934 : valid_97_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8491 = _T_12 ? _GEN_7935 : valid_98_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8492 = _T_12 ? _GEN_7936 : valid_98_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8493 = _T_12 ? _GEN_7937 : valid_99_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8494 = _T_12 ? _GEN_7938 : valid_99_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8495 = _T_12 ? _GEN_7939 : valid_100_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8496 = _T_12 ? _GEN_7940 : valid_100_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8497 = _T_12 ? _GEN_7941 : valid_101_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8498 = _T_12 ? _GEN_7942 : valid_101_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8499 = _T_12 ? _GEN_7943 : valid_102_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8500 = _T_12 ? _GEN_7944 : valid_102_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8501 = _T_12 ? _GEN_7945 : valid_103_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8502 = _T_12 ? _GEN_7946 : valid_103_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8503 = _T_12 ? _GEN_7947 : valid_104_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8504 = _T_12 ? _GEN_7948 : valid_104_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8505 = _T_12 ? _GEN_7949 : valid_105_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8506 = _T_12 ? _GEN_7950 : valid_105_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8507 = _T_12 ? _GEN_7951 : valid_106_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8508 = _T_12 ? _GEN_7952 : valid_106_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8509 = _T_12 ? _GEN_7953 : valid_107_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8510 = _T_12 ? _GEN_7954 : valid_107_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8511 = _T_12 ? _GEN_7955 : valid_108_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8512 = _T_12 ? _GEN_7956 : valid_108_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8513 = _T_12 ? _GEN_7957 : valid_109_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8514 = _T_12 ? _GEN_7958 : valid_109_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8515 = _T_12 ? _GEN_7959 : valid_110_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8516 = _T_12 ? _GEN_7960 : valid_110_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8517 = _T_12 ? _GEN_7961 : valid_111_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8518 = _T_12 ? _GEN_7962 : valid_111_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8519 = _T_12 ? _GEN_7963 : valid_112_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8520 = _T_12 ? _GEN_7964 : valid_112_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8521 = _T_12 ? _GEN_7965 : valid_113_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8522 = _T_12 ? _GEN_7966 : valid_113_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8523 = _T_12 ? _GEN_7967 : valid_114_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8524 = _T_12 ? _GEN_7968 : valid_114_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8525 = _T_12 ? _GEN_7969 : valid_115_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8526 = _T_12 ? _GEN_7970 : valid_115_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8527 = _T_12 ? _GEN_7971 : valid_116_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8528 = _T_12 ? _GEN_7972 : valid_116_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8529 = _T_12 ? _GEN_7973 : valid_117_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8530 = _T_12 ? _GEN_7974 : valid_117_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8531 = _T_12 ? _GEN_7975 : valid_118_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8532 = _T_12 ? _GEN_7976 : valid_118_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8533 = _T_12 ? _GEN_7977 : valid_119_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8534 = _T_12 ? _GEN_7978 : valid_119_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8535 = _T_12 ? _GEN_7979 : valid_120_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8536 = _T_12 ? _GEN_7980 : valid_120_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8537 = _T_12 ? _GEN_7981 : valid_121_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8538 = _T_12 ? _GEN_7982 : valid_121_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8539 = _T_12 ? _GEN_7983 : valid_122_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8540 = _T_12 ? _GEN_7984 : valid_122_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8541 = _T_12 ? _GEN_7985 : valid_123_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8542 = _T_12 ? _GEN_7986 : valid_123_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8543 = _T_12 ? _GEN_7987 : valid_124_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8544 = _T_12 ? _GEN_7988 : valid_124_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8545 = _T_12 ? _GEN_7989 : valid_125_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8546 = _T_12 ? _GEN_7990 : valid_125_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8547 = _T_12 ? _GEN_7991 : valid_126_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8548 = _T_12 ? _GEN_7992 : valid_126_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8549 = _T_12 ? _GEN_7993 : valid_127_0; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8550 = _T_12 ? _GEN_7994 : valid_127_1; // @[DCache.scala 418:67 68:22]
  wire  _GEN_8551 = _T_12 ? _GEN_7995 : replace_working; // @[DCache.scala 418:67 98:40]
  wire [2:0] _GEN_8552 = _T_12 ? _GEN_7996 : state; // @[DCache.scala 418:67 65:96]
  wire [2:0] _GEN_8553 = _T_10 ? 3'h0 : state; // @[DCache.scala 504:39 505:26 65:96]
  wire  _GEN_8554 = _T_10 ? 1'h0 : data_tlb_invalid; // @[DCache.scala 250:25 504:39 506:26]
  wire  _GEN_8555 = _T_10 ? 1'h0 : data_tlb_refill; // @[DCache.scala 250:25 504:39 507:26]
  wire  _GEN_8556 = _T_10 ? 1'h0 : data_tlb_mod; // @[DCache.scala 250:25 504:39 508:26]
  wire [2:0] _GEN_8557 = 3'h5 == state ? _GEN_8553 : state; // @[DCache.scala 260:17 65:96]
  wire  _GEN_8558 = 3'h5 == state ? _GEN_8554 : data_tlb_invalid; // @[DCache.scala 260:17 250:25]
  wire  _GEN_8559 = 3'h5 == state ? _GEN_8555 : data_tlb_refill; // @[DCache.scala 260:17 250:25]
  wire  _GEN_8560 = 3'h5 == state ? _GEN_8556 : data_tlb_mod; // @[DCache.scala 260:17 250:25]
  wire [9:0] _GEN_8561 = 3'h4 == state ? _GEN_7997 : bram_replace_addr; // @[DCache.scala 260:17 90:40]
  wire [9:0] _GEN_8562 = 3'h4 == state ? _GEN_7998 : bram_read_ready_addr; // @[DCache.scala 260:17 91:40]
  wire [31:0] _GEN_8563 = 3'h4 == state ? _GEN_7999 : bram_r_buffer_0; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8564 = 3'h4 == state ? _GEN_8000 : bram_r_buffer_1; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8565 = 3'h4 == state ? _GEN_8001 : bram_r_buffer_2; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8566 = 3'h4 == state ? _GEN_8002 : bram_r_buffer_3; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8567 = 3'h4 == state ? _GEN_8003 : bram_r_buffer_4; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8568 = 3'h4 == state ? _GEN_8004 : bram_r_buffer_5; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8569 = 3'h4 == state ? _GEN_8005 : bram_r_buffer_6; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8570 = 3'h4 == state ? _GEN_8006 : bram_r_buffer_7; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8571 = 3'h4 == state ? _GEN_8007 : bram_r_buffer_8; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8572 = 3'h4 == state ? _GEN_8008 : bram_r_buffer_9; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8573 = 3'h4 == state ? _GEN_8009 : bram_r_buffer_10; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8574 = 3'h4 == state ? _GEN_8010 : bram_r_buffer_11; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8575 = 3'h4 == state ? _GEN_8011 : bram_r_buffer_12; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8576 = 3'h4 == state ? _GEN_8012 : bram_r_buffer_13; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8577 = 3'h4 == state ? _GEN_8013 : bram_r_buffer_14; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8578 = 3'h4 == state ? _GEN_8014 : bram_r_buffer_15; // @[DCache.scala 260:17 94:40]
  wire [31:0] _GEN_8579 = 3'h4 == state ? _GEN_8015 : _GEN_281; // @[DCache.scala 260:17]
  wire [7:0] _GEN_8580 = 3'h4 == state ? _GEN_8016 : _GEN_285; // @[DCache.scala 260:17]
  wire [2:0] _GEN_8581 = 3'h4 == state ? _GEN_8017 : _GEN_282; // @[DCache.scala 260:17]
  wire  _GEN_8582 = 3'h4 == state ? _GEN_8018 : _GEN_276; // @[DCache.scala 260:17]
  wire [31:0] _GEN_8583 = 3'h4 == state ? _GEN_8019 : _GEN_283; // @[DCache.scala 260:17]
  wire [3:0] _GEN_8584 = 3'h4 == state ? _GEN_8020 : _GEN_284; // @[DCache.scala 260:17]
  wire  _GEN_8585 = 3'h4 == state ? _GEN_8021 : _GEN_278; // @[DCache.scala 260:17]
  wire  _GEN_8586 = 3'h4 == state ? _GEN_8022 : _GEN_277; // @[DCache.scala 260:17]
  wire  _GEN_8587 = 3'h4 == state ? _GEN_8023 : aw_handshake; // @[DCache.scala 260:17 100:40]
  wire [3:0] _GEN_8588 = 3'h4 == state ? _GEN_8024 : axi_wcnt; // @[DCache.scala 260:17 89:40]
  wire  _GEN_8589 = 3'h4 == state ? _GEN_8025 : dirty_0_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8590 = 3'h4 == state ? _GEN_8026 : dirty_0_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8591 = 3'h4 == state ? _GEN_8027 : dirty_1_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8592 = 3'h4 == state ? _GEN_8028 : dirty_1_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8593 = 3'h4 == state ? _GEN_8029 : dirty_2_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8594 = 3'h4 == state ? _GEN_8030 : dirty_2_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8595 = 3'h4 == state ? _GEN_8031 : dirty_3_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8596 = 3'h4 == state ? _GEN_8032 : dirty_3_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8597 = 3'h4 == state ? _GEN_8033 : dirty_4_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8598 = 3'h4 == state ? _GEN_8034 : dirty_4_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8599 = 3'h4 == state ? _GEN_8035 : dirty_5_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8600 = 3'h4 == state ? _GEN_8036 : dirty_5_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8601 = 3'h4 == state ? _GEN_8037 : dirty_6_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8602 = 3'h4 == state ? _GEN_8038 : dirty_6_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8603 = 3'h4 == state ? _GEN_8039 : dirty_7_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8604 = 3'h4 == state ? _GEN_8040 : dirty_7_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8605 = 3'h4 == state ? _GEN_8041 : dirty_8_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8606 = 3'h4 == state ? _GEN_8042 : dirty_8_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8607 = 3'h4 == state ? _GEN_8043 : dirty_9_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8608 = 3'h4 == state ? _GEN_8044 : dirty_9_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8609 = 3'h4 == state ? _GEN_8045 : dirty_10_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8610 = 3'h4 == state ? _GEN_8046 : dirty_10_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8611 = 3'h4 == state ? _GEN_8047 : dirty_11_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8612 = 3'h4 == state ? _GEN_8048 : dirty_11_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8613 = 3'h4 == state ? _GEN_8049 : dirty_12_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8614 = 3'h4 == state ? _GEN_8050 : dirty_12_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8615 = 3'h4 == state ? _GEN_8051 : dirty_13_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8616 = 3'h4 == state ? _GEN_8052 : dirty_13_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8617 = 3'h4 == state ? _GEN_8053 : dirty_14_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8618 = 3'h4 == state ? _GEN_8054 : dirty_14_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8619 = 3'h4 == state ? _GEN_8055 : dirty_15_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8620 = 3'h4 == state ? _GEN_8056 : dirty_15_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8621 = 3'h4 == state ? _GEN_8057 : dirty_16_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8622 = 3'h4 == state ? _GEN_8058 : dirty_16_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8623 = 3'h4 == state ? _GEN_8059 : dirty_17_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8624 = 3'h4 == state ? _GEN_8060 : dirty_17_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8625 = 3'h4 == state ? _GEN_8061 : dirty_18_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8626 = 3'h4 == state ? _GEN_8062 : dirty_18_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8627 = 3'h4 == state ? _GEN_8063 : dirty_19_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8628 = 3'h4 == state ? _GEN_8064 : dirty_19_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8629 = 3'h4 == state ? _GEN_8065 : dirty_20_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8630 = 3'h4 == state ? _GEN_8066 : dirty_20_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8631 = 3'h4 == state ? _GEN_8067 : dirty_21_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8632 = 3'h4 == state ? _GEN_8068 : dirty_21_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8633 = 3'h4 == state ? _GEN_8069 : dirty_22_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8634 = 3'h4 == state ? _GEN_8070 : dirty_22_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8635 = 3'h4 == state ? _GEN_8071 : dirty_23_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8636 = 3'h4 == state ? _GEN_8072 : dirty_23_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8637 = 3'h4 == state ? _GEN_8073 : dirty_24_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8638 = 3'h4 == state ? _GEN_8074 : dirty_24_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8639 = 3'h4 == state ? _GEN_8075 : dirty_25_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8640 = 3'h4 == state ? _GEN_8076 : dirty_25_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8641 = 3'h4 == state ? _GEN_8077 : dirty_26_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8642 = 3'h4 == state ? _GEN_8078 : dirty_26_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8643 = 3'h4 == state ? _GEN_8079 : dirty_27_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8644 = 3'h4 == state ? _GEN_8080 : dirty_27_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8645 = 3'h4 == state ? _GEN_8081 : dirty_28_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8646 = 3'h4 == state ? _GEN_8082 : dirty_28_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8647 = 3'h4 == state ? _GEN_8083 : dirty_29_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8648 = 3'h4 == state ? _GEN_8084 : dirty_29_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8649 = 3'h4 == state ? _GEN_8085 : dirty_30_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8650 = 3'h4 == state ? _GEN_8086 : dirty_30_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8651 = 3'h4 == state ? _GEN_8087 : dirty_31_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8652 = 3'h4 == state ? _GEN_8088 : dirty_31_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8653 = 3'h4 == state ? _GEN_8089 : dirty_32_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8654 = 3'h4 == state ? _GEN_8090 : dirty_32_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8655 = 3'h4 == state ? _GEN_8091 : dirty_33_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8656 = 3'h4 == state ? _GEN_8092 : dirty_33_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8657 = 3'h4 == state ? _GEN_8093 : dirty_34_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8658 = 3'h4 == state ? _GEN_8094 : dirty_34_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8659 = 3'h4 == state ? _GEN_8095 : dirty_35_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8660 = 3'h4 == state ? _GEN_8096 : dirty_35_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8661 = 3'h4 == state ? _GEN_8097 : dirty_36_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8662 = 3'h4 == state ? _GEN_8098 : dirty_36_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8663 = 3'h4 == state ? _GEN_8099 : dirty_37_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8664 = 3'h4 == state ? _GEN_8100 : dirty_37_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8665 = 3'h4 == state ? _GEN_8101 : dirty_38_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8666 = 3'h4 == state ? _GEN_8102 : dirty_38_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8667 = 3'h4 == state ? _GEN_8103 : dirty_39_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8668 = 3'h4 == state ? _GEN_8104 : dirty_39_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8669 = 3'h4 == state ? _GEN_8105 : dirty_40_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8670 = 3'h4 == state ? _GEN_8106 : dirty_40_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8671 = 3'h4 == state ? _GEN_8107 : dirty_41_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8672 = 3'h4 == state ? _GEN_8108 : dirty_41_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8673 = 3'h4 == state ? _GEN_8109 : dirty_42_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8674 = 3'h4 == state ? _GEN_8110 : dirty_42_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8675 = 3'h4 == state ? _GEN_8111 : dirty_43_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8676 = 3'h4 == state ? _GEN_8112 : dirty_43_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8677 = 3'h4 == state ? _GEN_8113 : dirty_44_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8678 = 3'h4 == state ? _GEN_8114 : dirty_44_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8679 = 3'h4 == state ? _GEN_8115 : dirty_45_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8680 = 3'h4 == state ? _GEN_8116 : dirty_45_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8681 = 3'h4 == state ? _GEN_8117 : dirty_46_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8682 = 3'h4 == state ? _GEN_8118 : dirty_46_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8683 = 3'h4 == state ? _GEN_8119 : dirty_47_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8684 = 3'h4 == state ? _GEN_8120 : dirty_47_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8685 = 3'h4 == state ? _GEN_8121 : dirty_48_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8686 = 3'h4 == state ? _GEN_8122 : dirty_48_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8687 = 3'h4 == state ? _GEN_8123 : dirty_49_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8688 = 3'h4 == state ? _GEN_8124 : dirty_49_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8689 = 3'h4 == state ? _GEN_8125 : dirty_50_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8690 = 3'h4 == state ? _GEN_8126 : dirty_50_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8691 = 3'h4 == state ? _GEN_8127 : dirty_51_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8692 = 3'h4 == state ? _GEN_8128 : dirty_51_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8693 = 3'h4 == state ? _GEN_8129 : dirty_52_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8694 = 3'h4 == state ? _GEN_8130 : dirty_52_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8695 = 3'h4 == state ? _GEN_8131 : dirty_53_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8696 = 3'h4 == state ? _GEN_8132 : dirty_53_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8697 = 3'h4 == state ? _GEN_8133 : dirty_54_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8698 = 3'h4 == state ? _GEN_8134 : dirty_54_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8699 = 3'h4 == state ? _GEN_8135 : dirty_55_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8700 = 3'h4 == state ? _GEN_8136 : dirty_55_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8701 = 3'h4 == state ? _GEN_8137 : dirty_56_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8702 = 3'h4 == state ? _GEN_8138 : dirty_56_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8703 = 3'h4 == state ? _GEN_8139 : dirty_57_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8704 = 3'h4 == state ? _GEN_8140 : dirty_57_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8705 = 3'h4 == state ? _GEN_8141 : dirty_58_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8706 = 3'h4 == state ? _GEN_8142 : dirty_58_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8707 = 3'h4 == state ? _GEN_8143 : dirty_59_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8708 = 3'h4 == state ? _GEN_8144 : dirty_59_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8709 = 3'h4 == state ? _GEN_8145 : dirty_60_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8710 = 3'h4 == state ? _GEN_8146 : dirty_60_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8711 = 3'h4 == state ? _GEN_8147 : dirty_61_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8712 = 3'h4 == state ? _GEN_8148 : dirty_61_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8713 = 3'h4 == state ? _GEN_8149 : dirty_62_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8714 = 3'h4 == state ? _GEN_8150 : dirty_62_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8715 = 3'h4 == state ? _GEN_8151 : dirty_63_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8716 = 3'h4 == state ? _GEN_8152 : dirty_63_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8717 = 3'h4 == state ? _GEN_8153 : dirty_64_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8718 = 3'h4 == state ? _GEN_8154 : dirty_64_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8719 = 3'h4 == state ? _GEN_8155 : dirty_65_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8720 = 3'h4 == state ? _GEN_8156 : dirty_65_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8721 = 3'h4 == state ? _GEN_8157 : dirty_66_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8722 = 3'h4 == state ? _GEN_8158 : dirty_66_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8723 = 3'h4 == state ? _GEN_8159 : dirty_67_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8724 = 3'h4 == state ? _GEN_8160 : dirty_67_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8725 = 3'h4 == state ? _GEN_8161 : dirty_68_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8726 = 3'h4 == state ? _GEN_8162 : dirty_68_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8727 = 3'h4 == state ? _GEN_8163 : dirty_69_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8728 = 3'h4 == state ? _GEN_8164 : dirty_69_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8729 = 3'h4 == state ? _GEN_8165 : dirty_70_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8730 = 3'h4 == state ? _GEN_8166 : dirty_70_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8731 = 3'h4 == state ? _GEN_8167 : dirty_71_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8732 = 3'h4 == state ? _GEN_8168 : dirty_71_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8733 = 3'h4 == state ? _GEN_8169 : dirty_72_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8734 = 3'h4 == state ? _GEN_8170 : dirty_72_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8735 = 3'h4 == state ? _GEN_8171 : dirty_73_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8736 = 3'h4 == state ? _GEN_8172 : dirty_73_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8737 = 3'h4 == state ? _GEN_8173 : dirty_74_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8738 = 3'h4 == state ? _GEN_8174 : dirty_74_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8739 = 3'h4 == state ? _GEN_8175 : dirty_75_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8740 = 3'h4 == state ? _GEN_8176 : dirty_75_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8741 = 3'h4 == state ? _GEN_8177 : dirty_76_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8742 = 3'h4 == state ? _GEN_8178 : dirty_76_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8743 = 3'h4 == state ? _GEN_8179 : dirty_77_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8744 = 3'h4 == state ? _GEN_8180 : dirty_77_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8745 = 3'h4 == state ? _GEN_8181 : dirty_78_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8746 = 3'h4 == state ? _GEN_8182 : dirty_78_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8747 = 3'h4 == state ? _GEN_8183 : dirty_79_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8748 = 3'h4 == state ? _GEN_8184 : dirty_79_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8749 = 3'h4 == state ? _GEN_8185 : dirty_80_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8750 = 3'h4 == state ? _GEN_8186 : dirty_80_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8751 = 3'h4 == state ? _GEN_8187 : dirty_81_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8752 = 3'h4 == state ? _GEN_8188 : dirty_81_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8753 = 3'h4 == state ? _GEN_8189 : dirty_82_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8754 = 3'h4 == state ? _GEN_8190 : dirty_82_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8755 = 3'h4 == state ? _GEN_8191 : dirty_83_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8756 = 3'h4 == state ? _GEN_8192 : dirty_83_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8757 = 3'h4 == state ? _GEN_8193 : dirty_84_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8758 = 3'h4 == state ? _GEN_8194 : dirty_84_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8759 = 3'h4 == state ? _GEN_8195 : dirty_85_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8760 = 3'h4 == state ? _GEN_8196 : dirty_85_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8761 = 3'h4 == state ? _GEN_8197 : dirty_86_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8762 = 3'h4 == state ? _GEN_8198 : dirty_86_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8763 = 3'h4 == state ? _GEN_8199 : dirty_87_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8764 = 3'h4 == state ? _GEN_8200 : dirty_87_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8765 = 3'h4 == state ? _GEN_8201 : dirty_88_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8766 = 3'h4 == state ? _GEN_8202 : dirty_88_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8767 = 3'h4 == state ? _GEN_8203 : dirty_89_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8768 = 3'h4 == state ? _GEN_8204 : dirty_89_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8769 = 3'h4 == state ? _GEN_8205 : dirty_90_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8770 = 3'h4 == state ? _GEN_8206 : dirty_90_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8771 = 3'h4 == state ? _GEN_8207 : dirty_91_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8772 = 3'h4 == state ? _GEN_8208 : dirty_91_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8773 = 3'h4 == state ? _GEN_8209 : dirty_92_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8774 = 3'h4 == state ? _GEN_8210 : dirty_92_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8775 = 3'h4 == state ? _GEN_8211 : dirty_93_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8776 = 3'h4 == state ? _GEN_8212 : dirty_93_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8777 = 3'h4 == state ? _GEN_8213 : dirty_94_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8778 = 3'h4 == state ? _GEN_8214 : dirty_94_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8779 = 3'h4 == state ? _GEN_8215 : dirty_95_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8780 = 3'h4 == state ? _GEN_8216 : dirty_95_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8781 = 3'h4 == state ? _GEN_8217 : dirty_96_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8782 = 3'h4 == state ? _GEN_8218 : dirty_96_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8783 = 3'h4 == state ? _GEN_8219 : dirty_97_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8784 = 3'h4 == state ? _GEN_8220 : dirty_97_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8785 = 3'h4 == state ? _GEN_8221 : dirty_98_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8786 = 3'h4 == state ? _GEN_8222 : dirty_98_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8787 = 3'h4 == state ? _GEN_8223 : dirty_99_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8788 = 3'h4 == state ? _GEN_8224 : dirty_99_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8789 = 3'h4 == state ? _GEN_8225 : dirty_100_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8790 = 3'h4 == state ? _GEN_8226 : dirty_100_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8791 = 3'h4 == state ? _GEN_8227 : dirty_101_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8792 = 3'h4 == state ? _GEN_8228 : dirty_101_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8793 = 3'h4 == state ? _GEN_8229 : dirty_102_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8794 = 3'h4 == state ? _GEN_8230 : dirty_102_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8795 = 3'h4 == state ? _GEN_8231 : dirty_103_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8796 = 3'h4 == state ? _GEN_8232 : dirty_103_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8797 = 3'h4 == state ? _GEN_8233 : dirty_104_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8798 = 3'h4 == state ? _GEN_8234 : dirty_104_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8799 = 3'h4 == state ? _GEN_8235 : dirty_105_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8800 = 3'h4 == state ? _GEN_8236 : dirty_105_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8801 = 3'h4 == state ? _GEN_8237 : dirty_106_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8802 = 3'h4 == state ? _GEN_8238 : dirty_106_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8803 = 3'h4 == state ? _GEN_8239 : dirty_107_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8804 = 3'h4 == state ? _GEN_8240 : dirty_107_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8805 = 3'h4 == state ? _GEN_8241 : dirty_108_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8806 = 3'h4 == state ? _GEN_8242 : dirty_108_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8807 = 3'h4 == state ? _GEN_8243 : dirty_109_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8808 = 3'h4 == state ? _GEN_8244 : dirty_109_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8809 = 3'h4 == state ? _GEN_8245 : dirty_110_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8810 = 3'h4 == state ? _GEN_8246 : dirty_110_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8811 = 3'h4 == state ? _GEN_8247 : dirty_111_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8812 = 3'h4 == state ? _GEN_8248 : dirty_111_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8813 = 3'h4 == state ? _GEN_8249 : dirty_112_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8814 = 3'h4 == state ? _GEN_8250 : dirty_112_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8815 = 3'h4 == state ? _GEN_8251 : dirty_113_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8816 = 3'h4 == state ? _GEN_8252 : dirty_113_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8817 = 3'h4 == state ? _GEN_8253 : dirty_114_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8818 = 3'h4 == state ? _GEN_8254 : dirty_114_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8819 = 3'h4 == state ? _GEN_8255 : dirty_115_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8820 = 3'h4 == state ? _GEN_8256 : dirty_115_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8821 = 3'h4 == state ? _GEN_8257 : dirty_116_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8822 = 3'h4 == state ? _GEN_8258 : dirty_116_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8823 = 3'h4 == state ? _GEN_8259 : dirty_117_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8824 = 3'h4 == state ? _GEN_8260 : dirty_117_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8825 = 3'h4 == state ? _GEN_8261 : dirty_118_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8826 = 3'h4 == state ? _GEN_8262 : dirty_118_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8827 = 3'h4 == state ? _GEN_8263 : dirty_119_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8828 = 3'h4 == state ? _GEN_8264 : dirty_119_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8829 = 3'h4 == state ? _GEN_8265 : dirty_120_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8830 = 3'h4 == state ? _GEN_8266 : dirty_120_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8831 = 3'h4 == state ? _GEN_8267 : dirty_121_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8832 = 3'h4 == state ? _GEN_8268 : dirty_121_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8833 = 3'h4 == state ? _GEN_8269 : dirty_122_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8834 = 3'h4 == state ? _GEN_8270 : dirty_122_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8835 = 3'h4 == state ? _GEN_8271 : dirty_123_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8836 = 3'h4 == state ? _GEN_8272 : dirty_123_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8837 = 3'h4 == state ? _GEN_8273 : dirty_124_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8838 = 3'h4 == state ? _GEN_8274 : dirty_124_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8839 = 3'h4 == state ? _GEN_8275 : dirty_125_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8840 = 3'h4 == state ? _GEN_8276 : dirty_125_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8841 = 3'h4 == state ? _GEN_8277 : dirty_126_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8842 = 3'h4 == state ? _GEN_8278 : dirty_126_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8843 = 3'h4 == state ? _GEN_8279 : dirty_127_0; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8844 = 3'h4 == state ? _GEN_8280 : dirty_127_1; // @[DCache.scala 260:17 69:22]
  wire  _GEN_8845 = 3'h4 == state ? _GEN_8281 : replace_writeback; // @[DCache.scala 260:17 101:40]
  wire [31:0] _GEN_8846 = 3'h4 == state ? _GEN_8282 : ar_addr; // @[DCache.scala 260:17 199:24]
  wire [7:0] _GEN_8847 = 3'h4 == state ? _GEN_8283 : ar_len; // @[DCache.scala 260:17 199:24]
  wire [2:0] _GEN_8848 = 3'h4 == state ? _GEN_8284 : ar_size; // @[DCache.scala 260:17 199:24]
  wire  _GEN_8849 = 3'h4 == state ? _GEN_8285 : arvalid; // @[DCache.scala 260:17 200:24]
  wire  _GEN_8850 = 3'h4 == state ? _GEN_8286 : rready; // @[DCache.scala 260:17 203:23]
  wire  _GEN_8851 = 3'h4 == state ? _GEN_8287 : ar_handshake; // @[DCache.scala 260:17 99:40]
  wire [3:0] _GEN_8852 = 3'h4 == state ? _GEN_8288 : bram_replace_wea_0; // @[DCache.scala 260:17 73:33]
  wire [3:0] _GEN_8853 = 3'h4 == state ? _GEN_8289 : bram_replace_wea_1; // @[DCache.scala 260:17 73:33]
  wire  _GEN_8854 = 3'h4 == state ? _GEN_8290 : tag_wstrb_0; // @[DCache.scala 260:17 72:33]
  wire  _GEN_8855 = 3'h4 == state ? _GEN_8291 : tag_wstrb_1; // @[DCache.scala 260:17 72:33]
  wire [19:0] _GEN_8856 = 3'h4 == state ? _GEN_8292 : tag_wdata; // @[DCache.scala 260:17 77:26]
  wire [9:0] _GEN_8857 = 3'h4 == state ? _GEN_8293 : bram_replace_write_addr; // @[DCache.scala 260:17 92:40]
  wire  _GEN_8858 = 3'h4 == state ? _GEN_8294 : bram_use_replace_addr; // @[DCache.scala 260:17 95:40]
  wire  _GEN_8859 = 3'h4 == state ? _GEN_8295 : valid_0_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8860 = 3'h4 == state ? _GEN_8296 : valid_0_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8861 = 3'h4 == state ? _GEN_8297 : valid_1_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8862 = 3'h4 == state ? _GEN_8298 : valid_1_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8863 = 3'h4 == state ? _GEN_8299 : valid_2_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8864 = 3'h4 == state ? _GEN_8300 : valid_2_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8865 = 3'h4 == state ? _GEN_8301 : valid_3_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8866 = 3'h4 == state ? _GEN_8302 : valid_3_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8867 = 3'h4 == state ? _GEN_8303 : valid_4_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8868 = 3'h4 == state ? _GEN_8304 : valid_4_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8869 = 3'h4 == state ? _GEN_8305 : valid_5_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8870 = 3'h4 == state ? _GEN_8306 : valid_5_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8871 = 3'h4 == state ? _GEN_8307 : valid_6_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8872 = 3'h4 == state ? _GEN_8308 : valid_6_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8873 = 3'h4 == state ? _GEN_8309 : valid_7_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8874 = 3'h4 == state ? _GEN_8310 : valid_7_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8875 = 3'h4 == state ? _GEN_8311 : valid_8_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8876 = 3'h4 == state ? _GEN_8312 : valid_8_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8877 = 3'h4 == state ? _GEN_8313 : valid_9_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8878 = 3'h4 == state ? _GEN_8314 : valid_9_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8879 = 3'h4 == state ? _GEN_8315 : valid_10_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8880 = 3'h4 == state ? _GEN_8316 : valid_10_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8881 = 3'h4 == state ? _GEN_8317 : valid_11_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8882 = 3'h4 == state ? _GEN_8318 : valid_11_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8883 = 3'h4 == state ? _GEN_8319 : valid_12_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8884 = 3'h4 == state ? _GEN_8320 : valid_12_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8885 = 3'h4 == state ? _GEN_8321 : valid_13_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8886 = 3'h4 == state ? _GEN_8322 : valid_13_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8887 = 3'h4 == state ? _GEN_8323 : valid_14_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8888 = 3'h4 == state ? _GEN_8324 : valid_14_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8889 = 3'h4 == state ? _GEN_8325 : valid_15_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8890 = 3'h4 == state ? _GEN_8326 : valid_15_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8891 = 3'h4 == state ? _GEN_8327 : valid_16_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8892 = 3'h4 == state ? _GEN_8328 : valid_16_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8893 = 3'h4 == state ? _GEN_8329 : valid_17_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8894 = 3'h4 == state ? _GEN_8330 : valid_17_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8895 = 3'h4 == state ? _GEN_8331 : valid_18_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8896 = 3'h4 == state ? _GEN_8332 : valid_18_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8897 = 3'h4 == state ? _GEN_8333 : valid_19_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8898 = 3'h4 == state ? _GEN_8334 : valid_19_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8899 = 3'h4 == state ? _GEN_8335 : valid_20_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8900 = 3'h4 == state ? _GEN_8336 : valid_20_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8901 = 3'h4 == state ? _GEN_8337 : valid_21_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8902 = 3'h4 == state ? _GEN_8338 : valid_21_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8903 = 3'h4 == state ? _GEN_8339 : valid_22_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8904 = 3'h4 == state ? _GEN_8340 : valid_22_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8905 = 3'h4 == state ? _GEN_8341 : valid_23_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8906 = 3'h4 == state ? _GEN_8342 : valid_23_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8907 = 3'h4 == state ? _GEN_8343 : valid_24_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8908 = 3'h4 == state ? _GEN_8344 : valid_24_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8909 = 3'h4 == state ? _GEN_8345 : valid_25_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8910 = 3'h4 == state ? _GEN_8346 : valid_25_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8911 = 3'h4 == state ? _GEN_8347 : valid_26_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8912 = 3'h4 == state ? _GEN_8348 : valid_26_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8913 = 3'h4 == state ? _GEN_8349 : valid_27_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8914 = 3'h4 == state ? _GEN_8350 : valid_27_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8915 = 3'h4 == state ? _GEN_8351 : valid_28_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8916 = 3'h4 == state ? _GEN_8352 : valid_28_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8917 = 3'h4 == state ? _GEN_8353 : valid_29_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8918 = 3'h4 == state ? _GEN_8354 : valid_29_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8919 = 3'h4 == state ? _GEN_8355 : valid_30_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8920 = 3'h4 == state ? _GEN_8356 : valid_30_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8921 = 3'h4 == state ? _GEN_8357 : valid_31_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8922 = 3'h4 == state ? _GEN_8358 : valid_31_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8923 = 3'h4 == state ? _GEN_8359 : valid_32_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8924 = 3'h4 == state ? _GEN_8360 : valid_32_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8925 = 3'h4 == state ? _GEN_8361 : valid_33_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8926 = 3'h4 == state ? _GEN_8362 : valid_33_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8927 = 3'h4 == state ? _GEN_8363 : valid_34_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8928 = 3'h4 == state ? _GEN_8364 : valid_34_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8929 = 3'h4 == state ? _GEN_8365 : valid_35_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8930 = 3'h4 == state ? _GEN_8366 : valid_35_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8931 = 3'h4 == state ? _GEN_8367 : valid_36_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8932 = 3'h4 == state ? _GEN_8368 : valid_36_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8933 = 3'h4 == state ? _GEN_8369 : valid_37_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8934 = 3'h4 == state ? _GEN_8370 : valid_37_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8935 = 3'h4 == state ? _GEN_8371 : valid_38_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8936 = 3'h4 == state ? _GEN_8372 : valid_38_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8937 = 3'h4 == state ? _GEN_8373 : valid_39_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8938 = 3'h4 == state ? _GEN_8374 : valid_39_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8939 = 3'h4 == state ? _GEN_8375 : valid_40_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8940 = 3'h4 == state ? _GEN_8376 : valid_40_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8941 = 3'h4 == state ? _GEN_8377 : valid_41_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8942 = 3'h4 == state ? _GEN_8378 : valid_41_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8943 = 3'h4 == state ? _GEN_8379 : valid_42_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8944 = 3'h4 == state ? _GEN_8380 : valid_42_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8945 = 3'h4 == state ? _GEN_8381 : valid_43_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8946 = 3'h4 == state ? _GEN_8382 : valid_43_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8947 = 3'h4 == state ? _GEN_8383 : valid_44_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8948 = 3'h4 == state ? _GEN_8384 : valid_44_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8949 = 3'h4 == state ? _GEN_8385 : valid_45_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8950 = 3'h4 == state ? _GEN_8386 : valid_45_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8951 = 3'h4 == state ? _GEN_8387 : valid_46_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8952 = 3'h4 == state ? _GEN_8388 : valid_46_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8953 = 3'h4 == state ? _GEN_8389 : valid_47_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8954 = 3'h4 == state ? _GEN_8390 : valid_47_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8955 = 3'h4 == state ? _GEN_8391 : valid_48_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8956 = 3'h4 == state ? _GEN_8392 : valid_48_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8957 = 3'h4 == state ? _GEN_8393 : valid_49_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8958 = 3'h4 == state ? _GEN_8394 : valid_49_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8959 = 3'h4 == state ? _GEN_8395 : valid_50_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8960 = 3'h4 == state ? _GEN_8396 : valid_50_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8961 = 3'h4 == state ? _GEN_8397 : valid_51_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8962 = 3'h4 == state ? _GEN_8398 : valid_51_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8963 = 3'h4 == state ? _GEN_8399 : valid_52_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8964 = 3'h4 == state ? _GEN_8400 : valid_52_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8965 = 3'h4 == state ? _GEN_8401 : valid_53_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8966 = 3'h4 == state ? _GEN_8402 : valid_53_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8967 = 3'h4 == state ? _GEN_8403 : valid_54_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8968 = 3'h4 == state ? _GEN_8404 : valid_54_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8969 = 3'h4 == state ? _GEN_8405 : valid_55_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8970 = 3'h4 == state ? _GEN_8406 : valid_55_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8971 = 3'h4 == state ? _GEN_8407 : valid_56_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8972 = 3'h4 == state ? _GEN_8408 : valid_56_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8973 = 3'h4 == state ? _GEN_8409 : valid_57_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8974 = 3'h4 == state ? _GEN_8410 : valid_57_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8975 = 3'h4 == state ? _GEN_8411 : valid_58_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8976 = 3'h4 == state ? _GEN_8412 : valid_58_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8977 = 3'h4 == state ? _GEN_8413 : valid_59_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8978 = 3'h4 == state ? _GEN_8414 : valid_59_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8979 = 3'h4 == state ? _GEN_8415 : valid_60_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8980 = 3'h4 == state ? _GEN_8416 : valid_60_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8981 = 3'h4 == state ? _GEN_8417 : valid_61_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8982 = 3'h4 == state ? _GEN_8418 : valid_61_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8983 = 3'h4 == state ? _GEN_8419 : valid_62_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8984 = 3'h4 == state ? _GEN_8420 : valid_62_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8985 = 3'h4 == state ? _GEN_8421 : valid_63_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8986 = 3'h4 == state ? _GEN_8422 : valid_63_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8987 = 3'h4 == state ? _GEN_8423 : valid_64_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8988 = 3'h4 == state ? _GEN_8424 : valid_64_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8989 = 3'h4 == state ? _GEN_8425 : valid_65_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8990 = 3'h4 == state ? _GEN_8426 : valid_65_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8991 = 3'h4 == state ? _GEN_8427 : valid_66_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8992 = 3'h4 == state ? _GEN_8428 : valid_66_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8993 = 3'h4 == state ? _GEN_8429 : valid_67_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8994 = 3'h4 == state ? _GEN_8430 : valid_67_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8995 = 3'h4 == state ? _GEN_8431 : valid_68_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8996 = 3'h4 == state ? _GEN_8432 : valid_68_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8997 = 3'h4 == state ? _GEN_8433 : valid_69_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8998 = 3'h4 == state ? _GEN_8434 : valid_69_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_8999 = 3'h4 == state ? _GEN_8435 : valid_70_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9000 = 3'h4 == state ? _GEN_8436 : valid_70_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9001 = 3'h4 == state ? _GEN_8437 : valid_71_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9002 = 3'h4 == state ? _GEN_8438 : valid_71_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9003 = 3'h4 == state ? _GEN_8439 : valid_72_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9004 = 3'h4 == state ? _GEN_8440 : valid_72_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9005 = 3'h4 == state ? _GEN_8441 : valid_73_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9006 = 3'h4 == state ? _GEN_8442 : valid_73_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9007 = 3'h4 == state ? _GEN_8443 : valid_74_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9008 = 3'h4 == state ? _GEN_8444 : valid_74_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9009 = 3'h4 == state ? _GEN_8445 : valid_75_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9010 = 3'h4 == state ? _GEN_8446 : valid_75_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9011 = 3'h4 == state ? _GEN_8447 : valid_76_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9012 = 3'h4 == state ? _GEN_8448 : valid_76_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9013 = 3'h4 == state ? _GEN_8449 : valid_77_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9014 = 3'h4 == state ? _GEN_8450 : valid_77_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9015 = 3'h4 == state ? _GEN_8451 : valid_78_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9016 = 3'h4 == state ? _GEN_8452 : valid_78_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9017 = 3'h4 == state ? _GEN_8453 : valid_79_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9018 = 3'h4 == state ? _GEN_8454 : valid_79_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9019 = 3'h4 == state ? _GEN_8455 : valid_80_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9020 = 3'h4 == state ? _GEN_8456 : valid_80_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9021 = 3'h4 == state ? _GEN_8457 : valid_81_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9022 = 3'h4 == state ? _GEN_8458 : valid_81_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9023 = 3'h4 == state ? _GEN_8459 : valid_82_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9024 = 3'h4 == state ? _GEN_8460 : valid_82_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9025 = 3'h4 == state ? _GEN_8461 : valid_83_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9026 = 3'h4 == state ? _GEN_8462 : valid_83_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9027 = 3'h4 == state ? _GEN_8463 : valid_84_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9028 = 3'h4 == state ? _GEN_8464 : valid_84_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9029 = 3'h4 == state ? _GEN_8465 : valid_85_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9030 = 3'h4 == state ? _GEN_8466 : valid_85_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9031 = 3'h4 == state ? _GEN_8467 : valid_86_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9032 = 3'h4 == state ? _GEN_8468 : valid_86_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9033 = 3'h4 == state ? _GEN_8469 : valid_87_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9034 = 3'h4 == state ? _GEN_8470 : valid_87_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9035 = 3'h4 == state ? _GEN_8471 : valid_88_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9036 = 3'h4 == state ? _GEN_8472 : valid_88_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9037 = 3'h4 == state ? _GEN_8473 : valid_89_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9038 = 3'h4 == state ? _GEN_8474 : valid_89_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9039 = 3'h4 == state ? _GEN_8475 : valid_90_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9040 = 3'h4 == state ? _GEN_8476 : valid_90_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9041 = 3'h4 == state ? _GEN_8477 : valid_91_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9042 = 3'h4 == state ? _GEN_8478 : valid_91_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9043 = 3'h4 == state ? _GEN_8479 : valid_92_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9044 = 3'h4 == state ? _GEN_8480 : valid_92_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9045 = 3'h4 == state ? _GEN_8481 : valid_93_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9046 = 3'h4 == state ? _GEN_8482 : valid_93_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9047 = 3'h4 == state ? _GEN_8483 : valid_94_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9048 = 3'h4 == state ? _GEN_8484 : valid_94_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9049 = 3'h4 == state ? _GEN_8485 : valid_95_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9050 = 3'h4 == state ? _GEN_8486 : valid_95_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9051 = 3'h4 == state ? _GEN_8487 : valid_96_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9052 = 3'h4 == state ? _GEN_8488 : valid_96_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9053 = 3'h4 == state ? _GEN_8489 : valid_97_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9054 = 3'h4 == state ? _GEN_8490 : valid_97_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9055 = 3'h4 == state ? _GEN_8491 : valid_98_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9056 = 3'h4 == state ? _GEN_8492 : valid_98_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9057 = 3'h4 == state ? _GEN_8493 : valid_99_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9058 = 3'h4 == state ? _GEN_8494 : valid_99_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9059 = 3'h4 == state ? _GEN_8495 : valid_100_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9060 = 3'h4 == state ? _GEN_8496 : valid_100_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9061 = 3'h4 == state ? _GEN_8497 : valid_101_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9062 = 3'h4 == state ? _GEN_8498 : valid_101_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9063 = 3'h4 == state ? _GEN_8499 : valid_102_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9064 = 3'h4 == state ? _GEN_8500 : valid_102_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9065 = 3'h4 == state ? _GEN_8501 : valid_103_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9066 = 3'h4 == state ? _GEN_8502 : valid_103_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9067 = 3'h4 == state ? _GEN_8503 : valid_104_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9068 = 3'h4 == state ? _GEN_8504 : valid_104_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9069 = 3'h4 == state ? _GEN_8505 : valid_105_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9070 = 3'h4 == state ? _GEN_8506 : valid_105_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9071 = 3'h4 == state ? _GEN_8507 : valid_106_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9072 = 3'h4 == state ? _GEN_8508 : valid_106_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9073 = 3'h4 == state ? _GEN_8509 : valid_107_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9074 = 3'h4 == state ? _GEN_8510 : valid_107_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9075 = 3'h4 == state ? _GEN_8511 : valid_108_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9076 = 3'h4 == state ? _GEN_8512 : valid_108_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9077 = 3'h4 == state ? _GEN_8513 : valid_109_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9078 = 3'h4 == state ? _GEN_8514 : valid_109_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9079 = 3'h4 == state ? _GEN_8515 : valid_110_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9080 = 3'h4 == state ? _GEN_8516 : valid_110_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9081 = 3'h4 == state ? _GEN_8517 : valid_111_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9082 = 3'h4 == state ? _GEN_8518 : valid_111_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9083 = 3'h4 == state ? _GEN_8519 : valid_112_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9084 = 3'h4 == state ? _GEN_8520 : valid_112_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9085 = 3'h4 == state ? _GEN_8521 : valid_113_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9086 = 3'h4 == state ? _GEN_8522 : valid_113_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9087 = 3'h4 == state ? _GEN_8523 : valid_114_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9088 = 3'h4 == state ? _GEN_8524 : valid_114_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9089 = 3'h4 == state ? _GEN_8525 : valid_115_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9090 = 3'h4 == state ? _GEN_8526 : valid_115_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9091 = 3'h4 == state ? _GEN_8527 : valid_116_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9092 = 3'h4 == state ? _GEN_8528 : valid_116_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9093 = 3'h4 == state ? _GEN_8529 : valid_117_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9094 = 3'h4 == state ? _GEN_8530 : valid_117_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9095 = 3'h4 == state ? _GEN_8531 : valid_118_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9096 = 3'h4 == state ? _GEN_8532 : valid_118_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9097 = 3'h4 == state ? _GEN_8533 : valid_119_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9098 = 3'h4 == state ? _GEN_8534 : valid_119_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9099 = 3'h4 == state ? _GEN_8535 : valid_120_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9100 = 3'h4 == state ? _GEN_8536 : valid_120_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9101 = 3'h4 == state ? _GEN_8537 : valid_121_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9102 = 3'h4 == state ? _GEN_8538 : valid_121_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9103 = 3'h4 == state ? _GEN_8539 : valid_122_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9104 = 3'h4 == state ? _GEN_8540 : valid_122_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9105 = 3'h4 == state ? _GEN_8541 : valid_123_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9106 = 3'h4 == state ? _GEN_8542 : valid_123_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9107 = 3'h4 == state ? _GEN_8543 : valid_124_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9108 = 3'h4 == state ? _GEN_8544 : valid_124_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9109 = 3'h4 == state ? _GEN_8545 : valid_125_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9110 = 3'h4 == state ? _GEN_8546 : valid_125_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9111 = 3'h4 == state ? _GEN_8547 : valid_126_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9112 = 3'h4 == state ? _GEN_8548 : valid_126_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9113 = 3'h4 == state ? _GEN_8549 : valid_127_0; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9114 = 3'h4 == state ? _GEN_8550 : valid_127_1; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9115 = 3'h4 == state ? _GEN_8551 : replace_working; // @[DCache.scala 260:17 98:40]
  wire [2:0] _GEN_9116 = 3'h4 == state ? _GEN_8552 : _GEN_8557; // @[DCache.scala 260:17]
  wire  _GEN_9117 = 3'h4 == state ? data_tlb_invalid : _GEN_8558; // @[DCache.scala 260:17 250:25]
  wire  _GEN_9118 = 3'h4 == state ? data_tlb_refill : _GEN_8559; // @[DCache.scala 260:17 250:25]
  wire  _GEN_9119 = 3'h4 == state ? data_tlb_mod : _GEN_8560; // @[DCache.scala 260:17 250:25]
  wire [9:0] _GEN_9120 = 3'h3 == state ? _GEN_5751 : _GEN_8561; // @[DCache.scala 260:17]
  wire [9:0] _GEN_9121 = 3'h3 == state ? _GEN_5752 : _GEN_8562; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9122 = 3'h3 == state ? _GEN_5753 : _GEN_8563; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9123 = 3'h3 == state ? _GEN_5754 : _GEN_8564; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9124 = 3'h3 == state ? _GEN_5755 : _GEN_8565; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9125 = 3'h3 == state ? _GEN_5756 : _GEN_8566; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9126 = 3'h3 == state ? _GEN_5757 : _GEN_8567; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9127 = 3'h3 == state ? _GEN_5758 : _GEN_8568; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9128 = 3'h3 == state ? _GEN_5759 : _GEN_8569; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9129 = 3'h3 == state ? _GEN_5760 : _GEN_8570; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9130 = 3'h3 == state ? _GEN_5761 : _GEN_8571; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9131 = 3'h3 == state ? _GEN_5762 : _GEN_8572; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9132 = 3'h3 == state ? _GEN_5763 : _GEN_8573; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9133 = 3'h3 == state ? _GEN_5764 : _GEN_8574; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9134 = 3'h3 == state ? _GEN_5765 : _GEN_8575; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9135 = 3'h3 == state ? _GEN_5766 : _GEN_8576; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9136 = 3'h3 == state ? _GEN_5767 : _GEN_8577; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9137 = 3'h3 == state ? _GEN_5768 : _GEN_8578; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9138 = 3'h3 == state ? _GEN_5769 : _GEN_8579; // @[DCache.scala 260:17]
  wire [7:0] _GEN_9139 = 3'h3 == state ? _GEN_5770 : _GEN_8580; // @[DCache.scala 260:17]
  wire [2:0] _GEN_9140 = 3'h3 == state ? _GEN_5771 : _GEN_8581; // @[DCache.scala 260:17]
  wire  _GEN_9141 = 3'h3 == state ? _GEN_5772 : _GEN_8582; // @[DCache.scala 260:17]
  wire [31:0] _GEN_9142 = 3'h3 == state ? _GEN_5773 : _GEN_8583; // @[DCache.scala 260:17]
  wire [3:0] _GEN_9143 = 3'h3 == state ? _GEN_5774 : _GEN_8584; // @[DCache.scala 260:17]
  wire  _GEN_9144 = 3'h3 == state ? _GEN_5775 : _GEN_8585; // @[DCache.scala 260:17]
  wire  _GEN_9145 = 3'h3 == state ? _GEN_5776 : _GEN_8586; // @[DCache.scala 260:17]
  wire  _GEN_9146 = 3'h3 == state ? _GEN_5777 : _GEN_8587; // @[DCache.scala 260:17]
  wire [3:0] _GEN_9147 = 3'h3 == state ? _GEN_5778 : _GEN_8588; // @[DCache.scala 260:17]
  wire  _GEN_9148 = 3'h3 == state ? _GEN_5779 : _GEN_8589; // @[DCache.scala 260:17]
  wire  _GEN_9149 = 3'h3 == state ? _GEN_5780 : _GEN_8590; // @[DCache.scala 260:17]
  wire  _GEN_9150 = 3'h3 == state ? _GEN_5781 : _GEN_8591; // @[DCache.scala 260:17]
  wire  _GEN_9151 = 3'h3 == state ? _GEN_5782 : _GEN_8592; // @[DCache.scala 260:17]
  wire  _GEN_9152 = 3'h3 == state ? _GEN_5783 : _GEN_8593; // @[DCache.scala 260:17]
  wire  _GEN_9153 = 3'h3 == state ? _GEN_5784 : _GEN_8594; // @[DCache.scala 260:17]
  wire  _GEN_9154 = 3'h3 == state ? _GEN_5785 : _GEN_8595; // @[DCache.scala 260:17]
  wire  _GEN_9155 = 3'h3 == state ? _GEN_5786 : _GEN_8596; // @[DCache.scala 260:17]
  wire  _GEN_9156 = 3'h3 == state ? _GEN_5787 : _GEN_8597; // @[DCache.scala 260:17]
  wire  _GEN_9157 = 3'h3 == state ? _GEN_5788 : _GEN_8598; // @[DCache.scala 260:17]
  wire  _GEN_9158 = 3'h3 == state ? _GEN_5789 : _GEN_8599; // @[DCache.scala 260:17]
  wire  _GEN_9159 = 3'h3 == state ? _GEN_5790 : _GEN_8600; // @[DCache.scala 260:17]
  wire  _GEN_9160 = 3'h3 == state ? _GEN_5791 : _GEN_8601; // @[DCache.scala 260:17]
  wire  _GEN_9161 = 3'h3 == state ? _GEN_5792 : _GEN_8602; // @[DCache.scala 260:17]
  wire  _GEN_9162 = 3'h3 == state ? _GEN_5793 : _GEN_8603; // @[DCache.scala 260:17]
  wire  _GEN_9163 = 3'h3 == state ? _GEN_5794 : _GEN_8604; // @[DCache.scala 260:17]
  wire  _GEN_9164 = 3'h3 == state ? _GEN_5795 : _GEN_8605; // @[DCache.scala 260:17]
  wire  _GEN_9165 = 3'h3 == state ? _GEN_5796 : _GEN_8606; // @[DCache.scala 260:17]
  wire  _GEN_9166 = 3'h3 == state ? _GEN_5797 : _GEN_8607; // @[DCache.scala 260:17]
  wire  _GEN_9167 = 3'h3 == state ? _GEN_5798 : _GEN_8608; // @[DCache.scala 260:17]
  wire  _GEN_9168 = 3'h3 == state ? _GEN_5799 : _GEN_8609; // @[DCache.scala 260:17]
  wire  _GEN_9169 = 3'h3 == state ? _GEN_5800 : _GEN_8610; // @[DCache.scala 260:17]
  wire  _GEN_9170 = 3'h3 == state ? _GEN_5801 : _GEN_8611; // @[DCache.scala 260:17]
  wire  _GEN_9171 = 3'h3 == state ? _GEN_5802 : _GEN_8612; // @[DCache.scala 260:17]
  wire  _GEN_9172 = 3'h3 == state ? _GEN_5803 : _GEN_8613; // @[DCache.scala 260:17]
  wire  _GEN_9173 = 3'h3 == state ? _GEN_5804 : _GEN_8614; // @[DCache.scala 260:17]
  wire  _GEN_9174 = 3'h3 == state ? _GEN_5805 : _GEN_8615; // @[DCache.scala 260:17]
  wire  _GEN_9175 = 3'h3 == state ? _GEN_5806 : _GEN_8616; // @[DCache.scala 260:17]
  wire  _GEN_9176 = 3'h3 == state ? _GEN_5807 : _GEN_8617; // @[DCache.scala 260:17]
  wire  _GEN_9177 = 3'h3 == state ? _GEN_5808 : _GEN_8618; // @[DCache.scala 260:17]
  wire  _GEN_9178 = 3'h3 == state ? _GEN_5809 : _GEN_8619; // @[DCache.scala 260:17]
  wire  _GEN_9179 = 3'h3 == state ? _GEN_5810 : _GEN_8620; // @[DCache.scala 260:17]
  wire  _GEN_9180 = 3'h3 == state ? _GEN_5811 : _GEN_8621; // @[DCache.scala 260:17]
  wire  _GEN_9181 = 3'h3 == state ? _GEN_5812 : _GEN_8622; // @[DCache.scala 260:17]
  wire  _GEN_9182 = 3'h3 == state ? _GEN_5813 : _GEN_8623; // @[DCache.scala 260:17]
  wire  _GEN_9183 = 3'h3 == state ? _GEN_5814 : _GEN_8624; // @[DCache.scala 260:17]
  wire  _GEN_9184 = 3'h3 == state ? _GEN_5815 : _GEN_8625; // @[DCache.scala 260:17]
  wire  _GEN_9185 = 3'h3 == state ? _GEN_5816 : _GEN_8626; // @[DCache.scala 260:17]
  wire  _GEN_9186 = 3'h3 == state ? _GEN_5817 : _GEN_8627; // @[DCache.scala 260:17]
  wire  _GEN_9187 = 3'h3 == state ? _GEN_5818 : _GEN_8628; // @[DCache.scala 260:17]
  wire  _GEN_9188 = 3'h3 == state ? _GEN_5819 : _GEN_8629; // @[DCache.scala 260:17]
  wire  _GEN_9189 = 3'h3 == state ? _GEN_5820 : _GEN_8630; // @[DCache.scala 260:17]
  wire  _GEN_9190 = 3'h3 == state ? _GEN_5821 : _GEN_8631; // @[DCache.scala 260:17]
  wire  _GEN_9191 = 3'h3 == state ? _GEN_5822 : _GEN_8632; // @[DCache.scala 260:17]
  wire  _GEN_9192 = 3'h3 == state ? _GEN_5823 : _GEN_8633; // @[DCache.scala 260:17]
  wire  _GEN_9193 = 3'h3 == state ? _GEN_5824 : _GEN_8634; // @[DCache.scala 260:17]
  wire  _GEN_9194 = 3'h3 == state ? _GEN_5825 : _GEN_8635; // @[DCache.scala 260:17]
  wire  _GEN_9195 = 3'h3 == state ? _GEN_5826 : _GEN_8636; // @[DCache.scala 260:17]
  wire  _GEN_9196 = 3'h3 == state ? _GEN_5827 : _GEN_8637; // @[DCache.scala 260:17]
  wire  _GEN_9197 = 3'h3 == state ? _GEN_5828 : _GEN_8638; // @[DCache.scala 260:17]
  wire  _GEN_9198 = 3'h3 == state ? _GEN_5829 : _GEN_8639; // @[DCache.scala 260:17]
  wire  _GEN_9199 = 3'h3 == state ? _GEN_5830 : _GEN_8640; // @[DCache.scala 260:17]
  wire  _GEN_9200 = 3'h3 == state ? _GEN_5831 : _GEN_8641; // @[DCache.scala 260:17]
  wire  _GEN_9201 = 3'h3 == state ? _GEN_5832 : _GEN_8642; // @[DCache.scala 260:17]
  wire  _GEN_9202 = 3'h3 == state ? _GEN_5833 : _GEN_8643; // @[DCache.scala 260:17]
  wire  _GEN_9203 = 3'h3 == state ? _GEN_5834 : _GEN_8644; // @[DCache.scala 260:17]
  wire  _GEN_9204 = 3'h3 == state ? _GEN_5835 : _GEN_8645; // @[DCache.scala 260:17]
  wire  _GEN_9205 = 3'h3 == state ? _GEN_5836 : _GEN_8646; // @[DCache.scala 260:17]
  wire  _GEN_9206 = 3'h3 == state ? _GEN_5837 : _GEN_8647; // @[DCache.scala 260:17]
  wire  _GEN_9207 = 3'h3 == state ? _GEN_5838 : _GEN_8648; // @[DCache.scala 260:17]
  wire  _GEN_9208 = 3'h3 == state ? _GEN_5839 : _GEN_8649; // @[DCache.scala 260:17]
  wire  _GEN_9209 = 3'h3 == state ? _GEN_5840 : _GEN_8650; // @[DCache.scala 260:17]
  wire  _GEN_9210 = 3'h3 == state ? _GEN_5841 : _GEN_8651; // @[DCache.scala 260:17]
  wire  _GEN_9211 = 3'h3 == state ? _GEN_5842 : _GEN_8652; // @[DCache.scala 260:17]
  wire  _GEN_9212 = 3'h3 == state ? _GEN_5843 : _GEN_8653; // @[DCache.scala 260:17]
  wire  _GEN_9213 = 3'h3 == state ? _GEN_5844 : _GEN_8654; // @[DCache.scala 260:17]
  wire  _GEN_9214 = 3'h3 == state ? _GEN_5845 : _GEN_8655; // @[DCache.scala 260:17]
  wire  _GEN_9215 = 3'h3 == state ? _GEN_5846 : _GEN_8656; // @[DCache.scala 260:17]
  wire  _GEN_9216 = 3'h3 == state ? _GEN_5847 : _GEN_8657; // @[DCache.scala 260:17]
  wire  _GEN_9217 = 3'h3 == state ? _GEN_5848 : _GEN_8658; // @[DCache.scala 260:17]
  wire  _GEN_9218 = 3'h3 == state ? _GEN_5849 : _GEN_8659; // @[DCache.scala 260:17]
  wire  _GEN_9219 = 3'h3 == state ? _GEN_5850 : _GEN_8660; // @[DCache.scala 260:17]
  wire  _GEN_9220 = 3'h3 == state ? _GEN_5851 : _GEN_8661; // @[DCache.scala 260:17]
  wire  _GEN_9221 = 3'h3 == state ? _GEN_5852 : _GEN_8662; // @[DCache.scala 260:17]
  wire  _GEN_9222 = 3'h3 == state ? _GEN_5853 : _GEN_8663; // @[DCache.scala 260:17]
  wire  _GEN_9223 = 3'h3 == state ? _GEN_5854 : _GEN_8664; // @[DCache.scala 260:17]
  wire  _GEN_9224 = 3'h3 == state ? _GEN_5855 : _GEN_8665; // @[DCache.scala 260:17]
  wire  _GEN_9225 = 3'h3 == state ? _GEN_5856 : _GEN_8666; // @[DCache.scala 260:17]
  wire  _GEN_9226 = 3'h3 == state ? _GEN_5857 : _GEN_8667; // @[DCache.scala 260:17]
  wire  _GEN_9227 = 3'h3 == state ? _GEN_5858 : _GEN_8668; // @[DCache.scala 260:17]
  wire  _GEN_9228 = 3'h3 == state ? _GEN_5859 : _GEN_8669; // @[DCache.scala 260:17]
  wire  _GEN_9229 = 3'h3 == state ? _GEN_5860 : _GEN_8670; // @[DCache.scala 260:17]
  wire  _GEN_9230 = 3'h3 == state ? _GEN_5861 : _GEN_8671; // @[DCache.scala 260:17]
  wire  _GEN_9231 = 3'h3 == state ? _GEN_5862 : _GEN_8672; // @[DCache.scala 260:17]
  wire  _GEN_9232 = 3'h3 == state ? _GEN_5863 : _GEN_8673; // @[DCache.scala 260:17]
  wire  _GEN_9233 = 3'h3 == state ? _GEN_5864 : _GEN_8674; // @[DCache.scala 260:17]
  wire  _GEN_9234 = 3'h3 == state ? _GEN_5865 : _GEN_8675; // @[DCache.scala 260:17]
  wire  _GEN_9235 = 3'h3 == state ? _GEN_5866 : _GEN_8676; // @[DCache.scala 260:17]
  wire  _GEN_9236 = 3'h3 == state ? _GEN_5867 : _GEN_8677; // @[DCache.scala 260:17]
  wire  _GEN_9237 = 3'h3 == state ? _GEN_5868 : _GEN_8678; // @[DCache.scala 260:17]
  wire  _GEN_9238 = 3'h3 == state ? _GEN_5869 : _GEN_8679; // @[DCache.scala 260:17]
  wire  _GEN_9239 = 3'h3 == state ? _GEN_5870 : _GEN_8680; // @[DCache.scala 260:17]
  wire  _GEN_9240 = 3'h3 == state ? _GEN_5871 : _GEN_8681; // @[DCache.scala 260:17]
  wire  _GEN_9241 = 3'h3 == state ? _GEN_5872 : _GEN_8682; // @[DCache.scala 260:17]
  wire  _GEN_9242 = 3'h3 == state ? _GEN_5873 : _GEN_8683; // @[DCache.scala 260:17]
  wire  _GEN_9243 = 3'h3 == state ? _GEN_5874 : _GEN_8684; // @[DCache.scala 260:17]
  wire  _GEN_9244 = 3'h3 == state ? _GEN_5875 : _GEN_8685; // @[DCache.scala 260:17]
  wire  _GEN_9245 = 3'h3 == state ? _GEN_5876 : _GEN_8686; // @[DCache.scala 260:17]
  wire  _GEN_9246 = 3'h3 == state ? _GEN_5877 : _GEN_8687; // @[DCache.scala 260:17]
  wire  _GEN_9247 = 3'h3 == state ? _GEN_5878 : _GEN_8688; // @[DCache.scala 260:17]
  wire  _GEN_9248 = 3'h3 == state ? _GEN_5879 : _GEN_8689; // @[DCache.scala 260:17]
  wire  _GEN_9249 = 3'h3 == state ? _GEN_5880 : _GEN_8690; // @[DCache.scala 260:17]
  wire  _GEN_9250 = 3'h3 == state ? _GEN_5881 : _GEN_8691; // @[DCache.scala 260:17]
  wire  _GEN_9251 = 3'h3 == state ? _GEN_5882 : _GEN_8692; // @[DCache.scala 260:17]
  wire  _GEN_9252 = 3'h3 == state ? _GEN_5883 : _GEN_8693; // @[DCache.scala 260:17]
  wire  _GEN_9253 = 3'h3 == state ? _GEN_5884 : _GEN_8694; // @[DCache.scala 260:17]
  wire  _GEN_9254 = 3'h3 == state ? _GEN_5885 : _GEN_8695; // @[DCache.scala 260:17]
  wire  _GEN_9255 = 3'h3 == state ? _GEN_5886 : _GEN_8696; // @[DCache.scala 260:17]
  wire  _GEN_9256 = 3'h3 == state ? _GEN_5887 : _GEN_8697; // @[DCache.scala 260:17]
  wire  _GEN_9257 = 3'h3 == state ? _GEN_5888 : _GEN_8698; // @[DCache.scala 260:17]
  wire  _GEN_9258 = 3'h3 == state ? _GEN_5889 : _GEN_8699; // @[DCache.scala 260:17]
  wire  _GEN_9259 = 3'h3 == state ? _GEN_5890 : _GEN_8700; // @[DCache.scala 260:17]
  wire  _GEN_9260 = 3'h3 == state ? _GEN_5891 : _GEN_8701; // @[DCache.scala 260:17]
  wire  _GEN_9261 = 3'h3 == state ? _GEN_5892 : _GEN_8702; // @[DCache.scala 260:17]
  wire  _GEN_9262 = 3'h3 == state ? _GEN_5893 : _GEN_8703; // @[DCache.scala 260:17]
  wire  _GEN_9263 = 3'h3 == state ? _GEN_5894 : _GEN_8704; // @[DCache.scala 260:17]
  wire  _GEN_9264 = 3'h3 == state ? _GEN_5895 : _GEN_8705; // @[DCache.scala 260:17]
  wire  _GEN_9265 = 3'h3 == state ? _GEN_5896 : _GEN_8706; // @[DCache.scala 260:17]
  wire  _GEN_9266 = 3'h3 == state ? _GEN_5897 : _GEN_8707; // @[DCache.scala 260:17]
  wire  _GEN_9267 = 3'h3 == state ? _GEN_5898 : _GEN_8708; // @[DCache.scala 260:17]
  wire  _GEN_9268 = 3'h3 == state ? _GEN_5899 : _GEN_8709; // @[DCache.scala 260:17]
  wire  _GEN_9269 = 3'h3 == state ? _GEN_5900 : _GEN_8710; // @[DCache.scala 260:17]
  wire  _GEN_9270 = 3'h3 == state ? _GEN_5901 : _GEN_8711; // @[DCache.scala 260:17]
  wire  _GEN_9271 = 3'h3 == state ? _GEN_5902 : _GEN_8712; // @[DCache.scala 260:17]
  wire  _GEN_9272 = 3'h3 == state ? _GEN_5903 : _GEN_8713; // @[DCache.scala 260:17]
  wire  _GEN_9273 = 3'h3 == state ? _GEN_5904 : _GEN_8714; // @[DCache.scala 260:17]
  wire  _GEN_9274 = 3'h3 == state ? _GEN_5905 : _GEN_8715; // @[DCache.scala 260:17]
  wire  _GEN_9275 = 3'h3 == state ? _GEN_5906 : _GEN_8716; // @[DCache.scala 260:17]
  wire  _GEN_9276 = 3'h3 == state ? _GEN_5907 : _GEN_8717; // @[DCache.scala 260:17]
  wire  _GEN_9277 = 3'h3 == state ? _GEN_5908 : _GEN_8718; // @[DCache.scala 260:17]
  wire  _GEN_9278 = 3'h3 == state ? _GEN_5909 : _GEN_8719; // @[DCache.scala 260:17]
  wire  _GEN_9279 = 3'h3 == state ? _GEN_5910 : _GEN_8720; // @[DCache.scala 260:17]
  wire  _GEN_9280 = 3'h3 == state ? _GEN_5911 : _GEN_8721; // @[DCache.scala 260:17]
  wire  _GEN_9281 = 3'h3 == state ? _GEN_5912 : _GEN_8722; // @[DCache.scala 260:17]
  wire  _GEN_9282 = 3'h3 == state ? _GEN_5913 : _GEN_8723; // @[DCache.scala 260:17]
  wire  _GEN_9283 = 3'h3 == state ? _GEN_5914 : _GEN_8724; // @[DCache.scala 260:17]
  wire  _GEN_9284 = 3'h3 == state ? _GEN_5915 : _GEN_8725; // @[DCache.scala 260:17]
  wire  _GEN_9285 = 3'h3 == state ? _GEN_5916 : _GEN_8726; // @[DCache.scala 260:17]
  wire  _GEN_9286 = 3'h3 == state ? _GEN_5917 : _GEN_8727; // @[DCache.scala 260:17]
  wire  _GEN_9287 = 3'h3 == state ? _GEN_5918 : _GEN_8728; // @[DCache.scala 260:17]
  wire  _GEN_9288 = 3'h3 == state ? _GEN_5919 : _GEN_8729; // @[DCache.scala 260:17]
  wire  _GEN_9289 = 3'h3 == state ? _GEN_5920 : _GEN_8730; // @[DCache.scala 260:17]
  wire  _GEN_9290 = 3'h3 == state ? _GEN_5921 : _GEN_8731; // @[DCache.scala 260:17]
  wire  _GEN_9291 = 3'h3 == state ? _GEN_5922 : _GEN_8732; // @[DCache.scala 260:17]
  wire  _GEN_9292 = 3'h3 == state ? _GEN_5923 : _GEN_8733; // @[DCache.scala 260:17]
  wire  _GEN_9293 = 3'h3 == state ? _GEN_5924 : _GEN_8734; // @[DCache.scala 260:17]
  wire  _GEN_9294 = 3'h3 == state ? _GEN_5925 : _GEN_8735; // @[DCache.scala 260:17]
  wire  _GEN_9295 = 3'h3 == state ? _GEN_5926 : _GEN_8736; // @[DCache.scala 260:17]
  wire  _GEN_9296 = 3'h3 == state ? _GEN_5927 : _GEN_8737; // @[DCache.scala 260:17]
  wire  _GEN_9297 = 3'h3 == state ? _GEN_5928 : _GEN_8738; // @[DCache.scala 260:17]
  wire  _GEN_9298 = 3'h3 == state ? _GEN_5929 : _GEN_8739; // @[DCache.scala 260:17]
  wire  _GEN_9299 = 3'h3 == state ? _GEN_5930 : _GEN_8740; // @[DCache.scala 260:17]
  wire  _GEN_9300 = 3'h3 == state ? _GEN_5931 : _GEN_8741; // @[DCache.scala 260:17]
  wire  _GEN_9301 = 3'h3 == state ? _GEN_5932 : _GEN_8742; // @[DCache.scala 260:17]
  wire  _GEN_9302 = 3'h3 == state ? _GEN_5933 : _GEN_8743; // @[DCache.scala 260:17]
  wire  _GEN_9303 = 3'h3 == state ? _GEN_5934 : _GEN_8744; // @[DCache.scala 260:17]
  wire  _GEN_9304 = 3'h3 == state ? _GEN_5935 : _GEN_8745; // @[DCache.scala 260:17]
  wire  _GEN_9305 = 3'h3 == state ? _GEN_5936 : _GEN_8746; // @[DCache.scala 260:17]
  wire  _GEN_9306 = 3'h3 == state ? _GEN_5937 : _GEN_8747; // @[DCache.scala 260:17]
  wire  _GEN_9307 = 3'h3 == state ? _GEN_5938 : _GEN_8748; // @[DCache.scala 260:17]
  wire  _GEN_9308 = 3'h3 == state ? _GEN_5939 : _GEN_8749; // @[DCache.scala 260:17]
  wire  _GEN_9309 = 3'h3 == state ? _GEN_5940 : _GEN_8750; // @[DCache.scala 260:17]
  wire  _GEN_9310 = 3'h3 == state ? _GEN_5941 : _GEN_8751; // @[DCache.scala 260:17]
  wire  _GEN_9311 = 3'h3 == state ? _GEN_5942 : _GEN_8752; // @[DCache.scala 260:17]
  wire  _GEN_9312 = 3'h3 == state ? _GEN_5943 : _GEN_8753; // @[DCache.scala 260:17]
  wire  _GEN_9313 = 3'h3 == state ? _GEN_5944 : _GEN_8754; // @[DCache.scala 260:17]
  wire  _GEN_9314 = 3'h3 == state ? _GEN_5945 : _GEN_8755; // @[DCache.scala 260:17]
  wire  _GEN_9315 = 3'h3 == state ? _GEN_5946 : _GEN_8756; // @[DCache.scala 260:17]
  wire  _GEN_9316 = 3'h3 == state ? _GEN_5947 : _GEN_8757; // @[DCache.scala 260:17]
  wire  _GEN_9317 = 3'h3 == state ? _GEN_5948 : _GEN_8758; // @[DCache.scala 260:17]
  wire  _GEN_9318 = 3'h3 == state ? _GEN_5949 : _GEN_8759; // @[DCache.scala 260:17]
  wire  _GEN_9319 = 3'h3 == state ? _GEN_5950 : _GEN_8760; // @[DCache.scala 260:17]
  wire  _GEN_9320 = 3'h3 == state ? _GEN_5951 : _GEN_8761; // @[DCache.scala 260:17]
  wire  _GEN_9321 = 3'h3 == state ? _GEN_5952 : _GEN_8762; // @[DCache.scala 260:17]
  wire  _GEN_9322 = 3'h3 == state ? _GEN_5953 : _GEN_8763; // @[DCache.scala 260:17]
  wire  _GEN_9323 = 3'h3 == state ? _GEN_5954 : _GEN_8764; // @[DCache.scala 260:17]
  wire  _GEN_9324 = 3'h3 == state ? _GEN_5955 : _GEN_8765; // @[DCache.scala 260:17]
  wire  _GEN_9325 = 3'h3 == state ? _GEN_5956 : _GEN_8766; // @[DCache.scala 260:17]
  wire  _GEN_9326 = 3'h3 == state ? _GEN_5957 : _GEN_8767; // @[DCache.scala 260:17]
  wire  _GEN_9327 = 3'h3 == state ? _GEN_5958 : _GEN_8768; // @[DCache.scala 260:17]
  wire  _GEN_9328 = 3'h3 == state ? _GEN_5959 : _GEN_8769; // @[DCache.scala 260:17]
  wire  _GEN_9329 = 3'h3 == state ? _GEN_5960 : _GEN_8770; // @[DCache.scala 260:17]
  wire  _GEN_9330 = 3'h3 == state ? _GEN_5961 : _GEN_8771; // @[DCache.scala 260:17]
  wire  _GEN_9331 = 3'h3 == state ? _GEN_5962 : _GEN_8772; // @[DCache.scala 260:17]
  wire  _GEN_9332 = 3'h3 == state ? _GEN_5963 : _GEN_8773; // @[DCache.scala 260:17]
  wire  _GEN_9333 = 3'h3 == state ? _GEN_5964 : _GEN_8774; // @[DCache.scala 260:17]
  wire  _GEN_9334 = 3'h3 == state ? _GEN_5965 : _GEN_8775; // @[DCache.scala 260:17]
  wire  _GEN_9335 = 3'h3 == state ? _GEN_5966 : _GEN_8776; // @[DCache.scala 260:17]
  wire  _GEN_9336 = 3'h3 == state ? _GEN_5967 : _GEN_8777; // @[DCache.scala 260:17]
  wire  _GEN_9337 = 3'h3 == state ? _GEN_5968 : _GEN_8778; // @[DCache.scala 260:17]
  wire  _GEN_9338 = 3'h3 == state ? _GEN_5969 : _GEN_8779; // @[DCache.scala 260:17]
  wire  _GEN_9339 = 3'h3 == state ? _GEN_5970 : _GEN_8780; // @[DCache.scala 260:17]
  wire  _GEN_9340 = 3'h3 == state ? _GEN_5971 : _GEN_8781; // @[DCache.scala 260:17]
  wire  _GEN_9341 = 3'h3 == state ? _GEN_5972 : _GEN_8782; // @[DCache.scala 260:17]
  wire  _GEN_9342 = 3'h3 == state ? _GEN_5973 : _GEN_8783; // @[DCache.scala 260:17]
  wire  _GEN_9343 = 3'h3 == state ? _GEN_5974 : _GEN_8784; // @[DCache.scala 260:17]
  wire  _GEN_9344 = 3'h3 == state ? _GEN_5975 : _GEN_8785; // @[DCache.scala 260:17]
  wire  _GEN_9345 = 3'h3 == state ? _GEN_5976 : _GEN_8786; // @[DCache.scala 260:17]
  wire  _GEN_9346 = 3'h3 == state ? _GEN_5977 : _GEN_8787; // @[DCache.scala 260:17]
  wire  _GEN_9347 = 3'h3 == state ? _GEN_5978 : _GEN_8788; // @[DCache.scala 260:17]
  wire  _GEN_9348 = 3'h3 == state ? _GEN_5979 : _GEN_8789; // @[DCache.scala 260:17]
  wire  _GEN_9349 = 3'h3 == state ? _GEN_5980 : _GEN_8790; // @[DCache.scala 260:17]
  wire  _GEN_9350 = 3'h3 == state ? _GEN_5981 : _GEN_8791; // @[DCache.scala 260:17]
  wire  _GEN_9351 = 3'h3 == state ? _GEN_5982 : _GEN_8792; // @[DCache.scala 260:17]
  wire  _GEN_9352 = 3'h3 == state ? _GEN_5983 : _GEN_8793; // @[DCache.scala 260:17]
  wire  _GEN_9353 = 3'h3 == state ? _GEN_5984 : _GEN_8794; // @[DCache.scala 260:17]
  wire  _GEN_9354 = 3'h3 == state ? _GEN_5985 : _GEN_8795; // @[DCache.scala 260:17]
  wire  _GEN_9355 = 3'h3 == state ? _GEN_5986 : _GEN_8796; // @[DCache.scala 260:17]
  wire  _GEN_9356 = 3'h3 == state ? _GEN_5987 : _GEN_8797; // @[DCache.scala 260:17]
  wire  _GEN_9357 = 3'h3 == state ? _GEN_5988 : _GEN_8798; // @[DCache.scala 260:17]
  wire  _GEN_9358 = 3'h3 == state ? _GEN_5989 : _GEN_8799; // @[DCache.scala 260:17]
  wire  _GEN_9359 = 3'h3 == state ? _GEN_5990 : _GEN_8800; // @[DCache.scala 260:17]
  wire  _GEN_9360 = 3'h3 == state ? _GEN_5991 : _GEN_8801; // @[DCache.scala 260:17]
  wire  _GEN_9361 = 3'h3 == state ? _GEN_5992 : _GEN_8802; // @[DCache.scala 260:17]
  wire  _GEN_9362 = 3'h3 == state ? _GEN_5993 : _GEN_8803; // @[DCache.scala 260:17]
  wire  _GEN_9363 = 3'h3 == state ? _GEN_5994 : _GEN_8804; // @[DCache.scala 260:17]
  wire  _GEN_9364 = 3'h3 == state ? _GEN_5995 : _GEN_8805; // @[DCache.scala 260:17]
  wire  _GEN_9365 = 3'h3 == state ? _GEN_5996 : _GEN_8806; // @[DCache.scala 260:17]
  wire  _GEN_9366 = 3'h3 == state ? _GEN_5997 : _GEN_8807; // @[DCache.scala 260:17]
  wire  _GEN_9367 = 3'h3 == state ? _GEN_5998 : _GEN_8808; // @[DCache.scala 260:17]
  wire  _GEN_9368 = 3'h3 == state ? _GEN_5999 : _GEN_8809; // @[DCache.scala 260:17]
  wire  _GEN_9369 = 3'h3 == state ? _GEN_6000 : _GEN_8810; // @[DCache.scala 260:17]
  wire  _GEN_9370 = 3'h3 == state ? _GEN_6001 : _GEN_8811; // @[DCache.scala 260:17]
  wire  _GEN_9371 = 3'h3 == state ? _GEN_6002 : _GEN_8812; // @[DCache.scala 260:17]
  wire  _GEN_9372 = 3'h3 == state ? _GEN_6003 : _GEN_8813; // @[DCache.scala 260:17]
  wire  _GEN_9373 = 3'h3 == state ? _GEN_6004 : _GEN_8814; // @[DCache.scala 260:17]
  wire  _GEN_9374 = 3'h3 == state ? _GEN_6005 : _GEN_8815; // @[DCache.scala 260:17]
  wire  _GEN_9375 = 3'h3 == state ? _GEN_6006 : _GEN_8816; // @[DCache.scala 260:17]
  wire  _GEN_9376 = 3'h3 == state ? _GEN_6007 : _GEN_8817; // @[DCache.scala 260:17]
  wire  _GEN_9377 = 3'h3 == state ? _GEN_6008 : _GEN_8818; // @[DCache.scala 260:17]
  wire  _GEN_9378 = 3'h3 == state ? _GEN_6009 : _GEN_8819; // @[DCache.scala 260:17]
  wire  _GEN_9379 = 3'h3 == state ? _GEN_6010 : _GEN_8820; // @[DCache.scala 260:17]
  wire  _GEN_9380 = 3'h3 == state ? _GEN_6011 : _GEN_8821; // @[DCache.scala 260:17]
  wire  _GEN_9381 = 3'h3 == state ? _GEN_6012 : _GEN_8822; // @[DCache.scala 260:17]
  wire  _GEN_9382 = 3'h3 == state ? _GEN_6013 : _GEN_8823; // @[DCache.scala 260:17]
  wire  _GEN_9383 = 3'h3 == state ? _GEN_6014 : _GEN_8824; // @[DCache.scala 260:17]
  wire  _GEN_9384 = 3'h3 == state ? _GEN_6015 : _GEN_8825; // @[DCache.scala 260:17]
  wire  _GEN_9385 = 3'h3 == state ? _GEN_6016 : _GEN_8826; // @[DCache.scala 260:17]
  wire  _GEN_9386 = 3'h3 == state ? _GEN_6017 : _GEN_8827; // @[DCache.scala 260:17]
  wire  _GEN_9387 = 3'h3 == state ? _GEN_6018 : _GEN_8828; // @[DCache.scala 260:17]
  wire  _GEN_9388 = 3'h3 == state ? _GEN_6019 : _GEN_8829; // @[DCache.scala 260:17]
  wire  _GEN_9389 = 3'h3 == state ? _GEN_6020 : _GEN_8830; // @[DCache.scala 260:17]
  wire  _GEN_9390 = 3'h3 == state ? _GEN_6021 : _GEN_8831; // @[DCache.scala 260:17]
  wire  _GEN_9391 = 3'h3 == state ? _GEN_6022 : _GEN_8832; // @[DCache.scala 260:17]
  wire  _GEN_9392 = 3'h3 == state ? _GEN_6023 : _GEN_8833; // @[DCache.scala 260:17]
  wire  _GEN_9393 = 3'h3 == state ? _GEN_6024 : _GEN_8834; // @[DCache.scala 260:17]
  wire  _GEN_9394 = 3'h3 == state ? _GEN_6025 : _GEN_8835; // @[DCache.scala 260:17]
  wire  _GEN_9395 = 3'h3 == state ? _GEN_6026 : _GEN_8836; // @[DCache.scala 260:17]
  wire  _GEN_9396 = 3'h3 == state ? _GEN_6027 : _GEN_8837; // @[DCache.scala 260:17]
  wire  _GEN_9397 = 3'h3 == state ? _GEN_6028 : _GEN_8838; // @[DCache.scala 260:17]
  wire  _GEN_9398 = 3'h3 == state ? _GEN_6029 : _GEN_8839; // @[DCache.scala 260:17]
  wire  _GEN_9399 = 3'h3 == state ? _GEN_6030 : _GEN_8840; // @[DCache.scala 260:17]
  wire  _GEN_9400 = 3'h3 == state ? _GEN_6031 : _GEN_8841; // @[DCache.scala 260:17]
  wire  _GEN_9401 = 3'h3 == state ? _GEN_6032 : _GEN_8842; // @[DCache.scala 260:17]
  wire  _GEN_9402 = 3'h3 == state ? _GEN_6033 : _GEN_8843; // @[DCache.scala 260:17]
  wire  _GEN_9403 = 3'h3 == state ? _GEN_6034 : _GEN_8844; // @[DCache.scala 260:17]
  wire  _GEN_9404 = 3'h3 == state ? _GEN_6035 : fence_working; // @[DCache.scala 260:17 97:40]
  wire  _GEN_9405 = 3'h3 == state ? _GEN_6036 : _GEN_8858; // @[DCache.scala 260:17]
  wire [2:0] _GEN_9406 = 3'h3 == state ? _GEN_6037 : _GEN_9116; // @[DCache.scala 260:17]
  wire  _GEN_9407 = 3'h3 == state ? replace_writeback : _GEN_8845; // @[DCache.scala 260:17 101:40]
  wire [31:0] _GEN_9408 = 3'h3 == state ? ar_addr : _GEN_8846; // @[DCache.scala 260:17 199:24]
  wire [7:0] _GEN_9409 = 3'h3 == state ? ar_len : _GEN_8847; // @[DCache.scala 260:17 199:24]
  wire [2:0] _GEN_9410 = 3'h3 == state ? ar_size : _GEN_8848; // @[DCache.scala 260:17 199:24]
  wire  _GEN_9411 = 3'h3 == state ? arvalid : _GEN_8849; // @[DCache.scala 260:17 200:24]
  wire  _GEN_9412 = 3'h3 == state ? rready : _GEN_8850; // @[DCache.scala 260:17 203:23]
  wire  _GEN_9413 = 3'h3 == state ? ar_handshake : _GEN_8851; // @[DCache.scala 260:17 99:40]
  wire [3:0] _GEN_9414 = 3'h3 == state ? bram_replace_wea_0 : _GEN_8852; // @[DCache.scala 260:17 73:33]
  wire [3:0] _GEN_9415 = 3'h3 == state ? bram_replace_wea_1 : _GEN_8853; // @[DCache.scala 260:17 73:33]
  wire  _GEN_9416 = 3'h3 == state ? tag_wstrb_0 : _GEN_8854; // @[DCache.scala 260:17 72:33]
  wire  _GEN_9417 = 3'h3 == state ? tag_wstrb_1 : _GEN_8855; // @[DCache.scala 260:17 72:33]
  wire [19:0] _GEN_9418 = 3'h3 == state ? tag_wdata : _GEN_8856; // @[DCache.scala 260:17 77:26]
  wire [9:0] _GEN_9419 = 3'h3 == state ? bram_replace_write_addr : _GEN_8857; // @[DCache.scala 260:17 92:40]
  wire  _GEN_9420 = 3'h3 == state ? valid_0_0 : _GEN_8859; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9421 = 3'h3 == state ? valid_0_1 : _GEN_8860; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9422 = 3'h3 == state ? valid_1_0 : _GEN_8861; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9423 = 3'h3 == state ? valid_1_1 : _GEN_8862; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9424 = 3'h3 == state ? valid_2_0 : _GEN_8863; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9425 = 3'h3 == state ? valid_2_1 : _GEN_8864; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9426 = 3'h3 == state ? valid_3_0 : _GEN_8865; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9427 = 3'h3 == state ? valid_3_1 : _GEN_8866; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9428 = 3'h3 == state ? valid_4_0 : _GEN_8867; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9429 = 3'h3 == state ? valid_4_1 : _GEN_8868; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9430 = 3'h3 == state ? valid_5_0 : _GEN_8869; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9431 = 3'h3 == state ? valid_5_1 : _GEN_8870; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9432 = 3'h3 == state ? valid_6_0 : _GEN_8871; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9433 = 3'h3 == state ? valid_6_1 : _GEN_8872; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9434 = 3'h3 == state ? valid_7_0 : _GEN_8873; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9435 = 3'h3 == state ? valid_7_1 : _GEN_8874; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9436 = 3'h3 == state ? valid_8_0 : _GEN_8875; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9437 = 3'h3 == state ? valid_8_1 : _GEN_8876; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9438 = 3'h3 == state ? valid_9_0 : _GEN_8877; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9439 = 3'h3 == state ? valid_9_1 : _GEN_8878; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9440 = 3'h3 == state ? valid_10_0 : _GEN_8879; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9441 = 3'h3 == state ? valid_10_1 : _GEN_8880; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9442 = 3'h3 == state ? valid_11_0 : _GEN_8881; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9443 = 3'h3 == state ? valid_11_1 : _GEN_8882; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9444 = 3'h3 == state ? valid_12_0 : _GEN_8883; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9445 = 3'h3 == state ? valid_12_1 : _GEN_8884; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9446 = 3'h3 == state ? valid_13_0 : _GEN_8885; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9447 = 3'h3 == state ? valid_13_1 : _GEN_8886; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9448 = 3'h3 == state ? valid_14_0 : _GEN_8887; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9449 = 3'h3 == state ? valid_14_1 : _GEN_8888; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9450 = 3'h3 == state ? valid_15_0 : _GEN_8889; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9451 = 3'h3 == state ? valid_15_1 : _GEN_8890; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9452 = 3'h3 == state ? valid_16_0 : _GEN_8891; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9453 = 3'h3 == state ? valid_16_1 : _GEN_8892; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9454 = 3'h3 == state ? valid_17_0 : _GEN_8893; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9455 = 3'h3 == state ? valid_17_1 : _GEN_8894; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9456 = 3'h3 == state ? valid_18_0 : _GEN_8895; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9457 = 3'h3 == state ? valid_18_1 : _GEN_8896; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9458 = 3'h3 == state ? valid_19_0 : _GEN_8897; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9459 = 3'h3 == state ? valid_19_1 : _GEN_8898; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9460 = 3'h3 == state ? valid_20_0 : _GEN_8899; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9461 = 3'h3 == state ? valid_20_1 : _GEN_8900; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9462 = 3'h3 == state ? valid_21_0 : _GEN_8901; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9463 = 3'h3 == state ? valid_21_1 : _GEN_8902; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9464 = 3'h3 == state ? valid_22_0 : _GEN_8903; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9465 = 3'h3 == state ? valid_22_1 : _GEN_8904; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9466 = 3'h3 == state ? valid_23_0 : _GEN_8905; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9467 = 3'h3 == state ? valid_23_1 : _GEN_8906; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9468 = 3'h3 == state ? valid_24_0 : _GEN_8907; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9469 = 3'h3 == state ? valid_24_1 : _GEN_8908; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9470 = 3'h3 == state ? valid_25_0 : _GEN_8909; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9471 = 3'h3 == state ? valid_25_1 : _GEN_8910; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9472 = 3'h3 == state ? valid_26_0 : _GEN_8911; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9473 = 3'h3 == state ? valid_26_1 : _GEN_8912; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9474 = 3'h3 == state ? valid_27_0 : _GEN_8913; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9475 = 3'h3 == state ? valid_27_1 : _GEN_8914; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9476 = 3'h3 == state ? valid_28_0 : _GEN_8915; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9477 = 3'h3 == state ? valid_28_1 : _GEN_8916; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9478 = 3'h3 == state ? valid_29_0 : _GEN_8917; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9479 = 3'h3 == state ? valid_29_1 : _GEN_8918; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9480 = 3'h3 == state ? valid_30_0 : _GEN_8919; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9481 = 3'h3 == state ? valid_30_1 : _GEN_8920; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9482 = 3'h3 == state ? valid_31_0 : _GEN_8921; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9483 = 3'h3 == state ? valid_31_1 : _GEN_8922; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9484 = 3'h3 == state ? valid_32_0 : _GEN_8923; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9485 = 3'h3 == state ? valid_32_1 : _GEN_8924; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9486 = 3'h3 == state ? valid_33_0 : _GEN_8925; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9487 = 3'h3 == state ? valid_33_1 : _GEN_8926; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9488 = 3'h3 == state ? valid_34_0 : _GEN_8927; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9489 = 3'h3 == state ? valid_34_1 : _GEN_8928; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9490 = 3'h3 == state ? valid_35_0 : _GEN_8929; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9491 = 3'h3 == state ? valid_35_1 : _GEN_8930; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9492 = 3'h3 == state ? valid_36_0 : _GEN_8931; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9493 = 3'h3 == state ? valid_36_1 : _GEN_8932; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9494 = 3'h3 == state ? valid_37_0 : _GEN_8933; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9495 = 3'h3 == state ? valid_37_1 : _GEN_8934; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9496 = 3'h3 == state ? valid_38_0 : _GEN_8935; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9497 = 3'h3 == state ? valid_38_1 : _GEN_8936; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9498 = 3'h3 == state ? valid_39_0 : _GEN_8937; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9499 = 3'h3 == state ? valid_39_1 : _GEN_8938; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9500 = 3'h3 == state ? valid_40_0 : _GEN_8939; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9501 = 3'h3 == state ? valid_40_1 : _GEN_8940; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9502 = 3'h3 == state ? valid_41_0 : _GEN_8941; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9503 = 3'h3 == state ? valid_41_1 : _GEN_8942; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9504 = 3'h3 == state ? valid_42_0 : _GEN_8943; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9505 = 3'h3 == state ? valid_42_1 : _GEN_8944; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9506 = 3'h3 == state ? valid_43_0 : _GEN_8945; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9507 = 3'h3 == state ? valid_43_1 : _GEN_8946; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9508 = 3'h3 == state ? valid_44_0 : _GEN_8947; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9509 = 3'h3 == state ? valid_44_1 : _GEN_8948; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9510 = 3'h3 == state ? valid_45_0 : _GEN_8949; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9511 = 3'h3 == state ? valid_45_1 : _GEN_8950; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9512 = 3'h3 == state ? valid_46_0 : _GEN_8951; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9513 = 3'h3 == state ? valid_46_1 : _GEN_8952; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9514 = 3'h3 == state ? valid_47_0 : _GEN_8953; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9515 = 3'h3 == state ? valid_47_1 : _GEN_8954; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9516 = 3'h3 == state ? valid_48_0 : _GEN_8955; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9517 = 3'h3 == state ? valid_48_1 : _GEN_8956; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9518 = 3'h3 == state ? valid_49_0 : _GEN_8957; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9519 = 3'h3 == state ? valid_49_1 : _GEN_8958; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9520 = 3'h3 == state ? valid_50_0 : _GEN_8959; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9521 = 3'h3 == state ? valid_50_1 : _GEN_8960; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9522 = 3'h3 == state ? valid_51_0 : _GEN_8961; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9523 = 3'h3 == state ? valid_51_1 : _GEN_8962; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9524 = 3'h3 == state ? valid_52_0 : _GEN_8963; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9525 = 3'h3 == state ? valid_52_1 : _GEN_8964; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9526 = 3'h3 == state ? valid_53_0 : _GEN_8965; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9527 = 3'h3 == state ? valid_53_1 : _GEN_8966; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9528 = 3'h3 == state ? valid_54_0 : _GEN_8967; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9529 = 3'h3 == state ? valid_54_1 : _GEN_8968; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9530 = 3'h3 == state ? valid_55_0 : _GEN_8969; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9531 = 3'h3 == state ? valid_55_1 : _GEN_8970; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9532 = 3'h3 == state ? valid_56_0 : _GEN_8971; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9533 = 3'h3 == state ? valid_56_1 : _GEN_8972; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9534 = 3'h3 == state ? valid_57_0 : _GEN_8973; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9535 = 3'h3 == state ? valid_57_1 : _GEN_8974; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9536 = 3'h3 == state ? valid_58_0 : _GEN_8975; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9537 = 3'h3 == state ? valid_58_1 : _GEN_8976; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9538 = 3'h3 == state ? valid_59_0 : _GEN_8977; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9539 = 3'h3 == state ? valid_59_1 : _GEN_8978; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9540 = 3'h3 == state ? valid_60_0 : _GEN_8979; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9541 = 3'h3 == state ? valid_60_1 : _GEN_8980; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9542 = 3'h3 == state ? valid_61_0 : _GEN_8981; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9543 = 3'h3 == state ? valid_61_1 : _GEN_8982; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9544 = 3'h3 == state ? valid_62_0 : _GEN_8983; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9545 = 3'h3 == state ? valid_62_1 : _GEN_8984; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9546 = 3'h3 == state ? valid_63_0 : _GEN_8985; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9547 = 3'h3 == state ? valid_63_1 : _GEN_8986; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9548 = 3'h3 == state ? valid_64_0 : _GEN_8987; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9549 = 3'h3 == state ? valid_64_1 : _GEN_8988; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9550 = 3'h3 == state ? valid_65_0 : _GEN_8989; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9551 = 3'h3 == state ? valid_65_1 : _GEN_8990; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9552 = 3'h3 == state ? valid_66_0 : _GEN_8991; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9553 = 3'h3 == state ? valid_66_1 : _GEN_8992; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9554 = 3'h3 == state ? valid_67_0 : _GEN_8993; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9555 = 3'h3 == state ? valid_67_1 : _GEN_8994; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9556 = 3'h3 == state ? valid_68_0 : _GEN_8995; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9557 = 3'h3 == state ? valid_68_1 : _GEN_8996; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9558 = 3'h3 == state ? valid_69_0 : _GEN_8997; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9559 = 3'h3 == state ? valid_69_1 : _GEN_8998; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9560 = 3'h3 == state ? valid_70_0 : _GEN_8999; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9561 = 3'h3 == state ? valid_70_1 : _GEN_9000; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9562 = 3'h3 == state ? valid_71_0 : _GEN_9001; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9563 = 3'h3 == state ? valid_71_1 : _GEN_9002; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9564 = 3'h3 == state ? valid_72_0 : _GEN_9003; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9565 = 3'h3 == state ? valid_72_1 : _GEN_9004; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9566 = 3'h3 == state ? valid_73_0 : _GEN_9005; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9567 = 3'h3 == state ? valid_73_1 : _GEN_9006; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9568 = 3'h3 == state ? valid_74_0 : _GEN_9007; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9569 = 3'h3 == state ? valid_74_1 : _GEN_9008; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9570 = 3'h3 == state ? valid_75_0 : _GEN_9009; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9571 = 3'h3 == state ? valid_75_1 : _GEN_9010; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9572 = 3'h3 == state ? valid_76_0 : _GEN_9011; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9573 = 3'h3 == state ? valid_76_1 : _GEN_9012; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9574 = 3'h3 == state ? valid_77_0 : _GEN_9013; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9575 = 3'h3 == state ? valid_77_1 : _GEN_9014; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9576 = 3'h3 == state ? valid_78_0 : _GEN_9015; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9577 = 3'h3 == state ? valid_78_1 : _GEN_9016; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9578 = 3'h3 == state ? valid_79_0 : _GEN_9017; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9579 = 3'h3 == state ? valid_79_1 : _GEN_9018; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9580 = 3'h3 == state ? valid_80_0 : _GEN_9019; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9581 = 3'h3 == state ? valid_80_1 : _GEN_9020; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9582 = 3'h3 == state ? valid_81_0 : _GEN_9021; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9583 = 3'h3 == state ? valid_81_1 : _GEN_9022; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9584 = 3'h3 == state ? valid_82_0 : _GEN_9023; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9585 = 3'h3 == state ? valid_82_1 : _GEN_9024; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9586 = 3'h3 == state ? valid_83_0 : _GEN_9025; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9587 = 3'h3 == state ? valid_83_1 : _GEN_9026; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9588 = 3'h3 == state ? valid_84_0 : _GEN_9027; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9589 = 3'h3 == state ? valid_84_1 : _GEN_9028; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9590 = 3'h3 == state ? valid_85_0 : _GEN_9029; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9591 = 3'h3 == state ? valid_85_1 : _GEN_9030; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9592 = 3'h3 == state ? valid_86_0 : _GEN_9031; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9593 = 3'h3 == state ? valid_86_1 : _GEN_9032; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9594 = 3'h3 == state ? valid_87_0 : _GEN_9033; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9595 = 3'h3 == state ? valid_87_1 : _GEN_9034; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9596 = 3'h3 == state ? valid_88_0 : _GEN_9035; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9597 = 3'h3 == state ? valid_88_1 : _GEN_9036; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9598 = 3'h3 == state ? valid_89_0 : _GEN_9037; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9599 = 3'h3 == state ? valid_89_1 : _GEN_9038; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9600 = 3'h3 == state ? valid_90_0 : _GEN_9039; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9601 = 3'h3 == state ? valid_90_1 : _GEN_9040; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9602 = 3'h3 == state ? valid_91_0 : _GEN_9041; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9603 = 3'h3 == state ? valid_91_1 : _GEN_9042; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9604 = 3'h3 == state ? valid_92_0 : _GEN_9043; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9605 = 3'h3 == state ? valid_92_1 : _GEN_9044; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9606 = 3'h3 == state ? valid_93_0 : _GEN_9045; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9607 = 3'h3 == state ? valid_93_1 : _GEN_9046; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9608 = 3'h3 == state ? valid_94_0 : _GEN_9047; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9609 = 3'h3 == state ? valid_94_1 : _GEN_9048; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9610 = 3'h3 == state ? valid_95_0 : _GEN_9049; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9611 = 3'h3 == state ? valid_95_1 : _GEN_9050; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9612 = 3'h3 == state ? valid_96_0 : _GEN_9051; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9613 = 3'h3 == state ? valid_96_1 : _GEN_9052; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9614 = 3'h3 == state ? valid_97_0 : _GEN_9053; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9615 = 3'h3 == state ? valid_97_1 : _GEN_9054; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9616 = 3'h3 == state ? valid_98_0 : _GEN_9055; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9617 = 3'h3 == state ? valid_98_1 : _GEN_9056; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9618 = 3'h3 == state ? valid_99_0 : _GEN_9057; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9619 = 3'h3 == state ? valid_99_1 : _GEN_9058; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9620 = 3'h3 == state ? valid_100_0 : _GEN_9059; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9621 = 3'h3 == state ? valid_100_1 : _GEN_9060; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9622 = 3'h3 == state ? valid_101_0 : _GEN_9061; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9623 = 3'h3 == state ? valid_101_1 : _GEN_9062; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9624 = 3'h3 == state ? valid_102_0 : _GEN_9063; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9625 = 3'h3 == state ? valid_102_1 : _GEN_9064; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9626 = 3'h3 == state ? valid_103_0 : _GEN_9065; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9627 = 3'h3 == state ? valid_103_1 : _GEN_9066; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9628 = 3'h3 == state ? valid_104_0 : _GEN_9067; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9629 = 3'h3 == state ? valid_104_1 : _GEN_9068; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9630 = 3'h3 == state ? valid_105_0 : _GEN_9069; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9631 = 3'h3 == state ? valid_105_1 : _GEN_9070; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9632 = 3'h3 == state ? valid_106_0 : _GEN_9071; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9633 = 3'h3 == state ? valid_106_1 : _GEN_9072; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9634 = 3'h3 == state ? valid_107_0 : _GEN_9073; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9635 = 3'h3 == state ? valid_107_1 : _GEN_9074; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9636 = 3'h3 == state ? valid_108_0 : _GEN_9075; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9637 = 3'h3 == state ? valid_108_1 : _GEN_9076; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9638 = 3'h3 == state ? valid_109_0 : _GEN_9077; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9639 = 3'h3 == state ? valid_109_1 : _GEN_9078; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9640 = 3'h3 == state ? valid_110_0 : _GEN_9079; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9641 = 3'h3 == state ? valid_110_1 : _GEN_9080; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9642 = 3'h3 == state ? valid_111_0 : _GEN_9081; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9643 = 3'h3 == state ? valid_111_1 : _GEN_9082; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9644 = 3'h3 == state ? valid_112_0 : _GEN_9083; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9645 = 3'h3 == state ? valid_112_1 : _GEN_9084; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9646 = 3'h3 == state ? valid_113_0 : _GEN_9085; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9647 = 3'h3 == state ? valid_113_1 : _GEN_9086; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9648 = 3'h3 == state ? valid_114_0 : _GEN_9087; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9649 = 3'h3 == state ? valid_114_1 : _GEN_9088; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9650 = 3'h3 == state ? valid_115_0 : _GEN_9089; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9651 = 3'h3 == state ? valid_115_1 : _GEN_9090; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9652 = 3'h3 == state ? valid_116_0 : _GEN_9091; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9653 = 3'h3 == state ? valid_116_1 : _GEN_9092; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9654 = 3'h3 == state ? valid_117_0 : _GEN_9093; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9655 = 3'h3 == state ? valid_117_1 : _GEN_9094; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9656 = 3'h3 == state ? valid_118_0 : _GEN_9095; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9657 = 3'h3 == state ? valid_118_1 : _GEN_9096; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9658 = 3'h3 == state ? valid_119_0 : _GEN_9097; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9659 = 3'h3 == state ? valid_119_1 : _GEN_9098; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9660 = 3'h3 == state ? valid_120_0 : _GEN_9099; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9661 = 3'h3 == state ? valid_120_1 : _GEN_9100; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9662 = 3'h3 == state ? valid_121_0 : _GEN_9101; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9663 = 3'h3 == state ? valid_121_1 : _GEN_9102; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9664 = 3'h3 == state ? valid_122_0 : _GEN_9103; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9665 = 3'h3 == state ? valid_122_1 : _GEN_9104; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9666 = 3'h3 == state ? valid_123_0 : _GEN_9105; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9667 = 3'h3 == state ? valid_123_1 : _GEN_9106; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9668 = 3'h3 == state ? valid_124_0 : _GEN_9107; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9669 = 3'h3 == state ? valid_124_1 : _GEN_9108; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9670 = 3'h3 == state ? valid_125_0 : _GEN_9109; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9671 = 3'h3 == state ? valid_125_1 : _GEN_9110; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9672 = 3'h3 == state ? valid_126_0 : _GEN_9111; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9673 = 3'h3 == state ? valid_126_1 : _GEN_9112; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9674 = 3'h3 == state ? valid_127_0 : _GEN_9113; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9675 = 3'h3 == state ? valid_127_1 : _GEN_9114; // @[DCache.scala 260:17 68:22]
  wire  _GEN_9676 = 3'h3 == state ? replace_working : _GEN_9115; // @[DCache.scala 260:17 98:40]
  wire  _GEN_9677 = 3'h3 == state ? data_tlb_invalid : _GEN_9117; // @[DCache.scala 260:17 250:25]
  wire  _GEN_9678 = 3'h3 == state ? data_tlb_refill : _GEN_9118; // @[DCache.scala 260:17 250:25]
  wire  _GEN_9679 = 3'h3 == state ? data_tlb_mod : _GEN_9119; // @[DCache.scala 260:17 250:25]
  wire [19:0] _GEN_10809 = 3'h0 == state ? _GEN_4491 : {{1'd0}, tlb2_vpn}; // @[DCache.scala 260:17 245:21]
  wire [19:0] _GEN_15206 = reset ? 20'h0 : _GEN_10809; // @[DCache.scala 245:{21,21}]
  Queue write_buffer ( // @[DCache.scala 82:28]
    .clock(write_buffer_clock),
    .reset(write_buffer_reset),
    .io_enq_ready(write_buffer_io_enq_ready),
    .io_enq_valid(write_buffer_io_enq_valid),
    .io_enq_bits_data(write_buffer_io_enq_bits_data),
    .io_enq_bits_addr(write_buffer_io_enq_bits_addr),
    .io_enq_bits_strb(write_buffer_io_enq_bits_strb),
    .io_enq_bits_size(write_buffer_io_enq_bits_size),
    .io_deq_ready(write_buffer_io_deq_ready),
    .io_deq_valid(write_buffer_io_deq_valid),
    .io_deq_bits_data(write_buffer_io_deq_bits_data),
    .io_deq_bits_addr(write_buffer_io_deq_bits_addr),
    .io_deq_bits_strb(write_buffer_io_deq_bits_strb),
    .io_deq_bits_size(write_buffer_io_deq_bits_size)
  );
  SimpleDualPortRam_8 bank_ram ( // @[DCache.scala 153:26]
    .clock(bank_ram_clock),
    .reset(bank_ram_reset),
    .io_raddr(bank_ram_io_raddr),
    .io_rdata(bank_ram_io_rdata),
    .io_waddr(bank_ram_io_waddr),
    .io_wen(bank_ram_io_wen),
    .io_wstrb(bank_ram_io_wstrb),
    .io_wdata(bank_ram_io_wdata)
  );
  SimpleDualPortRam_9 tag_ram ( // @[DCache.scala 163:25]
    .clock(tag_ram_clock),
    .reset(tag_ram_reset),
    .io_raddr(tag_ram_io_raddr),
    .io_rdata(tag_ram_io_rdata),
    .io_waddr(tag_ram_io_waddr),
    .io_wen(tag_ram_io_wen),
    .io_wstrb(tag_ram_io_wstrb),
    .io_wdata(tag_ram_io_wdata)
  );
  SimpleDualPortRam_8 bank_ram_1 ( // @[DCache.scala 153:26]
    .clock(bank_ram_1_clock),
    .reset(bank_ram_1_reset),
    .io_raddr(bank_ram_1_io_raddr),
    .io_rdata(bank_ram_1_io_rdata),
    .io_waddr(bank_ram_1_io_waddr),
    .io_wen(bank_ram_1_io_wen),
    .io_wstrb(bank_ram_1_io_wstrb),
    .io_wdata(bank_ram_1_io_wdata)
  );
  SimpleDualPortRam_9 tag_ram_1 ( // @[DCache.scala 163:25]
    .clock(tag_ram_1_clock),
    .reset(tag_ram_1_reset),
    .io_raddr(tag_ram_1_io_raddr),
    .io_rdata(tag_ram_1_io_rdata),
    .io_waddr(tag_ram_1_io_waddr),
    .io_wen(tag_ram_1_io_wen),
    .io_wstrb(tag_ram_1_io_wstrb),
    .io_wdata(tag_ram_1_io_wdata)
  );
  assign io_cpu_dstall = _io_cpu_dstall_T ? _io_cpu_dstall_T_4 : _bram_addr_choose_T_1; // @[DCache.scala 135:23]
  assign io_cpu_M_rdata = state == 3'h5 ? saved_rdata : _GEN_1; // @[DCache.scala 149:24]
  assign io_cpu_tlb_vpn2 = tlb2_vpn; // @[DCache.scala 248:19]
  assign io_cpu_data_tlb_refill = data_tlb_refill; // @[DCache.scala 256:27]
  assign io_cpu_data_tlb_invalid = data_tlb_invalid; // @[DCache.scala 257:27]
  assign io_cpu_data_tlb_mod = data_tlb_mod; // @[DCache.scala 258:27]
  assign io_axi_ar_valid = arvalid; // @[DCache.scala 202:19]
  assign io_axi_ar_bits_addr = ar_addr; // @[DCache.scala 201:18]
  assign io_axi_ar_bits_len = ar_len; // @[DCache.scala 201:18]
  assign io_axi_ar_bits_size = ar_size; // @[DCache.scala 201:18]
  assign io_axi_r_ready = rready; // @[DCache.scala 204:18]
  assign io_axi_aw_valid = awvalid; // @[DCache.scala 208:19]
  assign io_axi_aw_bits_addr = aw_addr; // @[DCache.scala 207:18]
  assign io_axi_aw_bits_len = aw_len; // @[DCache.scala 207:18]
  assign io_axi_aw_bits_size = aw_size; // @[DCache.scala 207:18]
  assign io_axi_w_valid = wvalid; // @[DCache.scala 212:18]
  assign io_axi_w_bits_data = w_data; // @[DCache.scala 211:17]
  assign io_axi_w_bits_strb = w_strb; // @[DCache.scala 211:17]
  assign io_axi_w_bits_last = w_last; // @[DCache.scala 211:17]
  assign io_axi_b_ready = 1'h1; // @[DCache.scala 214:18]
  assign write_buffer_clock = clock;
  assign write_buffer_reset = reset;
  assign write_buffer_io_enq_valid = 3'h0 == state & _GEN_4492; // @[DCache.scala 260:17 83:29]
  assign write_buffer_io_enq_bits_data = 3'h0 == state ? _GEN_4496 : 32'h0; // @[DCache.scala 260:17 84:29]
  assign write_buffer_io_enq_bits_addr = 3'h0 == state ? _GEN_4493 : 32'h0; // @[DCache.scala 260:17 84:29]
  assign write_buffer_io_enq_bits_strb = 3'h0 == state ? _GEN_4495 : 4'h0; // @[DCache.scala 260:17 84:29]
  assign write_buffer_io_enq_bits_size = 3'h0 == state ? _GEN_4494 : 2'h0; // @[DCache.scala 260:17 84:29]
  assign write_buffer_io_deq_ready = write_buffer_axi_busy ? 1'h0 : _GEN_266; // @[DCache.scala 219:31 85:29]
  assign bank_ram_clock = clock;
  assign bank_ram_reset = reset;
  assign bank_ram_io_raddr = bram_use_replace_addr ? bram_replace_addr : _data_raddr_T_2; // @[DCache.scala 104:23]
  assign bank_ram_io_waddr = bram_use_replace_addr ? bram_replace_write_addr : io_cpu_M_mem_va[11:2]; // @[DCache.scala 114:23]
  assign bank_ram_io_wen = |data_wstrb_0; // @[DCache.scala 158:40]
  assign bank_ram_io_wstrb = _data_wstrb_0_T_5 ? io_cpu_M_wmask : bram_replace_wea_0; // @[DCache.scala 180:25]
  assign bank_ram_io_wdata = data_bram_wdata_sel ? io_axi_r_bits_data : io_cpu_M_wdata; // @[DCache.scala 117:32]
  assign tag_ram_clock = clock;
  assign tag_ram_reset = reset;
  assign tag_ram_io_raddr = {{1'd0}, tag_raddr}; // @[DCache.scala 165:22]
  assign tag_ram_io_waddr = {{1'd0}, bram_replace_addr[9:4]}; // @[DCache.scala 170:22]
  assign tag_ram_io_wen = |tag_wstrb_0; // @[DCache.scala 168:38]
  assign tag_ram_io_wstrb = tag_wstrb_0; // @[DCache.scala 169:22]
  assign tag_ram_io_wdata = tag_wdata; // @[DCache.scala 171:22]
  assign bank_ram_1_clock = clock;
  assign bank_ram_1_reset = reset;
  assign bank_ram_1_io_raddr = bram_use_replace_addr ? bram_replace_addr : _data_raddr_T_2; // @[DCache.scala 104:23]
  assign bank_ram_1_io_waddr = bram_use_replace_addr ? bram_replace_write_addr : io_cpu_M_mem_va[11:2]; // @[DCache.scala 114:23]
  assign bank_ram_1_io_wen = |data_wstrb_1; // @[DCache.scala 158:40]
  assign bank_ram_1_io_wstrb = _data_wstrb_1_T_5 ? io_cpu_M_wmask : bram_replace_wea_1; // @[DCache.scala 180:25]
  assign bank_ram_1_io_wdata = data_bram_wdata_sel ? io_axi_r_bits_data : io_cpu_M_wdata; // @[DCache.scala 117:32]
  assign tag_ram_1_clock = clock;
  assign tag_ram_1_reset = reset;
  assign tag_ram_1_io_raddr = {{1'd0}, tag_raddr}; // @[DCache.scala 165:22]
  assign tag_ram_1_io_waddr = {{1'd0}, bram_replace_addr[9:4]}; // @[DCache.scala 170:22]
  assign tag_ram_1_io_wen = |tag_wstrb_1; // @[DCache.scala 168:38]
  assign tag_ram_1_io_wstrb = tag_wstrb_1; // @[DCache.scala 169:22]
  assign tag_ram_1_io_wdata = tag_wdata; // @[DCache.scala 171:22]
  always @(posedge clock) begin
    if (reset) begin // @[DCache.scala 46:20]
      tlb_vpn <= 20'h0; // @[DCache.scala 46:20]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (3'h1 == state) begin // @[DCache.scala 260:17]
        if (io_cpu_tlb_found) begin // @[DCache.scala 343:30]
          tlb_vpn <= _GEN_5158;
        end
      end
    end
    if (reset) begin // @[DCache.scala 46:20]
      tlb_ppn <= 20'h0; // @[DCache.scala 46:20]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (3'h1 == state) begin // @[DCache.scala 260:17]
        if (io_cpu_tlb_found) begin // @[DCache.scala 343:30]
          tlb_ppn <= _GEN_5159;
        end
      end
    end
    if (reset) begin // @[DCache.scala 46:20]
      tlb_uncached <= 1'h0; // @[DCache.scala 46:20]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (3'h1 == state) begin // @[DCache.scala 260:17]
        if (io_cpu_tlb_found) begin // @[DCache.scala 343:30]
          tlb_uncached <= _GEN_5160;
        end
      end
    end
    if (reset) begin // @[DCache.scala 46:20]
      tlb_dirty <= 1'h0; // @[DCache.scala 46:20]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (3'h1 == state) begin // @[DCache.scala 260:17]
        if (io_cpu_tlb_found) begin // @[DCache.scala 343:30]
          tlb_dirty <= _GEN_5161;
        end
      end
    end
    if (reset) begin // @[DCache.scala 46:20]
      tlb_valid <= 1'h0; // @[DCache.scala 46:20]
    end else if (io_cpu_fence_tlb) begin // @[DCache.scala 513:26]
      tlb_valid <= 1'h0; // @[DCache.scala 514:15]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (3'h1 == state) begin // @[DCache.scala 260:17]
        tlb_valid <= _GEN_5169;
      end
    end
    if (reset) begin // @[DCache.scala 65:96]
      state <= 3'h0; // @[DCache.scala 65:96]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (tlb_stall) begin // @[DCache.scala 263:31]
          state <= _GEN_286;
        end else begin
          state <= _GEN_2130;
        end
      end else if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
        state <= _GEN_3963;
      end
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_tlb_found) begin // @[DCache.scala 343:30]
        state <= _GEN_5163;
      end else begin
        state <= 3'h5; // @[DCache.scala 356:25]
      end
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      state <= _GEN_5175;
    end else begin
      state <= _GEN_9406;
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_0_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_0_0 <= _GEN_3970;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_0_0 <= _GEN_9420;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_0_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_0_1 <= _GEN_4098;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_0_1 <= _GEN_9421;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_1_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_1_0 <= _GEN_3971;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_1_0 <= _GEN_9422;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_1_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_1_1 <= _GEN_4099;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_1_1 <= _GEN_9423;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_2_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_2_0 <= _GEN_3972;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_2_0 <= _GEN_9424;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_2_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_2_1 <= _GEN_4100;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_2_1 <= _GEN_9425;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_3_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_3_0 <= _GEN_3973;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_3_0 <= _GEN_9426;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_3_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_3_1 <= _GEN_4101;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_3_1 <= _GEN_9427;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_4_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_4_0 <= _GEN_3974;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_4_0 <= _GEN_9428;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_4_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_4_1 <= _GEN_4102;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_4_1 <= _GEN_9429;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_5_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_5_0 <= _GEN_3975;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_5_0 <= _GEN_9430;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_5_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_5_1 <= _GEN_4103;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_5_1 <= _GEN_9431;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_6_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_6_0 <= _GEN_3976;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_6_0 <= _GEN_9432;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_6_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_6_1 <= _GEN_4104;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_6_1 <= _GEN_9433;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_7_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_7_0 <= _GEN_3977;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_7_0 <= _GEN_9434;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_7_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_7_1 <= _GEN_4105;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_7_1 <= _GEN_9435;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_8_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_8_0 <= _GEN_3978;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_8_0 <= _GEN_9436;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_8_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_8_1 <= _GEN_4106;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_8_1 <= _GEN_9437;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_9_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_9_0 <= _GEN_3979;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_9_0 <= _GEN_9438;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_9_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_9_1 <= _GEN_4107;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_9_1 <= _GEN_9439;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_10_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_10_0 <= _GEN_3980;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_10_0 <= _GEN_9440;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_10_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_10_1 <= _GEN_4108;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_10_1 <= _GEN_9441;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_11_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_11_0 <= _GEN_3981;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_11_0 <= _GEN_9442;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_11_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_11_1 <= _GEN_4109;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_11_1 <= _GEN_9443;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_12_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_12_0 <= _GEN_3982;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_12_0 <= _GEN_9444;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_12_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_12_1 <= _GEN_4110;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_12_1 <= _GEN_9445;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_13_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_13_0 <= _GEN_3983;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_13_0 <= _GEN_9446;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_13_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_13_1 <= _GEN_4111;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_13_1 <= _GEN_9447;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_14_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_14_0 <= _GEN_3984;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_14_0 <= _GEN_9448;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_14_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_14_1 <= _GEN_4112;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_14_1 <= _GEN_9449;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_15_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_15_0 <= _GEN_3985;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_15_0 <= _GEN_9450;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_15_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_15_1 <= _GEN_4113;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_15_1 <= _GEN_9451;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_16_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_16_0 <= _GEN_3986;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_16_0 <= _GEN_9452;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_16_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_16_1 <= _GEN_4114;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_16_1 <= _GEN_9453;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_17_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_17_0 <= _GEN_3987;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_17_0 <= _GEN_9454;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_17_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_17_1 <= _GEN_4115;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_17_1 <= _GEN_9455;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_18_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_18_0 <= _GEN_3988;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_18_0 <= _GEN_9456;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_18_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_18_1 <= _GEN_4116;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_18_1 <= _GEN_9457;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_19_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_19_0 <= _GEN_3989;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_19_0 <= _GEN_9458;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_19_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_19_1 <= _GEN_4117;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_19_1 <= _GEN_9459;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_20_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_20_0 <= _GEN_3990;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_20_0 <= _GEN_9460;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_20_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_20_1 <= _GEN_4118;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_20_1 <= _GEN_9461;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_21_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_21_0 <= _GEN_3991;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_21_0 <= _GEN_9462;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_21_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_21_1 <= _GEN_4119;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_21_1 <= _GEN_9463;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_22_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_22_0 <= _GEN_3992;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_22_0 <= _GEN_9464;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_22_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_22_1 <= _GEN_4120;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_22_1 <= _GEN_9465;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_23_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_23_0 <= _GEN_3993;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_23_0 <= _GEN_9466;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_23_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_23_1 <= _GEN_4121;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_23_1 <= _GEN_9467;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_24_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_24_0 <= _GEN_3994;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_24_0 <= _GEN_9468;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_24_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_24_1 <= _GEN_4122;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_24_1 <= _GEN_9469;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_25_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_25_0 <= _GEN_3995;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_25_0 <= _GEN_9470;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_25_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_25_1 <= _GEN_4123;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_25_1 <= _GEN_9471;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_26_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_26_0 <= _GEN_3996;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_26_0 <= _GEN_9472;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_26_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_26_1 <= _GEN_4124;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_26_1 <= _GEN_9473;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_27_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_27_0 <= _GEN_3997;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_27_0 <= _GEN_9474;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_27_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_27_1 <= _GEN_4125;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_27_1 <= _GEN_9475;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_28_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_28_0 <= _GEN_3998;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_28_0 <= _GEN_9476;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_28_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_28_1 <= _GEN_4126;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_28_1 <= _GEN_9477;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_29_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_29_0 <= _GEN_3999;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_29_0 <= _GEN_9478;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_29_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_29_1 <= _GEN_4127;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_29_1 <= _GEN_9479;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_30_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_30_0 <= _GEN_4000;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_30_0 <= _GEN_9480;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_30_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_30_1 <= _GEN_4128;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_30_1 <= _GEN_9481;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_31_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_31_0 <= _GEN_4001;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_31_0 <= _GEN_9482;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_31_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_31_1 <= _GEN_4129;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_31_1 <= _GEN_9483;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_32_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_32_0 <= _GEN_4002;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_32_0 <= _GEN_9484;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_32_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_32_1 <= _GEN_4130;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_32_1 <= _GEN_9485;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_33_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_33_0 <= _GEN_4003;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_33_0 <= _GEN_9486;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_33_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_33_1 <= _GEN_4131;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_33_1 <= _GEN_9487;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_34_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_34_0 <= _GEN_4004;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_34_0 <= _GEN_9488;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_34_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_34_1 <= _GEN_4132;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_34_1 <= _GEN_9489;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_35_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_35_0 <= _GEN_4005;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_35_0 <= _GEN_9490;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_35_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_35_1 <= _GEN_4133;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_35_1 <= _GEN_9491;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_36_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_36_0 <= _GEN_4006;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_36_0 <= _GEN_9492;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_36_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_36_1 <= _GEN_4134;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_36_1 <= _GEN_9493;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_37_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_37_0 <= _GEN_4007;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_37_0 <= _GEN_9494;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_37_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_37_1 <= _GEN_4135;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_37_1 <= _GEN_9495;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_38_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_38_0 <= _GEN_4008;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_38_0 <= _GEN_9496;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_38_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_38_1 <= _GEN_4136;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_38_1 <= _GEN_9497;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_39_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_39_0 <= _GEN_4009;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_39_0 <= _GEN_9498;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_39_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_39_1 <= _GEN_4137;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_39_1 <= _GEN_9499;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_40_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_40_0 <= _GEN_4010;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_40_0 <= _GEN_9500;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_40_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_40_1 <= _GEN_4138;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_40_1 <= _GEN_9501;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_41_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_41_0 <= _GEN_4011;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_41_0 <= _GEN_9502;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_41_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_41_1 <= _GEN_4139;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_41_1 <= _GEN_9503;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_42_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_42_0 <= _GEN_4012;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_42_0 <= _GEN_9504;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_42_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_42_1 <= _GEN_4140;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_42_1 <= _GEN_9505;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_43_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_43_0 <= _GEN_4013;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_43_0 <= _GEN_9506;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_43_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_43_1 <= _GEN_4141;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_43_1 <= _GEN_9507;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_44_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_44_0 <= _GEN_4014;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_44_0 <= _GEN_9508;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_44_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_44_1 <= _GEN_4142;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_44_1 <= _GEN_9509;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_45_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_45_0 <= _GEN_4015;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_45_0 <= _GEN_9510;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_45_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_45_1 <= _GEN_4143;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_45_1 <= _GEN_9511;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_46_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_46_0 <= _GEN_4016;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_46_0 <= _GEN_9512;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_46_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_46_1 <= _GEN_4144;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_46_1 <= _GEN_9513;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_47_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_47_0 <= _GEN_4017;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_47_0 <= _GEN_9514;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_47_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_47_1 <= _GEN_4145;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_47_1 <= _GEN_9515;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_48_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_48_0 <= _GEN_4018;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_48_0 <= _GEN_9516;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_48_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_48_1 <= _GEN_4146;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_48_1 <= _GEN_9517;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_49_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_49_0 <= _GEN_4019;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_49_0 <= _GEN_9518;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_49_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_49_1 <= _GEN_4147;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_49_1 <= _GEN_9519;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_50_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_50_0 <= _GEN_4020;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_50_0 <= _GEN_9520;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_50_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_50_1 <= _GEN_4148;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_50_1 <= _GEN_9521;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_51_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_51_0 <= _GEN_4021;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_51_0 <= _GEN_9522;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_51_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_51_1 <= _GEN_4149;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_51_1 <= _GEN_9523;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_52_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_52_0 <= _GEN_4022;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_52_0 <= _GEN_9524;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_52_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_52_1 <= _GEN_4150;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_52_1 <= _GEN_9525;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_53_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_53_0 <= _GEN_4023;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_53_0 <= _GEN_9526;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_53_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_53_1 <= _GEN_4151;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_53_1 <= _GEN_9527;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_54_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_54_0 <= _GEN_4024;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_54_0 <= _GEN_9528;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_54_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_54_1 <= _GEN_4152;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_54_1 <= _GEN_9529;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_55_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_55_0 <= _GEN_4025;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_55_0 <= _GEN_9530;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_55_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_55_1 <= _GEN_4153;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_55_1 <= _GEN_9531;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_56_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_56_0 <= _GEN_4026;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_56_0 <= _GEN_9532;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_56_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_56_1 <= _GEN_4154;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_56_1 <= _GEN_9533;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_57_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_57_0 <= _GEN_4027;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_57_0 <= _GEN_9534;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_57_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_57_1 <= _GEN_4155;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_57_1 <= _GEN_9535;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_58_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_58_0 <= _GEN_4028;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_58_0 <= _GEN_9536;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_58_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_58_1 <= _GEN_4156;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_58_1 <= _GEN_9537;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_59_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_59_0 <= _GEN_4029;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_59_0 <= _GEN_9538;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_59_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_59_1 <= _GEN_4157;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_59_1 <= _GEN_9539;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_60_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_60_0 <= _GEN_4030;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_60_0 <= _GEN_9540;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_60_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_60_1 <= _GEN_4158;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_60_1 <= _GEN_9541;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_61_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_61_0 <= _GEN_4031;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_61_0 <= _GEN_9542;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_61_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_61_1 <= _GEN_4159;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_61_1 <= _GEN_9543;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_62_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_62_0 <= _GEN_4032;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_62_0 <= _GEN_9544;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_62_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_62_1 <= _GEN_4160;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_62_1 <= _GEN_9545;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_63_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_63_0 <= _GEN_4033;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_63_0 <= _GEN_9546;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_63_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_63_1 <= _GEN_4161;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_63_1 <= _GEN_9547;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_64_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_64_0 <= _GEN_4034;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_64_0 <= _GEN_9548;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_64_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_64_1 <= _GEN_4162;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_64_1 <= _GEN_9549;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_65_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_65_0 <= _GEN_4035;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_65_0 <= _GEN_9550;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_65_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_65_1 <= _GEN_4163;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_65_1 <= _GEN_9551;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_66_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_66_0 <= _GEN_4036;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_66_0 <= _GEN_9552;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_66_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_66_1 <= _GEN_4164;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_66_1 <= _GEN_9553;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_67_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_67_0 <= _GEN_4037;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_67_0 <= _GEN_9554;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_67_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_67_1 <= _GEN_4165;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_67_1 <= _GEN_9555;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_68_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_68_0 <= _GEN_4038;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_68_0 <= _GEN_9556;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_68_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_68_1 <= _GEN_4166;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_68_1 <= _GEN_9557;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_69_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_69_0 <= _GEN_4039;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_69_0 <= _GEN_9558;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_69_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_69_1 <= _GEN_4167;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_69_1 <= _GEN_9559;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_70_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_70_0 <= _GEN_4040;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_70_0 <= _GEN_9560;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_70_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_70_1 <= _GEN_4168;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_70_1 <= _GEN_9561;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_71_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_71_0 <= _GEN_4041;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_71_0 <= _GEN_9562;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_71_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_71_1 <= _GEN_4169;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_71_1 <= _GEN_9563;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_72_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_72_0 <= _GEN_4042;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_72_0 <= _GEN_9564;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_72_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_72_1 <= _GEN_4170;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_72_1 <= _GEN_9565;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_73_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_73_0 <= _GEN_4043;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_73_0 <= _GEN_9566;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_73_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_73_1 <= _GEN_4171;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_73_1 <= _GEN_9567;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_74_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_74_0 <= _GEN_4044;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_74_0 <= _GEN_9568;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_74_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_74_1 <= _GEN_4172;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_74_1 <= _GEN_9569;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_75_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_75_0 <= _GEN_4045;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_75_0 <= _GEN_9570;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_75_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_75_1 <= _GEN_4173;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_75_1 <= _GEN_9571;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_76_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_76_0 <= _GEN_4046;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_76_0 <= _GEN_9572;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_76_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_76_1 <= _GEN_4174;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_76_1 <= _GEN_9573;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_77_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_77_0 <= _GEN_4047;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_77_0 <= _GEN_9574;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_77_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_77_1 <= _GEN_4175;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_77_1 <= _GEN_9575;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_78_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_78_0 <= _GEN_4048;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_78_0 <= _GEN_9576;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_78_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_78_1 <= _GEN_4176;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_78_1 <= _GEN_9577;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_79_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_79_0 <= _GEN_4049;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_79_0 <= _GEN_9578;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_79_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_79_1 <= _GEN_4177;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_79_1 <= _GEN_9579;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_80_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_80_0 <= _GEN_4050;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_80_0 <= _GEN_9580;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_80_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_80_1 <= _GEN_4178;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_80_1 <= _GEN_9581;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_81_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_81_0 <= _GEN_4051;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_81_0 <= _GEN_9582;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_81_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_81_1 <= _GEN_4179;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_81_1 <= _GEN_9583;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_82_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_82_0 <= _GEN_4052;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_82_0 <= _GEN_9584;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_82_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_82_1 <= _GEN_4180;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_82_1 <= _GEN_9585;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_83_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_83_0 <= _GEN_4053;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_83_0 <= _GEN_9586;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_83_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_83_1 <= _GEN_4181;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_83_1 <= _GEN_9587;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_84_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_84_0 <= _GEN_4054;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_84_0 <= _GEN_9588;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_84_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_84_1 <= _GEN_4182;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_84_1 <= _GEN_9589;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_85_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_85_0 <= _GEN_4055;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_85_0 <= _GEN_9590;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_85_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_85_1 <= _GEN_4183;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_85_1 <= _GEN_9591;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_86_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_86_0 <= _GEN_4056;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_86_0 <= _GEN_9592;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_86_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_86_1 <= _GEN_4184;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_86_1 <= _GEN_9593;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_87_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_87_0 <= _GEN_4057;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_87_0 <= _GEN_9594;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_87_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_87_1 <= _GEN_4185;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_87_1 <= _GEN_9595;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_88_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_88_0 <= _GEN_4058;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_88_0 <= _GEN_9596;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_88_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_88_1 <= _GEN_4186;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_88_1 <= _GEN_9597;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_89_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_89_0 <= _GEN_4059;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_89_0 <= _GEN_9598;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_89_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_89_1 <= _GEN_4187;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_89_1 <= _GEN_9599;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_90_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_90_0 <= _GEN_4060;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_90_0 <= _GEN_9600;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_90_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_90_1 <= _GEN_4188;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_90_1 <= _GEN_9601;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_91_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_91_0 <= _GEN_4061;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_91_0 <= _GEN_9602;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_91_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_91_1 <= _GEN_4189;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_91_1 <= _GEN_9603;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_92_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_92_0 <= _GEN_4062;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_92_0 <= _GEN_9604;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_92_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_92_1 <= _GEN_4190;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_92_1 <= _GEN_9605;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_93_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_93_0 <= _GEN_4063;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_93_0 <= _GEN_9606;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_93_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_93_1 <= _GEN_4191;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_93_1 <= _GEN_9607;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_94_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_94_0 <= _GEN_4064;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_94_0 <= _GEN_9608;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_94_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_94_1 <= _GEN_4192;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_94_1 <= _GEN_9609;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_95_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_95_0 <= _GEN_4065;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_95_0 <= _GEN_9610;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_95_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_95_1 <= _GEN_4193;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_95_1 <= _GEN_9611;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_96_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_96_0 <= _GEN_4066;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_96_0 <= _GEN_9612;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_96_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_96_1 <= _GEN_4194;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_96_1 <= _GEN_9613;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_97_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_97_0 <= _GEN_4067;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_97_0 <= _GEN_9614;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_97_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_97_1 <= _GEN_4195;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_97_1 <= _GEN_9615;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_98_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_98_0 <= _GEN_4068;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_98_0 <= _GEN_9616;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_98_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_98_1 <= _GEN_4196;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_98_1 <= _GEN_9617;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_99_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_99_0 <= _GEN_4069;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_99_0 <= _GEN_9618;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_99_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_99_1 <= _GEN_4197;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_99_1 <= _GEN_9619;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_100_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_100_0 <= _GEN_4070;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_100_0 <= _GEN_9620;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_100_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_100_1 <= _GEN_4198;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_100_1 <= _GEN_9621;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_101_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_101_0 <= _GEN_4071;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_101_0 <= _GEN_9622;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_101_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_101_1 <= _GEN_4199;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_101_1 <= _GEN_9623;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_102_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_102_0 <= _GEN_4072;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_102_0 <= _GEN_9624;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_102_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_102_1 <= _GEN_4200;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_102_1 <= _GEN_9625;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_103_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_103_0 <= _GEN_4073;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_103_0 <= _GEN_9626;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_103_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_103_1 <= _GEN_4201;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_103_1 <= _GEN_9627;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_104_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_104_0 <= _GEN_4074;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_104_0 <= _GEN_9628;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_104_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_104_1 <= _GEN_4202;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_104_1 <= _GEN_9629;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_105_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_105_0 <= _GEN_4075;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_105_0 <= _GEN_9630;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_105_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_105_1 <= _GEN_4203;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_105_1 <= _GEN_9631;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_106_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_106_0 <= _GEN_4076;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_106_0 <= _GEN_9632;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_106_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_106_1 <= _GEN_4204;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_106_1 <= _GEN_9633;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_107_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_107_0 <= _GEN_4077;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_107_0 <= _GEN_9634;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_107_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_107_1 <= _GEN_4205;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_107_1 <= _GEN_9635;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_108_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_108_0 <= _GEN_4078;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_108_0 <= _GEN_9636;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_108_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_108_1 <= _GEN_4206;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_108_1 <= _GEN_9637;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_109_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_109_0 <= _GEN_4079;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_109_0 <= _GEN_9638;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_109_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_109_1 <= _GEN_4207;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_109_1 <= _GEN_9639;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_110_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_110_0 <= _GEN_4080;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_110_0 <= _GEN_9640;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_110_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_110_1 <= _GEN_4208;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_110_1 <= _GEN_9641;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_111_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_111_0 <= _GEN_4081;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_111_0 <= _GEN_9642;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_111_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_111_1 <= _GEN_4209;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_111_1 <= _GEN_9643;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_112_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_112_0 <= _GEN_4082;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_112_0 <= _GEN_9644;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_112_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_112_1 <= _GEN_4210;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_112_1 <= _GEN_9645;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_113_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_113_0 <= _GEN_4083;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_113_0 <= _GEN_9646;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_113_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_113_1 <= _GEN_4211;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_113_1 <= _GEN_9647;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_114_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_114_0 <= _GEN_4084;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_114_0 <= _GEN_9648;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_114_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_114_1 <= _GEN_4212;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_114_1 <= _GEN_9649;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_115_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_115_0 <= _GEN_4085;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_115_0 <= _GEN_9650;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_115_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_115_1 <= _GEN_4213;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_115_1 <= _GEN_9651;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_116_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_116_0 <= _GEN_4086;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_116_0 <= _GEN_9652;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_116_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_116_1 <= _GEN_4214;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_116_1 <= _GEN_9653;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_117_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_117_0 <= _GEN_4087;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_117_0 <= _GEN_9654;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_117_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_117_1 <= _GEN_4215;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_117_1 <= _GEN_9655;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_118_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_118_0 <= _GEN_4088;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_118_0 <= _GEN_9656;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_118_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_118_1 <= _GEN_4216;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_118_1 <= _GEN_9657;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_119_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_119_0 <= _GEN_4089;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_119_0 <= _GEN_9658;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_119_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_119_1 <= _GEN_4217;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_119_1 <= _GEN_9659;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_120_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_120_0 <= _GEN_4090;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_120_0 <= _GEN_9660;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_120_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_120_1 <= _GEN_4218;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_120_1 <= _GEN_9661;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_121_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_121_0 <= _GEN_4091;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_121_0 <= _GEN_9662;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_121_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_121_1 <= _GEN_4219;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_121_1 <= _GEN_9663;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_122_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_122_0 <= _GEN_4092;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_122_0 <= _GEN_9664;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_122_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_122_1 <= _GEN_4220;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_122_1 <= _GEN_9665;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_123_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_123_0 <= _GEN_4093;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_123_0 <= _GEN_9666;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_123_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_123_1 <= _GEN_4221;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_123_1 <= _GEN_9667;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_124_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_124_0 <= _GEN_4094;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_124_0 <= _GEN_9668;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_124_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_124_1 <= _GEN_4222;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_124_1 <= _GEN_9669;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_125_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_125_0 <= _GEN_4095;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_125_0 <= _GEN_9670;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_125_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_125_1 <= _GEN_4223;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_125_1 <= _GEN_9671;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_126_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_126_0 <= _GEN_4096;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_126_0 <= _GEN_9672;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_126_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_126_1 <= _GEN_4224;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_126_1 <= _GEN_9673;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_127_0 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_127_0 <= _GEN_4097;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_127_0 <= _GEN_9674;
      end
    end
    if (reset) begin // @[DCache.scala 68:22]
      valid_127_1 <= 1'h0; // @[DCache.scala 68:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (!(io_cpu_M_mem_en)) begin // @[DCache.scala 262:22]
        if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
          valid_127_1 <= _GEN_4225;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        valid_127_1 <= _GEN_9675;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_0_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_0_0 <= _GEN_2268;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_0_0 <= _GEN_9148;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_0_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_0_1 <= _GEN_2269;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_0_1 <= _GEN_9149;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_1_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_1_0 <= _GEN_2270;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_1_0 <= _GEN_9150;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_1_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_1_1 <= _GEN_2271;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_1_1 <= _GEN_9151;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_2_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_2_0 <= _GEN_2272;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_2_0 <= _GEN_9152;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_2_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_2_1 <= _GEN_2273;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_2_1 <= _GEN_9153;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_3_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_3_0 <= _GEN_2274;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_3_0 <= _GEN_9154;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_3_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_3_1 <= _GEN_2275;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_3_1 <= _GEN_9155;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_4_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_4_0 <= _GEN_2276;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_4_0 <= _GEN_9156;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_4_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_4_1 <= _GEN_2277;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_4_1 <= _GEN_9157;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_5_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_5_0 <= _GEN_2278;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_5_0 <= _GEN_9158;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_5_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_5_1 <= _GEN_2279;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_5_1 <= _GEN_9159;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_6_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_6_0 <= _GEN_2280;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_6_0 <= _GEN_9160;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_6_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_6_1 <= _GEN_2281;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_6_1 <= _GEN_9161;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_7_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_7_0 <= _GEN_2282;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_7_0 <= _GEN_9162;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_7_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_7_1 <= _GEN_2283;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_7_1 <= _GEN_9163;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_8_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_8_0 <= _GEN_2284;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_8_0 <= _GEN_9164;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_8_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_8_1 <= _GEN_2285;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_8_1 <= _GEN_9165;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_9_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_9_0 <= _GEN_2286;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_9_0 <= _GEN_9166;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_9_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_9_1 <= _GEN_2287;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_9_1 <= _GEN_9167;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_10_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_10_0 <= _GEN_2288;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_10_0 <= _GEN_9168;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_10_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_10_1 <= _GEN_2289;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_10_1 <= _GEN_9169;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_11_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_11_0 <= _GEN_2290;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_11_0 <= _GEN_9170;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_11_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_11_1 <= _GEN_2291;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_11_1 <= _GEN_9171;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_12_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_12_0 <= _GEN_2292;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_12_0 <= _GEN_9172;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_12_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_12_1 <= _GEN_2293;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_12_1 <= _GEN_9173;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_13_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_13_0 <= _GEN_2294;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_13_0 <= _GEN_9174;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_13_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_13_1 <= _GEN_2295;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_13_1 <= _GEN_9175;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_14_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_14_0 <= _GEN_2296;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_14_0 <= _GEN_9176;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_14_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_14_1 <= _GEN_2297;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_14_1 <= _GEN_9177;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_15_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_15_0 <= _GEN_2298;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_15_0 <= _GEN_9178;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_15_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_15_1 <= _GEN_2299;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_15_1 <= _GEN_9179;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_16_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_16_0 <= _GEN_2300;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_16_0 <= _GEN_9180;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_16_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_16_1 <= _GEN_2301;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_16_1 <= _GEN_9181;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_17_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_17_0 <= _GEN_2302;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_17_0 <= _GEN_9182;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_17_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_17_1 <= _GEN_2303;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_17_1 <= _GEN_9183;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_18_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_18_0 <= _GEN_2304;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_18_0 <= _GEN_9184;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_18_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_18_1 <= _GEN_2305;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_18_1 <= _GEN_9185;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_19_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_19_0 <= _GEN_2306;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_19_0 <= _GEN_9186;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_19_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_19_1 <= _GEN_2307;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_19_1 <= _GEN_9187;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_20_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_20_0 <= _GEN_2308;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_20_0 <= _GEN_9188;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_20_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_20_1 <= _GEN_2309;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_20_1 <= _GEN_9189;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_21_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_21_0 <= _GEN_2310;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_21_0 <= _GEN_9190;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_21_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_21_1 <= _GEN_2311;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_21_1 <= _GEN_9191;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_22_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_22_0 <= _GEN_2312;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_22_0 <= _GEN_9192;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_22_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_22_1 <= _GEN_2313;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_22_1 <= _GEN_9193;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_23_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_23_0 <= _GEN_2314;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_23_0 <= _GEN_9194;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_23_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_23_1 <= _GEN_2315;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_23_1 <= _GEN_9195;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_24_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_24_0 <= _GEN_2316;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_24_0 <= _GEN_9196;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_24_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_24_1 <= _GEN_2317;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_24_1 <= _GEN_9197;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_25_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_25_0 <= _GEN_2318;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_25_0 <= _GEN_9198;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_25_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_25_1 <= _GEN_2319;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_25_1 <= _GEN_9199;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_26_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_26_0 <= _GEN_2320;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_26_0 <= _GEN_9200;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_26_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_26_1 <= _GEN_2321;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_26_1 <= _GEN_9201;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_27_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_27_0 <= _GEN_2322;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_27_0 <= _GEN_9202;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_27_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_27_1 <= _GEN_2323;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_27_1 <= _GEN_9203;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_28_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_28_0 <= _GEN_2324;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_28_0 <= _GEN_9204;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_28_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_28_1 <= _GEN_2325;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_28_1 <= _GEN_9205;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_29_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_29_0 <= _GEN_2326;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_29_0 <= _GEN_9206;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_29_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_29_1 <= _GEN_2327;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_29_1 <= _GEN_9207;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_30_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_30_0 <= _GEN_2328;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_30_0 <= _GEN_9208;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_30_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_30_1 <= _GEN_2329;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_30_1 <= _GEN_9209;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_31_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_31_0 <= _GEN_2330;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_31_0 <= _GEN_9210;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_31_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_31_1 <= _GEN_2331;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_31_1 <= _GEN_9211;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_32_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_32_0 <= _GEN_2332;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_32_0 <= _GEN_9212;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_32_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_32_1 <= _GEN_2333;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_32_1 <= _GEN_9213;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_33_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_33_0 <= _GEN_2334;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_33_0 <= _GEN_9214;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_33_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_33_1 <= _GEN_2335;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_33_1 <= _GEN_9215;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_34_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_34_0 <= _GEN_2336;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_34_0 <= _GEN_9216;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_34_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_34_1 <= _GEN_2337;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_34_1 <= _GEN_9217;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_35_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_35_0 <= _GEN_2338;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_35_0 <= _GEN_9218;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_35_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_35_1 <= _GEN_2339;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_35_1 <= _GEN_9219;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_36_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_36_0 <= _GEN_2340;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_36_0 <= _GEN_9220;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_36_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_36_1 <= _GEN_2341;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_36_1 <= _GEN_9221;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_37_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_37_0 <= _GEN_2342;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_37_0 <= _GEN_9222;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_37_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_37_1 <= _GEN_2343;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_37_1 <= _GEN_9223;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_38_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_38_0 <= _GEN_2344;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_38_0 <= _GEN_9224;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_38_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_38_1 <= _GEN_2345;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_38_1 <= _GEN_9225;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_39_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_39_0 <= _GEN_2346;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_39_0 <= _GEN_9226;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_39_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_39_1 <= _GEN_2347;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_39_1 <= _GEN_9227;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_40_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_40_0 <= _GEN_2348;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_40_0 <= _GEN_9228;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_40_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_40_1 <= _GEN_2349;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_40_1 <= _GEN_9229;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_41_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_41_0 <= _GEN_2350;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_41_0 <= _GEN_9230;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_41_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_41_1 <= _GEN_2351;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_41_1 <= _GEN_9231;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_42_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_42_0 <= _GEN_2352;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_42_0 <= _GEN_9232;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_42_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_42_1 <= _GEN_2353;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_42_1 <= _GEN_9233;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_43_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_43_0 <= _GEN_2354;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_43_0 <= _GEN_9234;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_43_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_43_1 <= _GEN_2355;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_43_1 <= _GEN_9235;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_44_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_44_0 <= _GEN_2356;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_44_0 <= _GEN_9236;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_44_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_44_1 <= _GEN_2357;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_44_1 <= _GEN_9237;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_45_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_45_0 <= _GEN_2358;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_45_0 <= _GEN_9238;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_45_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_45_1 <= _GEN_2359;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_45_1 <= _GEN_9239;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_46_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_46_0 <= _GEN_2360;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_46_0 <= _GEN_9240;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_46_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_46_1 <= _GEN_2361;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_46_1 <= _GEN_9241;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_47_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_47_0 <= _GEN_2362;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_47_0 <= _GEN_9242;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_47_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_47_1 <= _GEN_2363;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_47_1 <= _GEN_9243;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_48_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_48_0 <= _GEN_2364;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_48_0 <= _GEN_9244;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_48_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_48_1 <= _GEN_2365;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_48_1 <= _GEN_9245;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_49_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_49_0 <= _GEN_2366;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_49_0 <= _GEN_9246;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_49_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_49_1 <= _GEN_2367;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_49_1 <= _GEN_9247;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_50_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_50_0 <= _GEN_2368;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_50_0 <= _GEN_9248;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_50_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_50_1 <= _GEN_2369;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_50_1 <= _GEN_9249;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_51_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_51_0 <= _GEN_2370;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_51_0 <= _GEN_9250;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_51_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_51_1 <= _GEN_2371;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_51_1 <= _GEN_9251;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_52_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_52_0 <= _GEN_2372;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_52_0 <= _GEN_9252;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_52_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_52_1 <= _GEN_2373;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_52_1 <= _GEN_9253;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_53_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_53_0 <= _GEN_2374;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_53_0 <= _GEN_9254;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_53_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_53_1 <= _GEN_2375;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_53_1 <= _GEN_9255;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_54_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_54_0 <= _GEN_2376;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_54_0 <= _GEN_9256;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_54_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_54_1 <= _GEN_2377;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_54_1 <= _GEN_9257;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_55_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_55_0 <= _GEN_2378;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_55_0 <= _GEN_9258;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_55_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_55_1 <= _GEN_2379;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_55_1 <= _GEN_9259;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_56_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_56_0 <= _GEN_2380;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_56_0 <= _GEN_9260;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_56_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_56_1 <= _GEN_2381;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_56_1 <= _GEN_9261;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_57_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_57_0 <= _GEN_2382;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_57_0 <= _GEN_9262;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_57_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_57_1 <= _GEN_2383;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_57_1 <= _GEN_9263;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_58_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_58_0 <= _GEN_2384;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_58_0 <= _GEN_9264;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_58_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_58_1 <= _GEN_2385;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_58_1 <= _GEN_9265;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_59_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_59_0 <= _GEN_2386;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_59_0 <= _GEN_9266;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_59_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_59_1 <= _GEN_2387;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_59_1 <= _GEN_9267;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_60_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_60_0 <= _GEN_2388;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_60_0 <= _GEN_9268;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_60_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_60_1 <= _GEN_2389;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_60_1 <= _GEN_9269;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_61_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_61_0 <= _GEN_2390;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_61_0 <= _GEN_9270;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_61_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_61_1 <= _GEN_2391;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_61_1 <= _GEN_9271;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_62_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_62_0 <= _GEN_2392;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_62_0 <= _GEN_9272;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_62_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_62_1 <= _GEN_2393;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_62_1 <= _GEN_9273;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_63_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_63_0 <= _GEN_2394;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_63_0 <= _GEN_9274;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_63_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_63_1 <= _GEN_2395;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_63_1 <= _GEN_9275;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_64_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_64_0 <= _GEN_2396;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_64_0 <= _GEN_9276;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_64_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_64_1 <= _GEN_2397;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_64_1 <= _GEN_9277;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_65_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_65_0 <= _GEN_2398;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_65_0 <= _GEN_9278;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_65_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_65_1 <= _GEN_2399;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_65_1 <= _GEN_9279;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_66_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_66_0 <= _GEN_2400;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_66_0 <= _GEN_9280;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_66_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_66_1 <= _GEN_2401;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_66_1 <= _GEN_9281;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_67_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_67_0 <= _GEN_2402;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_67_0 <= _GEN_9282;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_67_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_67_1 <= _GEN_2403;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_67_1 <= _GEN_9283;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_68_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_68_0 <= _GEN_2404;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_68_0 <= _GEN_9284;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_68_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_68_1 <= _GEN_2405;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_68_1 <= _GEN_9285;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_69_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_69_0 <= _GEN_2406;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_69_0 <= _GEN_9286;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_69_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_69_1 <= _GEN_2407;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_69_1 <= _GEN_9287;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_70_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_70_0 <= _GEN_2408;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_70_0 <= _GEN_9288;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_70_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_70_1 <= _GEN_2409;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_70_1 <= _GEN_9289;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_71_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_71_0 <= _GEN_2410;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_71_0 <= _GEN_9290;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_71_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_71_1 <= _GEN_2411;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_71_1 <= _GEN_9291;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_72_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_72_0 <= _GEN_2412;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_72_0 <= _GEN_9292;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_72_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_72_1 <= _GEN_2413;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_72_1 <= _GEN_9293;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_73_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_73_0 <= _GEN_2414;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_73_0 <= _GEN_9294;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_73_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_73_1 <= _GEN_2415;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_73_1 <= _GEN_9295;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_74_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_74_0 <= _GEN_2416;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_74_0 <= _GEN_9296;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_74_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_74_1 <= _GEN_2417;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_74_1 <= _GEN_9297;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_75_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_75_0 <= _GEN_2418;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_75_0 <= _GEN_9298;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_75_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_75_1 <= _GEN_2419;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_75_1 <= _GEN_9299;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_76_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_76_0 <= _GEN_2420;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_76_0 <= _GEN_9300;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_76_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_76_1 <= _GEN_2421;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_76_1 <= _GEN_9301;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_77_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_77_0 <= _GEN_2422;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_77_0 <= _GEN_9302;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_77_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_77_1 <= _GEN_2423;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_77_1 <= _GEN_9303;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_78_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_78_0 <= _GEN_2424;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_78_0 <= _GEN_9304;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_78_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_78_1 <= _GEN_2425;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_78_1 <= _GEN_9305;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_79_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_79_0 <= _GEN_2426;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_79_0 <= _GEN_9306;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_79_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_79_1 <= _GEN_2427;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_79_1 <= _GEN_9307;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_80_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_80_0 <= _GEN_2428;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_80_0 <= _GEN_9308;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_80_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_80_1 <= _GEN_2429;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_80_1 <= _GEN_9309;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_81_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_81_0 <= _GEN_2430;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_81_0 <= _GEN_9310;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_81_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_81_1 <= _GEN_2431;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_81_1 <= _GEN_9311;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_82_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_82_0 <= _GEN_2432;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_82_0 <= _GEN_9312;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_82_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_82_1 <= _GEN_2433;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_82_1 <= _GEN_9313;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_83_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_83_0 <= _GEN_2434;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_83_0 <= _GEN_9314;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_83_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_83_1 <= _GEN_2435;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_83_1 <= _GEN_9315;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_84_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_84_0 <= _GEN_2436;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_84_0 <= _GEN_9316;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_84_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_84_1 <= _GEN_2437;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_84_1 <= _GEN_9317;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_85_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_85_0 <= _GEN_2438;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_85_0 <= _GEN_9318;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_85_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_85_1 <= _GEN_2439;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_85_1 <= _GEN_9319;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_86_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_86_0 <= _GEN_2440;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_86_0 <= _GEN_9320;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_86_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_86_1 <= _GEN_2441;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_86_1 <= _GEN_9321;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_87_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_87_0 <= _GEN_2442;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_87_0 <= _GEN_9322;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_87_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_87_1 <= _GEN_2443;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_87_1 <= _GEN_9323;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_88_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_88_0 <= _GEN_2444;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_88_0 <= _GEN_9324;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_88_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_88_1 <= _GEN_2445;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_88_1 <= _GEN_9325;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_89_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_89_0 <= _GEN_2446;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_89_0 <= _GEN_9326;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_89_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_89_1 <= _GEN_2447;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_89_1 <= _GEN_9327;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_90_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_90_0 <= _GEN_2448;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_90_0 <= _GEN_9328;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_90_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_90_1 <= _GEN_2449;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_90_1 <= _GEN_9329;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_91_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_91_0 <= _GEN_2450;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_91_0 <= _GEN_9330;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_91_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_91_1 <= _GEN_2451;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_91_1 <= _GEN_9331;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_92_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_92_0 <= _GEN_2452;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_92_0 <= _GEN_9332;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_92_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_92_1 <= _GEN_2453;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_92_1 <= _GEN_9333;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_93_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_93_0 <= _GEN_2454;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_93_0 <= _GEN_9334;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_93_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_93_1 <= _GEN_2455;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_93_1 <= _GEN_9335;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_94_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_94_0 <= _GEN_2456;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_94_0 <= _GEN_9336;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_94_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_94_1 <= _GEN_2457;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_94_1 <= _GEN_9337;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_95_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_95_0 <= _GEN_2458;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_95_0 <= _GEN_9338;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_95_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_95_1 <= _GEN_2459;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_95_1 <= _GEN_9339;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_96_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_96_0 <= _GEN_2460;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_96_0 <= _GEN_9340;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_96_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_96_1 <= _GEN_2461;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_96_1 <= _GEN_9341;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_97_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_97_0 <= _GEN_2462;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_97_0 <= _GEN_9342;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_97_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_97_1 <= _GEN_2463;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_97_1 <= _GEN_9343;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_98_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_98_0 <= _GEN_2464;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_98_0 <= _GEN_9344;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_98_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_98_1 <= _GEN_2465;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_98_1 <= _GEN_9345;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_99_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_99_0 <= _GEN_2466;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_99_0 <= _GEN_9346;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_99_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_99_1 <= _GEN_2467;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_99_1 <= _GEN_9347;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_100_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_100_0 <= _GEN_2468;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_100_0 <= _GEN_9348;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_100_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_100_1 <= _GEN_2469;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_100_1 <= _GEN_9349;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_101_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_101_0 <= _GEN_2470;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_101_0 <= _GEN_9350;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_101_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_101_1 <= _GEN_2471;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_101_1 <= _GEN_9351;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_102_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_102_0 <= _GEN_2472;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_102_0 <= _GEN_9352;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_102_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_102_1 <= _GEN_2473;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_102_1 <= _GEN_9353;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_103_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_103_0 <= _GEN_2474;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_103_0 <= _GEN_9354;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_103_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_103_1 <= _GEN_2475;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_103_1 <= _GEN_9355;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_104_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_104_0 <= _GEN_2476;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_104_0 <= _GEN_9356;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_104_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_104_1 <= _GEN_2477;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_104_1 <= _GEN_9357;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_105_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_105_0 <= _GEN_2478;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_105_0 <= _GEN_9358;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_105_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_105_1 <= _GEN_2479;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_105_1 <= _GEN_9359;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_106_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_106_0 <= _GEN_2480;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_106_0 <= _GEN_9360;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_106_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_106_1 <= _GEN_2481;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_106_1 <= _GEN_9361;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_107_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_107_0 <= _GEN_2482;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_107_0 <= _GEN_9362;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_107_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_107_1 <= _GEN_2483;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_107_1 <= _GEN_9363;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_108_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_108_0 <= _GEN_2484;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_108_0 <= _GEN_9364;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_108_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_108_1 <= _GEN_2485;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_108_1 <= _GEN_9365;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_109_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_109_0 <= _GEN_2486;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_109_0 <= _GEN_9366;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_109_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_109_1 <= _GEN_2487;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_109_1 <= _GEN_9367;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_110_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_110_0 <= _GEN_2488;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_110_0 <= _GEN_9368;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_110_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_110_1 <= _GEN_2489;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_110_1 <= _GEN_9369;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_111_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_111_0 <= _GEN_2490;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_111_0 <= _GEN_9370;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_111_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_111_1 <= _GEN_2491;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_111_1 <= _GEN_9371;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_112_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_112_0 <= _GEN_2492;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_112_0 <= _GEN_9372;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_112_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_112_1 <= _GEN_2493;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_112_1 <= _GEN_9373;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_113_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_113_0 <= _GEN_2494;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_113_0 <= _GEN_9374;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_113_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_113_1 <= _GEN_2495;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_113_1 <= _GEN_9375;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_114_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_114_0 <= _GEN_2496;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_114_0 <= _GEN_9376;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_114_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_114_1 <= _GEN_2497;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_114_1 <= _GEN_9377;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_115_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_115_0 <= _GEN_2498;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_115_0 <= _GEN_9378;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_115_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_115_1 <= _GEN_2499;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_115_1 <= _GEN_9379;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_116_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_116_0 <= _GEN_2500;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_116_0 <= _GEN_9380;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_116_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_116_1 <= _GEN_2501;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_116_1 <= _GEN_9381;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_117_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_117_0 <= _GEN_2502;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_117_0 <= _GEN_9382;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_117_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_117_1 <= _GEN_2503;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_117_1 <= _GEN_9383;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_118_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_118_0 <= _GEN_2504;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_118_0 <= _GEN_9384;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_118_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_118_1 <= _GEN_2505;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_118_1 <= _GEN_9385;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_119_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_119_0 <= _GEN_2506;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_119_0 <= _GEN_9386;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_119_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_119_1 <= _GEN_2507;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_119_1 <= _GEN_9387;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_120_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_120_0 <= _GEN_2508;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_120_0 <= _GEN_9388;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_120_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_120_1 <= _GEN_2509;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_120_1 <= _GEN_9389;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_121_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_121_0 <= _GEN_2510;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_121_0 <= _GEN_9390;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_121_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_121_1 <= _GEN_2511;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_121_1 <= _GEN_9391;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_122_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_122_0 <= _GEN_2512;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_122_0 <= _GEN_9392;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_122_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_122_1 <= _GEN_2513;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_122_1 <= _GEN_9393;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_123_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_123_0 <= _GEN_2514;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_123_0 <= _GEN_9394;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_123_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_123_1 <= _GEN_2515;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_123_1 <= _GEN_9395;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_124_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_124_0 <= _GEN_2516;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_124_0 <= _GEN_9396;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_124_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_124_1 <= _GEN_2517;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_124_1 <= _GEN_9397;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_125_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_125_0 <= _GEN_2518;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_125_0 <= _GEN_9398;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_125_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_125_1 <= _GEN_2519;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_125_1 <= _GEN_9399;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_126_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_126_0 <= _GEN_2520;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_126_0 <= _GEN_9400;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_126_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_126_1 <= _GEN_2521;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_126_1 <= _GEN_9401;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_127_0 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_127_0 <= _GEN_2522;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_127_0 <= _GEN_9402;
      end
    end
    if (reset) begin // @[DCache.scala 69:22]
      dirty_127_1 <= 1'h0; // @[DCache.scala 69:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          dirty_127_1 <= _GEN_2523;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        dirty_127_1 <= _GEN_9403;
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_0 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_0 <= _GEN_2140;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_1 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_1 <= _GEN_2141;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_2 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_2 <= _GEN_2142;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_3 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_3 <= _GEN_2143;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_4 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_4 <= _GEN_2144;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_5 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_5 <= _GEN_2145;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_6 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_6 <= _GEN_2146;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_7 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_7 <= _GEN_2147;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_8 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_8 <= _GEN_2148;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_9 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_9 <= _GEN_2149;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_10 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_10 <= _GEN_2150;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_11 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_11 <= _GEN_2151;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_12 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_12 <= _GEN_2152;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_13 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_13 <= _GEN_2153;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_14 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_14 <= _GEN_2154;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_15 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_15 <= _GEN_2155;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_16 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_16 <= _GEN_2156;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_17 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_17 <= _GEN_2157;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_18 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_18 <= _GEN_2158;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_19 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_19 <= _GEN_2159;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_20 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_20 <= _GEN_2160;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_21 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_21 <= _GEN_2161;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_22 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_22 <= _GEN_2162;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_23 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_23 <= _GEN_2163;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_24 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_24 <= _GEN_2164;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_25 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_25 <= _GEN_2165;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_26 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_26 <= _GEN_2166;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_27 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_27 <= _GEN_2167;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_28 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_28 <= _GEN_2168;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_29 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_29 <= _GEN_2169;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_30 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_30 <= _GEN_2170;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_31 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_31 <= _GEN_2171;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_32 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_32 <= _GEN_2172;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_33 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_33 <= _GEN_2173;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_34 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_34 <= _GEN_2174;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_35 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_35 <= _GEN_2175;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_36 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_36 <= _GEN_2176;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_37 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_37 <= _GEN_2177;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_38 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_38 <= _GEN_2178;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_39 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_39 <= _GEN_2179;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_40 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_40 <= _GEN_2180;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_41 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_41 <= _GEN_2181;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_42 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_42 <= _GEN_2182;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_43 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_43 <= _GEN_2183;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_44 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_44 <= _GEN_2184;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_45 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_45 <= _GEN_2185;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_46 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_46 <= _GEN_2186;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_47 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_47 <= _GEN_2187;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_48 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_48 <= _GEN_2188;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_49 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_49 <= _GEN_2189;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_50 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_50 <= _GEN_2190;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_51 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_51 <= _GEN_2191;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_52 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_52 <= _GEN_2192;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_53 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_53 <= _GEN_2193;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_54 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_54 <= _GEN_2194;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_55 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_55 <= _GEN_2195;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_56 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_56 <= _GEN_2196;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_57 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_57 <= _GEN_2197;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_58 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_58 <= _GEN_2198;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_59 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_59 <= _GEN_2199;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_60 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_60 <= _GEN_2200;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_61 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_61 <= _GEN_2201;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_62 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_62 <= _GEN_2202;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_63 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_63 <= _GEN_2203;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_64 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_64 <= _GEN_2204;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_65 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_65 <= _GEN_2205;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_66 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_66 <= _GEN_2206;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_67 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_67 <= _GEN_2207;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_68 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_68 <= _GEN_2208;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_69 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_69 <= _GEN_2209;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_70 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_70 <= _GEN_2210;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_71 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_71 <= _GEN_2211;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_72 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_72 <= _GEN_2212;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_73 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_73 <= _GEN_2213;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_74 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_74 <= _GEN_2214;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_75 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_75 <= _GEN_2215;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_76 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_76 <= _GEN_2216;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_77 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_77 <= _GEN_2217;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_78 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_78 <= _GEN_2218;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_79 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_79 <= _GEN_2219;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_80 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_80 <= _GEN_2220;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_81 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_81 <= _GEN_2221;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_82 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_82 <= _GEN_2222;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_83 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_83 <= _GEN_2223;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_84 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_84 <= _GEN_2224;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_85 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_85 <= _GEN_2225;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_86 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_86 <= _GEN_2226;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_87 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_87 <= _GEN_2227;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_88 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_88 <= _GEN_2228;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_89 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_89 <= _GEN_2229;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_90 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_90 <= _GEN_2230;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_91 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_91 <= _GEN_2231;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_92 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_92 <= _GEN_2232;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_93 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_93 <= _GEN_2233;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_94 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_94 <= _GEN_2234;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_95 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_95 <= _GEN_2235;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_96 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_96 <= _GEN_2236;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_97 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_97 <= _GEN_2237;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_98 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_98 <= _GEN_2238;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_99 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_99 <= _GEN_2239;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_100 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_100 <= _GEN_2240;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_101 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_101 <= _GEN_2241;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_102 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_102 <= _GEN_2242;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_103 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_103 <= _GEN_2243;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_104 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_104 <= _GEN_2244;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_105 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_105 <= _GEN_2245;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_106 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_106 <= _GEN_2246;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_107 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_107 <= _GEN_2247;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_108 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_108 <= _GEN_2248;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_109 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_109 <= _GEN_2249;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_110 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_110 <= _GEN_2250;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_111 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_111 <= _GEN_2251;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_112 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_112 <= _GEN_2252;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_113 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_113 <= _GEN_2253;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_114 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_114 <= _GEN_2254;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_115 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_115 <= _GEN_2255;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_116 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_116 <= _GEN_2256;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_117 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_117 <= _GEN_2257;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_118 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_118 <= _GEN_2258;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_119 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_119 <= _GEN_2259;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_120 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_120 <= _GEN_2260;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_121 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_121 <= _GEN_2261;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_122 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_122 <= _GEN_2262;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_123 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_123 <= _GEN_2263;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_124 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_124 <= _GEN_2264;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_125 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_125 <= _GEN_2265;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_126 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_126 <= _GEN_2266;
        end
      end
    end
    if (reset) begin // @[DCache.scala 70:22]
      lru_127 <= 1'h0; // @[DCache.scala 70:22]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          lru_127 <= _GEN_2267;
        end
      end
    end
    if (reset) begin // @[DCache.scala 72:33]
      tag_wstrb_0 <= 1'h0; // @[DCache.scala 72:33]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          tag_wstrb_0 <= _GEN_9416;
        end
      end
    end
    if (reset) begin // @[DCache.scala 72:33]
      tag_wstrb_1 <= 1'h0; // @[DCache.scala 72:33]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          tag_wstrb_1 <= _GEN_9417;
        end
      end
    end
    if (reset) begin // @[DCache.scala 73:33]
      bram_replace_wea_0 <= 4'h0; // @[DCache.scala 73:33]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_replace_wea_0 <= _GEN_9414;
        end
      end
    end
    if (reset) begin // @[DCache.scala 73:33]
      bram_replace_wea_1 <= 4'h0; // @[DCache.scala 73:33]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_replace_wea_1 <= _GEN_9415;
        end
      end
    end
    if (reset) begin // @[DCache.scala 77:26]
      tag_wdata <= 20'h0; // @[DCache.scala 77:26]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          tag_wdata <= _GEN_9418;
        end
      end
    end
    if (reset) begin // @[DCache.scala 89:40]
      axi_wcnt <= 4'h0; // @[DCache.scala 89:40]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          axi_wcnt <= _GEN_2132;
        end
      end else if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
        axi_wcnt <= _GEN_3964;
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        axi_wcnt <= _GEN_9147;
      end
    end
    if (reset) begin // @[DCache.scala 90:40]
      bram_replace_addr <= 10'h0; // @[DCache.scala 90:40]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          bram_replace_addr <= _GEN_2133;
        end
      end else if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
        bram_replace_addr <= _GEN_3965;
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        bram_replace_addr <= _GEN_9120;
      end
    end
    if (reset) begin // @[DCache.scala 91:40]
      bram_read_ready_addr <= 10'h0; // @[DCache.scala 91:40]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          bram_read_ready_addr <= _GEN_2134;
        end
      end else if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
        bram_read_ready_addr <= _GEN_3966;
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        bram_read_ready_addr <= _GEN_9121;
      end
    end
    if (reset) begin // @[DCache.scala 92:40]
      bram_replace_write_addr <= 10'h0; // @[DCache.scala 92:40]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          bram_replace_write_addr <= _GEN_2135;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        bram_replace_write_addr <= _GEN_9419;
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_0 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_0 <= _GEN_9122;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_1 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_1 <= _GEN_9123;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_2 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_2 <= _GEN_9124;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_3 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_3 <= _GEN_9125;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_4 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_4 <= _GEN_9126;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_5 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_5 <= _GEN_9127;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_6 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_6 <= _GEN_9128;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_7 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_7 <= _GEN_9129;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_8 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_8 <= _GEN_9130;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_9 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_9 <= _GEN_9131;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_10 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_10 <= _GEN_9132;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_11 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_11 <= _GEN_9133;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_12 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_12 <= _GEN_9134;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_13 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_13 <= _GEN_9135;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_14 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_14 <= _GEN_9136;
        end
      end
    end
    if (reset) begin // @[DCache.scala 94:40]
      bram_r_buffer_15 <= 32'h0; // @[DCache.scala 94:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          bram_r_buffer_15 <= _GEN_9137;
        end
      end
    end
    if (reset) begin // @[DCache.scala 95:40]
      bram_use_replace_addr <= 1'h0; // @[DCache.scala 95:40]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          bram_use_replace_addr <= _GEN_2137;
        end
      end else if (io_cpu_M_fence_d) begin // @[DCache.scala 322:29]
        bram_use_replace_addr <= _GEN_3968;
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        bram_use_replace_addr <= _GEN_9405;
      end
    end
    if (reset) begin // @[DCache.scala 97:40]
      fence_working <= 1'h0; // @[DCache.scala 97:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          fence_working <= _GEN_9404;
        end
      end
    end
    if (reset) begin // @[DCache.scala 98:40]
      replace_working <= 1'h0; // @[DCache.scala 98:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          replace_working <= _GEN_9676;
        end
      end
    end
    if (reset) begin // @[DCache.scala 99:40]
      ar_handshake <= 1'h0; // @[DCache.scala 99:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          ar_handshake <= _GEN_9413;
        end
      end
    end
    if (reset) begin // @[DCache.scala 100:40]
      aw_handshake <= 1'h0; // @[DCache.scala 100:40]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
        if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
          aw_handshake <= _GEN_9146;
        end
      end
    end
    if (reset) begin // @[DCache.scala 101:40]
      replace_writeback <= 1'h0; // @[DCache.scala 101:40]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          replace_writeback <= _GEN_2139;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        replace_writeback <= _GEN_9407;
      end
    end
    if (reset) begin // @[DCache.scala 141:28]
      saved_rdata <= 32'h0; // @[DCache.scala 141:28]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          saved_rdata <= _GEN_2524;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (3'h2 == state) begin // @[DCache.scala 260:17]
        saved_rdata <= _GEN_5174;
      end
    end
    if (reset) begin // @[DCache.scala 144:35]
      last_line_addr <= 10'h0; // @[DCache.scala 144:35]
    end else if (bram_use_replace_addr) begin // @[DCache.scala 114:23]
      last_line_addr <= bram_replace_write_addr;
    end else begin
      last_line_addr <= io_cpu_M_mem_va[11:2];
    end
    if (reset) begin // @[DCache.scala 145:35]
      last_wea_0 <= 32'h0; // @[DCache.scala 145:35]
    end else begin
      last_wea_0 <= _last_wea_0_T_12; // @[DCache.scala 186:17]
    end
    if (reset) begin // @[DCache.scala 145:35]
      last_wea_1 <= 32'h0; // @[DCache.scala 145:35]
    end else begin
      last_wea_1 <= _last_wea_1_T_12; // @[DCache.scala 186:17]
    end
    if (reset) begin // @[DCache.scala 146:35]
      last_wdata <= 32'h0; // @[DCache.scala 146:35]
    end else if (data_bram_wdata_sel) begin // @[DCache.scala 117:32]
      last_wdata <= io_axi_r_bits_data;
    end else begin
      last_wdata <= io_cpu_M_wdata;
    end
    if (reset) begin // @[DCache.scala 197:38]
      write_buffer_axi_busy <= 1'h0; // @[DCache.scala 197:38]
    end else if (write_buffer_axi_busy) begin // @[DCache.scala 219:31]
      if (_T_2) begin // @[DCache.scala 227:25]
        write_buffer_axi_busy <= 1'h0; // @[DCache.scala 228:29]
      end
    end else begin
      write_buffer_axi_busy <= _GEN_275;
    end
    if (reset) begin // @[DCache.scala 199:24]
      ar_addr <= 32'h0; // @[DCache.scala 199:24]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          ar_addr <= _GEN_2126;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        ar_addr <= _GEN_9408;
      end
    end
    if (reset) begin // @[DCache.scala 199:24]
      ar_len <= 8'h0; // @[DCache.scala 199:24]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          ar_len <= _GEN_2127;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        ar_len <= _GEN_9409;
      end
    end
    if (reset) begin // @[DCache.scala 199:24]
      ar_size <= 3'h0; // @[DCache.scala 199:24]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          ar_size <= _GEN_2128;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        ar_size <= _GEN_9410;
      end
    end
    if (reset) begin // @[DCache.scala 200:24]
      arvalid <= 1'h0; // @[DCache.scala 200:24]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          arvalid <= _GEN_2129;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (3'h2 == state) begin // @[DCache.scala 260:17]
        arvalid <= _GEN_5173;
      end else begin
        arvalid <= _GEN_9411;
      end
    end
    if (reset) begin // @[DCache.scala 203:23]
      rready <= 1'h0; // @[DCache.scala 203:23]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          rready <= _GEN_2131;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        rready <= _GEN_9412;
      end
    end
    if (reset) begin // @[DCache.scala 205:24]
      aw_addr <= 32'h0; // @[DCache.scala 205:24]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      aw_addr <= _GEN_281;
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      aw_addr <= _GEN_281;
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      aw_addr <= _GEN_281;
    end else begin
      aw_addr <= _GEN_9138;
    end
    if (reset) begin // @[DCache.scala 205:24]
      aw_len <= 8'h0; // @[DCache.scala 205:24]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      aw_len <= _GEN_285;
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      aw_len <= _GEN_285;
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      aw_len <= _GEN_285;
    end else begin
      aw_len <= _GEN_9139;
    end
    if (reset) begin // @[DCache.scala 205:24]
      aw_size <= 3'h0; // @[DCache.scala 205:24]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      aw_size <= _GEN_282;
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      aw_size <= _GEN_282;
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      aw_size <= _GEN_282;
    end else begin
      aw_size <= _GEN_9140;
    end
    if (reset) begin // @[DCache.scala 206:24]
      awvalid <= 1'h0; // @[DCache.scala 206:24]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      awvalid <= _GEN_276;
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      awvalid <= _GEN_276;
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      awvalid <= _GEN_276;
    end else begin
      awvalid <= _GEN_9141;
    end
    if (reset) begin // @[DCache.scala 209:23]
      w_data <= 32'h0; // @[DCache.scala 209:23]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      w_data <= _GEN_283;
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      w_data <= _GEN_283;
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      w_data <= _GEN_283;
    end else begin
      w_data <= _GEN_9142;
    end
    if (reset) begin // @[DCache.scala 209:23]
      w_strb <= 4'h0; // @[DCache.scala 209:23]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      w_strb <= _GEN_284;
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      w_strb <= _GEN_284;
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      w_strb <= _GEN_284;
    end else begin
      w_strb <= _GEN_9143;
    end
    if (reset) begin // @[DCache.scala 209:23]
      w_last <= 1'h0; // @[DCache.scala 209:23]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      w_last <= _GEN_278;
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      w_last <= _GEN_278;
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      w_last <= _GEN_278;
    end else begin
      w_last <= _GEN_9144;
    end
    if (reset) begin // @[DCache.scala 210:23]
      wvalid <= 1'h0; // @[DCache.scala 210:23]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      wvalid <= _GEN_277;
    end else if (3'h1 == state) begin // @[DCache.scala 260:17]
      wvalid <= _GEN_277;
    end else if (3'h2 == state) begin // @[DCache.scala 260:17]
      wvalid <= _GEN_277;
    end else begin
      wvalid <= _GEN_9145;
    end
    if (reset) begin // @[DCache.scala 216:41]
      current_mmio_write_saved <= 1'h0; // @[DCache.scala 216:41]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (!(tlb_stall)) begin // @[DCache.scala 263:31]
          current_mmio_write_saved <= _GEN_2125;
        end
      end
    end
    tlb2_vpn <= _GEN_15206[18:0]; // @[DCache.scala 245:{21,21}]
    if (reset) begin // @[DCache.scala 250:25]
      data_tlb_refill <= 1'h0; // @[DCache.scala 250:25]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (3'h1 == state) begin // @[DCache.scala 260:17]
        if (!(io_cpu_tlb_found)) begin // @[DCache.scala 343:30]
          data_tlb_refill <= 1'h1; // @[DCache.scala 357:25]
        end
      end else if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        data_tlb_refill <= _GEN_9678;
      end
    end
    if (reset) begin // @[DCache.scala 250:25]
      data_tlb_invalid <= 1'h0; // @[DCache.scala 250:25]
    end else if (!(3'h0 == state)) begin // @[DCache.scala 260:17]
      if (3'h1 == state) begin // @[DCache.scala 260:17]
        if (io_cpu_tlb_found) begin // @[DCache.scala 343:30]
          data_tlb_invalid <= _GEN_5164;
        end
      end else if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        data_tlb_invalid <= _GEN_9677;
      end
    end
    if (reset) begin // @[DCache.scala 250:25]
      data_tlb_mod <= 1'h0; // @[DCache.scala 250:25]
    end else if (3'h0 == state) begin // @[DCache.scala 260:17]
      if (io_cpu_M_mem_en) begin // @[DCache.scala 262:22]
        if (tlb_stall) begin // @[DCache.scala 263:31]
          data_tlb_mod <= _GEN_287;
        end
      end
    end else if (!(3'h1 == state)) begin // @[DCache.scala 260:17]
      if (!(3'h2 == state)) begin // @[DCache.scala 260:17]
        data_tlb_mod <= _GEN_9679;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlb_vpn = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  tlb_ppn = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  tlb_uncached = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  tlb_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  tlb_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  valid_0_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_0_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_1_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_2_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_2_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_3_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_3_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_4_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_4_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_5_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_5_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_6_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_6_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_7_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_7_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_8_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_8_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_9_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_9_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_10_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_10_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_11_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_11_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_12_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_12_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_13_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_13_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_14_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_14_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_15_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_15_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_16_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_16_1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_17_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_17_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_18_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_18_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_19_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_19_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_20_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_20_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_21_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_21_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_22_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_22_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_23_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_23_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_24_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_24_1 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_25_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_25_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_26_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_26_1 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_27_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_27_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_28_0 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_28_1 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_29_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_29_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_30_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_30_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_31_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_31_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_32_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_32_1 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_33_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_33_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_34_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_34_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_35_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_35_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_36_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_36_1 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_37_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_37_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_38_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_38_1 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_39_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_39_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_40_0 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_40_1 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_41_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_41_1 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_42_0 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_42_1 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_43_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_43_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_44_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_44_1 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_45_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_45_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_46_0 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_46_1 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_47_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_47_1 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_48_0 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_48_1 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_49_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_49_1 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_50_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_50_1 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_51_0 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_51_1 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_52_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_52_1 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_53_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_53_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_54_0 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_54_1 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_55_0 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_55_1 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_56_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_56_1 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_57_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_57_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_58_0 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_58_1 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_59_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_59_1 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_60_0 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_60_1 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_61_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_61_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_62_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_62_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_63_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_63_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_64_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_64_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_65_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_65_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_66_0 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_66_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_67_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_67_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_68_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_68_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_69_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_69_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_70_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_70_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_71_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_71_1 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_72_0 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_72_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_73_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_73_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_74_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_74_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_75_0 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_75_1 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_76_0 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_76_1 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_77_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_77_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_78_0 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_78_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_79_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_79_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_80_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_80_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_81_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_81_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_82_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_82_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_83_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_83_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_84_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_84_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_85_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_85_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_86_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_86_1 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_87_0 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_87_1 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_88_0 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_88_1 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_89_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_89_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_90_0 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_90_1 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_91_0 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_91_1 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_92_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_92_1 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_93_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_93_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_94_0 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_94_1 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_95_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_95_1 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_96_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_96_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_97_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_97_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_98_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_98_1 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_99_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_99_1 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_100_0 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_100_1 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_101_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_101_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_102_0 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_102_1 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_103_0 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_103_1 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_104_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_104_1 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_105_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_105_1 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_106_0 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_106_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_107_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_107_1 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_108_0 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_108_1 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_109_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_109_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_110_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_110_1 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_111_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_111_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_112_0 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_112_1 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_113_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_113_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_114_0 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_114_1 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_115_0 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_115_1 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_116_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_116_1 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_117_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_117_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_118_0 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_118_1 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_119_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_119_1 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_120_0 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_120_1 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_121_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_121_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_122_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_122_1 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_123_0 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_123_1 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_124_0 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_124_1 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_125_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_125_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_126_0 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_126_1 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_127_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_127_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  dirty_0_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  dirty_0_1 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  dirty_1_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  dirty_1_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  dirty_2_0 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  dirty_2_1 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  dirty_3_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  dirty_3_1 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  dirty_4_0 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  dirty_4_1 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  dirty_5_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  dirty_5_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  dirty_6_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  dirty_6_1 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  dirty_7_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  dirty_7_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  dirty_8_0 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  dirty_8_1 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  dirty_9_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  dirty_9_1 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  dirty_10_0 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  dirty_10_1 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  dirty_11_0 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  dirty_11_1 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  dirty_12_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  dirty_12_1 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  dirty_13_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  dirty_13_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  dirty_14_0 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  dirty_14_1 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  dirty_15_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  dirty_15_1 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  dirty_16_0 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  dirty_16_1 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  dirty_17_0 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  dirty_17_1 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  dirty_18_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  dirty_18_1 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  dirty_19_0 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  dirty_19_1 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  dirty_20_0 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  dirty_20_1 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  dirty_21_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  dirty_21_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  dirty_22_0 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  dirty_22_1 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  dirty_23_0 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  dirty_23_1 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  dirty_24_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  dirty_24_1 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  dirty_25_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  dirty_25_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  dirty_26_0 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  dirty_26_1 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  dirty_27_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  dirty_27_1 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  dirty_28_0 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  dirty_28_1 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  dirty_29_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  dirty_29_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  dirty_30_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  dirty_30_1 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  dirty_31_0 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  dirty_31_1 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  dirty_32_0 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  dirty_32_1 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  dirty_33_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  dirty_33_1 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  dirty_34_0 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  dirty_34_1 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  dirty_35_0 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  dirty_35_1 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  dirty_36_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  dirty_36_1 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  dirty_37_0 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  dirty_37_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  dirty_38_0 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  dirty_38_1 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  dirty_39_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  dirty_39_1 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  dirty_40_0 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  dirty_40_1 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  dirty_41_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  dirty_41_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  dirty_42_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  dirty_42_1 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  dirty_43_0 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  dirty_43_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  dirty_44_0 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  dirty_44_1 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  dirty_45_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  dirty_45_1 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  dirty_46_0 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  dirty_46_1 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  dirty_47_0 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  dirty_47_1 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  dirty_48_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  dirty_48_1 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  dirty_49_0 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  dirty_49_1 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  dirty_50_0 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  dirty_50_1 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  dirty_51_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  dirty_51_1 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  dirty_52_0 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  dirty_52_1 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  dirty_53_0 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  dirty_53_1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  dirty_54_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  dirty_54_1 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  dirty_55_0 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  dirty_55_1 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  dirty_56_0 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  dirty_56_1 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  dirty_57_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  dirty_57_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  dirty_58_0 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  dirty_58_1 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  dirty_59_0 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  dirty_59_1 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  dirty_60_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  dirty_60_1 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  dirty_61_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  dirty_61_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  dirty_62_0 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  dirty_62_1 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  dirty_63_0 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  dirty_63_1 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  dirty_64_0 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  dirty_64_1 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  dirty_65_0 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  dirty_65_1 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  dirty_66_0 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  dirty_66_1 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  dirty_67_0 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  dirty_67_1 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  dirty_68_0 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  dirty_68_1 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  dirty_69_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  dirty_69_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  dirty_70_0 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  dirty_70_1 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  dirty_71_0 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  dirty_71_1 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  dirty_72_0 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  dirty_72_1 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  dirty_73_0 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  dirty_73_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  dirty_74_0 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  dirty_74_1 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  dirty_75_0 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  dirty_75_1 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  dirty_76_0 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  dirty_76_1 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  dirty_77_0 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  dirty_77_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  dirty_78_0 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  dirty_78_1 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  dirty_79_0 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  dirty_79_1 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  dirty_80_0 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  dirty_80_1 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  dirty_81_0 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  dirty_81_1 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  dirty_82_0 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  dirty_82_1 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  dirty_83_0 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  dirty_83_1 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  dirty_84_0 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  dirty_84_1 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  dirty_85_0 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  dirty_85_1 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  dirty_86_0 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  dirty_86_1 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  dirty_87_0 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  dirty_87_1 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  dirty_88_0 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  dirty_88_1 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  dirty_89_0 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  dirty_89_1 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  dirty_90_0 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  dirty_90_1 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  dirty_91_0 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  dirty_91_1 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  dirty_92_0 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  dirty_92_1 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  dirty_93_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  dirty_93_1 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  dirty_94_0 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  dirty_94_1 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  dirty_95_0 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  dirty_95_1 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  dirty_96_0 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  dirty_96_1 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  dirty_97_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  dirty_97_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  dirty_98_0 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  dirty_98_1 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  dirty_99_0 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  dirty_99_1 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  dirty_100_0 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  dirty_100_1 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  dirty_101_0 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  dirty_101_1 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  dirty_102_0 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  dirty_102_1 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  dirty_103_0 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  dirty_103_1 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  dirty_104_0 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  dirty_104_1 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  dirty_105_0 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  dirty_105_1 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  dirty_106_0 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  dirty_106_1 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  dirty_107_0 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  dirty_107_1 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  dirty_108_0 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  dirty_108_1 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  dirty_109_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  dirty_109_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  dirty_110_0 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  dirty_110_1 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  dirty_111_0 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  dirty_111_1 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  dirty_112_0 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  dirty_112_1 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  dirty_113_0 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  dirty_113_1 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  dirty_114_0 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  dirty_114_1 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  dirty_115_0 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  dirty_115_1 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  dirty_116_0 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  dirty_116_1 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  dirty_117_0 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  dirty_117_1 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  dirty_118_0 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  dirty_118_1 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  dirty_119_0 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  dirty_119_1 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  dirty_120_0 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  dirty_120_1 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  dirty_121_0 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  dirty_121_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  dirty_122_0 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  dirty_122_1 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  dirty_123_0 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  dirty_123_1 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  dirty_124_0 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  dirty_124_1 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  dirty_125_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  dirty_125_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  dirty_126_0 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  dirty_126_1 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  dirty_127_0 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  dirty_127_1 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  lru_0 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  lru_1 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  lru_2 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  lru_3 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  lru_4 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  lru_5 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  lru_6 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  lru_7 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  lru_8 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  lru_9 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  lru_10 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  lru_11 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  lru_12 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  lru_13 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  lru_14 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  lru_15 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  lru_16 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  lru_17 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  lru_18 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  lru_19 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  lru_20 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  lru_21 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  lru_22 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  lru_23 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  lru_24 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  lru_25 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  lru_26 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  lru_27 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  lru_28 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  lru_29 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  lru_30 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  lru_31 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  lru_32 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  lru_33 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  lru_34 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  lru_35 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  lru_36 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  lru_37 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  lru_38 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  lru_39 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  lru_40 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  lru_41 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  lru_42 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  lru_43 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  lru_44 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  lru_45 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  lru_46 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  lru_47 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  lru_48 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  lru_49 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  lru_50 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  lru_51 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  lru_52 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  lru_53 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  lru_54 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  lru_55 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  lru_56 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  lru_57 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  lru_58 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  lru_59 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  lru_60 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  lru_61 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  lru_62 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  lru_63 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  lru_64 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  lru_65 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  lru_66 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  lru_67 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  lru_68 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  lru_69 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  lru_70 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  lru_71 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  lru_72 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  lru_73 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  lru_74 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  lru_75 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  lru_76 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  lru_77 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  lru_78 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  lru_79 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  lru_80 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  lru_81 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  lru_82 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  lru_83 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  lru_84 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  lru_85 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  lru_86 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  lru_87 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  lru_88 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  lru_89 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  lru_90 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  lru_91 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  lru_92 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  lru_93 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  lru_94 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  lru_95 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  lru_96 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  lru_97 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  lru_98 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  lru_99 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  lru_100 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  lru_101 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  lru_102 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  lru_103 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  lru_104 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  lru_105 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  lru_106 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  lru_107 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  lru_108 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  lru_109 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  lru_110 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  lru_111 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  lru_112 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  lru_113 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  lru_114 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  lru_115 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  lru_116 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  lru_117 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  lru_118 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  lru_119 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  lru_120 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  lru_121 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  lru_122 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  lru_123 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  lru_124 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  lru_125 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  lru_126 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  lru_127 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  tag_wstrb_0 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  tag_wstrb_1 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  bram_replace_wea_0 = _RAND_648[3:0];
  _RAND_649 = {1{`RANDOM}};
  bram_replace_wea_1 = _RAND_649[3:0];
  _RAND_650 = {1{`RANDOM}};
  tag_wdata = _RAND_650[19:0];
  _RAND_651 = {1{`RANDOM}};
  axi_wcnt = _RAND_651[3:0];
  _RAND_652 = {1{`RANDOM}};
  bram_replace_addr = _RAND_652[9:0];
  _RAND_653 = {1{`RANDOM}};
  bram_read_ready_addr = _RAND_653[9:0];
  _RAND_654 = {1{`RANDOM}};
  bram_replace_write_addr = _RAND_654[9:0];
  _RAND_655 = {1{`RANDOM}};
  bram_r_buffer_0 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  bram_r_buffer_1 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  bram_r_buffer_2 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  bram_r_buffer_3 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  bram_r_buffer_4 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  bram_r_buffer_5 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  bram_r_buffer_6 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  bram_r_buffer_7 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  bram_r_buffer_8 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  bram_r_buffer_9 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  bram_r_buffer_10 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  bram_r_buffer_11 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  bram_r_buffer_12 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  bram_r_buffer_13 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  bram_r_buffer_14 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  bram_r_buffer_15 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  bram_use_replace_addr = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  fence_working = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  replace_working = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  ar_handshake = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  aw_handshake = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  replace_writeback = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  saved_rdata = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  last_line_addr = _RAND_678[9:0];
  _RAND_679 = {1{`RANDOM}};
  last_wea_0 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  last_wea_1 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  last_wdata = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  write_buffer_axi_busy = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  ar_addr = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  ar_len = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  ar_size = _RAND_685[2:0];
  _RAND_686 = {1{`RANDOM}};
  arvalid = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  rready = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  aw_addr = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  aw_len = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  aw_size = _RAND_690[2:0];
  _RAND_691 = {1{`RANDOM}};
  awvalid = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  w_data = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  w_strb = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  w_last = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  wvalid = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  current_mmio_write_saved = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  tlb2_vpn = _RAND_697[18:0];
  _RAND_698 = {1{`RANDOM}};
  data_tlb_refill = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  data_tlb_invalid = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  data_tlb_mod = _RAND_700[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheAXIInterface(
  input         clock,
  input         reset,
  output        io_icache_ar_ready,
  input         io_icache_ar_valid,
  input  [31:0] io_icache_ar_bits_addr,
  input  [7:0]  io_icache_ar_bits_len,
  input  [2:0]  io_icache_ar_bits_size,
  input         io_icache_r_ready,
  output        io_icache_r_valid,
  output [31:0] io_icache_r_bits_data,
  output        io_icache_r_bits_last,
  output        io_dcache_ar_ready,
  input         io_dcache_ar_valid,
  input  [31:0] io_dcache_ar_bits_addr,
  input  [7:0]  io_dcache_ar_bits_len,
  input  [2:0]  io_dcache_ar_bits_size,
  input         io_dcache_r_ready,
  output        io_dcache_r_valid,
  output [31:0] io_dcache_r_bits_data,
  output        io_dcache_r_bits_last,
  output        io_dcache_aw_ready,
  input         io_dcache_aw_valid,
  input  [31:0] io_dcache_aw_bits_addr,
  input  [7:0]  io_dcache_aw_bits_len,
  input  [2:0]  io_dcache_aw_bits_size,
  output        io_dcache_w_ready,
  input         io_dcache_w_valid,
  input  [31:0] io_dcache_w_bits_data,
  input  [3:0]  io_dcache_w_bits_strb,
  input         io_dcache_w_bits_last,
  output        io_dcache_b_valid,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [3:0]  io_axi_ar_bits_id,
  output [31:0] io_axi_ar_bits_addr,
  output [7:0]  io_axi_ar_bits_len,
  output [2:0]  io_axi_ar_bits_size,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [3:0]  io_axi_r_bits_id,
  input  [31:0] io_axi_r_bits_data,
  input         io_axi_r_bits_last,
  input         io_axi_aw_ready,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  output [7:0]  io_axi_aw_bits_len,
  output [2:0]  io_axi_aw_bits_size,
  input         io_axi_w_ready,
  output        io_axi_w_valid,
  output [31:0] io_axi_w_bits_data,
  output [3:0]  io_axi_w_bits_strb,
  output        io_axi_w_bits_last,
  input         io_axi_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  ar_sel_lock; // @[CacheAXIInterface.scala 14:32]
  reg  ar_sel_lock_val; // @[CacheAXIInterface.scala 15:32]
  wire  ar_sel = ar_sel_lock ? ar_sel_lock_val : ~io_icache_ar_valid & io_dcache_ar_valid; // @[CacheAXIInterface.scala 25:16]
  wire  r_sel = io_axi_r_bits_id[0]; // @[CacheAXIInterface.scala 26:31]
  wire  _io_icache_r_bits_data_T = ~r_sel; // @[CacheAXIInterface.scala 44:32]
  assign io_icache_ar_ready = io_axi_ar_ready & ~ar_sel; // @[CacheAXIInterface.scala 43:44]
  assign io_icache_r_valid = _io_icache_r_bits_data_T & io_axi_r_valid; // @[CacheAXIInterface.scala 46:31]
  assign io_icache_r_bits_data = ~r_sel ? io_axi_r_bits_data : 32'h0; // @[CacheAXIInterface.scala 44:31]
  assign io_icache_r_bits_last = _io_icache_r_bits_data_T & io_axi_r_bits_last; // @[CacheAXIInterface.scala 45:31]
  assign io_dcache_ar_ready = io_axi_ar_ready & ar_sel; // @[CacheAXIInterface.scala 31:44]
  assign io_dcache_r_valid = r_sel & io_axi_r_valid; // @[CacheAXIInterface.scala 34:31]
  assign io_dcache_r_bits_data = r_sel ? io_axi_r_bits_data : 32'h0; // @[CacheAXIInterface.scala 32:31]
  assign io_dcache_r_bits_last = r_sel & io_axi_r_bits_last; // @[CacheAXIInterface.scala 33:31]
  assign io_dcache_aw_ready = io_axi_aw_ready; // @[CacheAXIInterface.scala 36:22]
  assign io_dcache_w_ready = io_axi_w_ready; // @[CacheAXIInterface.scala 37:22]
  assign io_dcache_b_valid = io_axi_b_valid; // @[CacheAXIInterface.scala 38:22]
  assign io_axi_ar_valid = ar_sel ? io_dcache_ar_valid : io_icache_ar_valid; // @[CacheAXIInterface.scala 59:30]
  assign io_axi_ar_bits_id = {{3'd0}, ar_sel}; // @[CacheAXIInterface.scala 51:24]
  assign io_axi_ar_bits_addr = ar_sel ? io_dcache_ar_bits_addr : io_icache_ar_bits_addr; // @[CacheAXIInterface.scala 52:30]
  assign io_axi_ar_bits_len = ar_sel ? io_dcache_ar_bits_len : io_icache_ar_bits_len; // @[CacheAXIInterface.scala 53:30]
  assign io_axi_ar_bits_size = ar_sel ? io_dcache_ar_bits_size : io_icache_ar_bits_size; // @[CacheAXIInterface.scala 54:30]
  assign io_axi_r_ready = _io_icache_r_bits_data_T ? io_icache_r_ready : io_dcache_r_ready; // @[CacheAXIInterface.scala 61:24]
  assign io_axi_aw_valid = io_dcache_aw_valid; // @[CacheAXIInterface.scala 71:24]
  assign io_axi_aw_bits_addr = io_dcache_aw_bits_addr; // @[CacheAXIInterface.scala 64:24]
  assign io_axi_aw_bits_len = io_dcache_aw_bits_len; // @[CacheAXIInterface.scala 65:24]
  assign io_axi_aw_bits_size = io_dcache_aw_bits_size; // @[CacheAXIInterface.scala 66:24]
  assign io_axi_w_valid = io_dcache_w_valid; // @[CacheAXIInterface.scala 77:22]
  assign io_axi_w_bits_data = io_dcache_w_bits_data; // @[CacheAXIInterface.scala 74:22]
  assign io_axi_w_bits_strb = io_dcache_w_bits_strb; // @[CacheAXIInterface.scala 75:22]
  assign io_axi_w_bits_last = io_dcache_w_bits_last; // @[CacheAXIInterface.scala 76:22]
  always @(posedge clock) begin
    if (reset) begin // @[CacheAXIInterface.scala 14:32]
      ar_sel_lock <= 1'h0; // @[CacheAXIInterface.scala 14:32]
    end else if (io_axi_ar_valid) begin // @[CacheAXIInterface.scala 16:25]
      if (io_axi_ar_ready) begin // @[CacheAXIInterface.scala 17:27]
        ar_sel_lock <= 1'h0; // @[CacheAXIInterface.scala 18:19]
      end else begin
        ar_sel_lock <= 1'h1; // @[CacheAXIInterface.scala 20:23]
      end
    end
    if (reset) begin // @[CacheAXIInterface.scala 15:32]
      ar_sel_lock_val <= 1'h0; // @[CacheAXIInterface.scala 15:32]
    end else if (io_axi_ar_valid) begin // @[CacheAXIInterface.scala 16:25]
      if (!(io_axi_ar_ready)) begin // @[CacheAXIInterface.scala 17:27]
        if (!(ar_sel_lock)) begin // @[CacheAXIInterface.scala 25:16]
          ar_sel_lock_val <= ~io_icache_ar_valid & io_dcache_ar_valid;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ar_sel_lock = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ar_sel_lock_val = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache(
  input         clock,
  input         reset,
  input         io_inst_req,
  input  [31:0] io_inst_addr_0,
  input  [31:0] io_inst_addr_1,
  output [31:0] io_inst_inst_0,
  output [31:0] io_inst_inst_1,
  output        io_inst_inst_valid_0,
  output        io_inst_inst_valid_1,
  input         io_inst_cpu_stall,
  output        io_inst_icache_stall,
  output        io_inst_tlb1_invalid,
  output [18:0] io_inst_tlb2_vpn,
  input         io_inst_tlb2_found,
  input  [19:0] io_inst_tlb2_entry_pfn_0,
  input  [19:0] io_inst_tlb2_entry_pfn_1,
  input         io_inst_tlb2_entry_c_0,
  input         io_inst_tlb2_entry_c_1,
  input         io_inst_tlb2_entry_v_0,
  input         io_inst_tlb2_entry_v_1,
  input         io_inst_fence_value,
  input  [31:0] io_inst_fence_addr,
  input         io_inst_fence_tlb,
  input         io_data_stallM,
  output        io_data_dstall,
  input  [31:0] io_data_E_mem_va,
  input  [31:0] io_data_M_mem_va,
  input  [31:0] io_data_M_fence_addr,
  input         io_data_M_fence_d,
  input         io_data_M_mem_en,
  input         io_data_M_mem_write,
  input  [3:0]  io_data_M_wmask,
  input  [1:0]  io_data_M_mem_size,
  input  [31:0] io_data_M_wdata,
  output [31:0] io_data_M_rdata,
  output [18:0] io_data_tlb_vpn2,
  input         io_data_tlb_found,
  input  [19:0] io_data_tlb_entry_pfn_0,
  input  [19:0] io_data_tlb_entry_pfn_1,
  input         io_data_tlb_entry_c_0,
  input         io_data_tlb_entry_c_1,
  input         io_data_tlb_entry_d_0,
  input         io_data_tlb_entry_d_1,
  input         io_data_tlb_entry_v_0,
  input         io_data_tlb_entry_v_1,
  input         io_data_fence_tlb,
  output        io_data_data_tlb_refill,
  output        io_data_data_tlb_invalid,
  output        io_data_data_tlb_mod,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [3:0]  io_axi_ar_bits_id,
  output [31:0] io_axi_ar_bits_addr,
  output [7:0]  io_axi_ar_bits_len,
  output [2:0]  io_axi_ar_bits_size,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [3:0]  io_axi_r_bits_id,
  input  [31:0] io_axi_r_bits_data,
  input         io_axi_r_bits_last,
  input         io_axi_aw_ready,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  output [7:0]  io_axi_aw_bits_len,
  output [2:0]  io_axi_aw_bits_size,
  input         io_axi_w_ready,
  output        io_axi_w_valid,
  output [31:0] io_axi_w_bits_data,
  output [3:0]  io_axi_w_bits_strb,
  output        io_axi_w_bits_last,
  input         io_axi_b_valid
);
  wire  icache_clock; // @[Cache.scala 17:29]
  wire  icache_reset; // @[Cache.scala 17:29]
  wire  icache_io_cpu_req; // @[Cache.scala 17:29]
  wire [31:0] icache_io_cpu_addr_0; // @[Cache.scala 17:29]
  wire [31:0] icache_io_cpu_addr_1; // @[Cache.scala 17:29]
  wire [31:0] icache_io_cpu_inst_0; // @[Cache.scala 17:29]
  wire [31:0] icache_io_cpu_inst_1; // @[Cache.scala 17:29]
  wire  icache_io_cpu_inst_valid_0; // @[Cache.scala 17:29]
  wire  icache_io_cpu_inst_valid_1; // @[Cache.scala 17:29]
  wire  icache_io_cpu_cpu_stall; // @[Cache.scala 17:29]
  wire  icache_io_cpu_icache_stall; // @[Cache.scala 17:29]
  wire  icache_io_cpu_tlb1_invalid; // @[Cache.scala 17:29]
  wire [18:0] icache_io_cpu_tlb2_vpn; // @[Cache.scala 17:29]
  wire  icache_io_cpu_tlb2_found; // @[Cache.scala 17:29]
  wire [19:0] icache_io_cpu_tlb2_entry_pfn_0; // @[Cache.scala 17:29]
  wire [19:0] icache_io_cpu_tlb2_entry_pfn_1; // @[Cache.scala 17:29]
  wire  icache_io_cpu_tlb2_entry_c_0; // @[Cache.scala 17:29]
  wire  icache_io_cpu_tlb2_entry_c_1; // @[Cache.scala 17:29]
  wire  icache_io_cpu_tlb2_entry_v_0; // @[Cache.scala 17:29]
  wire  icache_io_cpu_tlb2_entry_v_1; // @[Cache.scala 17:29]
  wire  icache_io_cpu_fence_value; // @[Cache.scala 17:29]
  wire [31:0] icache_io_cpu_fence_addr; // @[Cache.scala 17:29]
  wire  icache_io_cpu_fence_tlb; // @[Cache.scala 17:29]
  wire  icache_io_axi_ar_ready; // @[Cache.scala 17:29]
  wire  icache_io_axi_ar_valid; // @[Cache.scala 17:29]
  wire [31:0] icache_io_axi_ar_bits_addr; // @[Cache.scala 17:29]
  wire [7:0] icache_io_axi_ar_bits_len; // @[Cache.scala 17:29]
  wire [2:0] icache_io_axi_ar_bits_size; // @[Cache.scala 17:29]
  wire  icache_io_axi_r_ready; // @[Cache.scala 17:29]
  wire  icache_io_axi_r_valid; // @[Cache.scala 17:29]
  wire [31:0] icache_io_axi_r_bits_data; // @[Cache.scala 17:29]
  wire  icache_io_axi_r_bits_last; // @[Cache.scala 17:29]
  wire  dcache_clock; // @[Cache.scala 18:29]
  wire  dcache_reset; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_stallM; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_dstall; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_cpu_E_mem_va; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_cpu_M_mem_va; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_cpu_M_fence_addr; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_M_fence_d; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_M_mem_en; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_M_mem_write; // @[Cache.scala 18:29]
  wire [3:0] dcache_io_cpu_M_wmask; // @[Cache.scala 18:29]
  wire [1:0] dcache_io_cpu_M_mem_size; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_cpu_M_wdata; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_cpu_M_rdata; // @[Cache.scala 18:29]
  wire [18:0] dcache_io_cpu_tlb_vpn2; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_tlb_found; // @[Cache.scala 18:29]
  wire [19:0] dcache_io_cpu_tlb_entry_pfn_0; // @[Cache.scala 18:29]
  wire [19:0] dcache_io_cpu_tlb_entry_pfn_1; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_tlb_entry_c_0; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_tlb_entry_c_1; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_tlb_entry_d_0; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_tlb_entry_d_1; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_tlb_entry_v_0; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_tlb_entry_v_1; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_fence_tlb; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_data_tlb_refill; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_data_tlb_invalid; // @[Cache.scala 18:29]
  wire  dcache_io_cpu_data_tlb_mod; // @[Cache.scala 18:29]
  wire  dcache_io_axi_ar_ready; // @[Cache.scala 18:29]
  wire  dcache_io_axi_ar_valid; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_axi_ar_bits_addr; // @[Cache.scala 18:29]
  wire [7:0] dcache_io_axi_ar_bits_len; // @[Cache.scala 18:29]
  wire [2:0] dcache_io_axi_ar_bits_size; // @[Cache.scala 18:29]
  wire  dcache_io_axi_r_ready; // @[Cache.scala 18:29]
  wire  dcache_io_axi_r_valid; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_axi_r_bits_data; // @[Cache.scala 18:29]
  wire  dcache_io_axi_r_bits_last; // @[Cache.scala 18:29]
  wire  dcache_io_axi_aw_ready; // @[Cache.scala 18:29]
  wire  dcache_io_axi_aw_valid; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_axi_aw_bits_addr; // @[Cache.scala 18:29]
  wire [7:0] dcache_io_axi_aw_bits_len; // @[Cache.scala 18:29]
  wire [2:0] dcache_io_axi_aw_bits_size; // @[Cache.scala 18:29]
  wire  dcache_io_axi_w_ready; // @[Cache.scala 18:29]
  wire  dcache_io_axi_w_valid; // @[Cache.scala 18:29]
  wire [31:0] dcache_io_axi_w_bits_data; // @[Cache.scala 18:29]
  wire [3:0] dcache_io_axi_w_bits_strb; // @[Cache.scala 18:29]
  wire  dcache_io_axi_w_bits_last; // @[Cache.scala 18:29]
  wire  dcache_io_axi_b_ready; // @[Cache.scala 18:29]
  wire  dcache_io_axi_b_valid; // @[Cache.scala 18:29]
  wire  axi_interface_clock; // @[Cache.scala 19:29]
  wire  axi_interface_reset; // @[Cache.scala 19:29]
  wire  axi_interface_io_icache_ar_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_icache_ar_valid; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_icache_ar_bits_addr; // @[Cache.scala 19:29]
  wire [7:0] axi_interface_io_icache_ar_bits_len; // @[Cache.scala 19:29]
  wire [2:0] axi_interface_io_icache_ar_bits_size; // @[Cache.scala 19:29]
  wire  axi_interface_io_icache_r_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_icache_r_valid; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_icache_r_bits_data; // @[Cache.scala 19:29]
  wire  axi_interface_io_icache_r_bits_last; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_ar_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_ar_valid; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_dcache_ar_bits_addr; // @[Cache.scala 19:29]
  wire [7:0] axi_interface_io_dcache_ar_bits_len; // @[Cache.scala 19:29]
  wire [2:0] axi_interface_io_dcache_ar_bits_size; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_r_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_r_valid; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_dcache_r_bits_data; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_r_bits_last; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_aw_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_aw_valid; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_dcache_aw_bits_addr; // @[Cache.scala 19:29]
  wire [7:0] axi_interface_io_dcache_aw_bits_len; // @[Cache.scala 19:29]
  wire [2:0] axi_interface_io_dcache_aw_bits_size; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_w_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_w_valid; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_dcache_w_bits_data; // @[Cache.scala 19:29]
  wire [3:0] axi_interface_io_dcache_w_bits_strb; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_w_bits_last; // @[Cache.scala 19:29]
  wire  axi_interface_io_dcache_b_valid; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_ar_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_ar_valid; // @[Cache.scala 19:29]
  wire [3:0] axi_interface_io_axi_ar_bits_id; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_axi_ar_bits_addr; // @[Cache.scala 19:29]
  wire [7:0] axi_interface_io_axi_ar_bits_len; // @[Cache.scala 19:29]
  wire [2:0] axi_interface_io_axi_ar_bits_size; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_r_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_r_valid; // @[Cache.scala 19:29]
  wire [3:0] axi_interface_io_axi_r_bits_id; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_axi_r_bits_data; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_r_bits_last; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_aw_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_aw_valid; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_axi_aw_bits_addr; // @[Cache.scala 19:29]
  wire [7:0] axi_interface_io_axi_aw_bits_len; // @[Cache.scala 19:29]
  wire [2:0] axi_interface_io_axi_aw_bits_size; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_w_ready; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_w_valid; // @[Cache.scala 19:29]
  wire [31:0] axi_interface_io_axi_w_bits_data; // @[Cache.scala 19:29]
  wire [3:0] axi_interface_io_axi_w_bits_strb; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_w_bits_last; // @[Cache.scala 19:29]
  wire  axi_interface_io_axi_b_valid; // @[Cache.scala 19:29]
  ICache icache ( // @[Cache.scala 17:29]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_cpu_req(icache_io_cpu_req),
    .io_cpu_addr_0(icache_io_cpu_addr_0),
    .io_cpu_addr_1(icache_io_cpu_addr_1),
    .io_cpu_inst_0(icache_io_cpu_inst_0),
    .io_cpu_inst_1(icache_io_cpu_inst_1),
    .io_cpu_inst_valid_0(icache_io_cpu_inst_valid_0),
    .io_cpu_inst_valid_1(icache_io_cpu_inst_valid_1),
    .io_cpu_cpu_stall(icache_io_cpu_cpu_stall),
    .io_cpu_icache_stall(icache_io_cpu_icache_stall),
    .io_cpu_tlb1_invalid(icache_io_cpu_tlb1_invalid),
    .io_cpu_tlb2_vpn(icache_io_cpu_tlb2_vpn),
    .io_cpu_tlb2_found(icache_io_cpu_tlb2_found),
    .io_cpu_tlb2_entry_pfn_0(icache_io_cpu_tlb2_entry_pfn_0),
    .io_cpu_tlb2_entry_pfn_1(icache_io_cpu_tlb2_entry_pfn_1),
    .io_cpu_tlb2_entry_c_0(icache_io_cpu_tlb2_entry_c_0),
    .io_cpu_tlb2_entry_c_1(icache_io_cpu_tlb2_entry_c_1),
    .io_cpu_tlb2_entry_v_0(icache_io_cpu_tlb2_entry_v_0),
    .io_cpu_tlb2_entry_v_1(icache_io_cpu_tlb2_entry_v_1),
    .io_cpu_fence_value(icache_io_cpu_fence_value),
    .io_cpu_fence_addr(icache_io_cpu_fence_addr),
    .io_cpu_fence_tlb(icache_io_cpu_fence_tlb),
    .io_axi_ar_ready(icache_io_axi_ar_ready),
    .io_axi_ar_valid(icache_io_axi_ar_valid),
    .io_axi_ar_bits_addr(icache_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(icache_io_axi_ar_bits_len),
    .io_axi_ar_bits_size(icache_io_axi_ar_bits_size),
    .io_axi_r_ready(icache_io_axi_r_ready),
    .io_axi_r_valid(icache_io_axi_r_valid),
    .io_axi_r_bits_data(icache_io_axi_r_bits_data),
    .io_axi_r_bits_last(icache_io_axi_r_bits_last)
  );
  DCache dcache ( // @[Cache.scala 18:29]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_cpu_stallM(dcache_io_cpu_stallM),
    .io_cpu_dstall(dcache_io_cpu_dstall),
    .io_cpu_E_mem_va(dcache_io_cpu_E_mem_va),
    .io_cpu_M_mem_va(dcache_io_cpu_M_mem_va),
    .io_cpu_M_fence_addr(dcache_io_cpu_M_fence_addr),
    .io_cpu_M_fence_d(dcache_io_cpu_M_fence_d),
    .io_cpu_M_mem_en(dcache_io_cpu_M_mem_en),
    .io_cpu_M_mem_write(dcache_io_cpu_M_mem_write),
    .io_cpu_M_wmask(dcache_io_cpu_M_wmask),
    .io_cpu_M_mem_size(dcache_io_cpu_M_mem_size),
    .io_cpu_M_wdata(dcache_io_cpu_M_wdata),
    .io_cpu_M_rdata(dcache_io_cpu_M_rdata),
    .io_cpu_tlb_vpn2(dcache_io_cpu_tlb_vpn2),
    .io_cpu_tlb_found(dcache_io_cpu_tlb_found),
    .io_cpu_tlb_entry_pfn_0(dcache_io_cpu_tlb_entry_pfn_0),
    .io_cpu_tlb_entry_pfn_1(dcache_io_cpu_tlb_entry_pfn_1),
    .io_cpu_tlb_entry_c_0(dcache_io_cpu_tlb_entry_c_0),
    .io_cpu_tlb_entry_c_1(dcache_io_cpu_tlb_entry_c_1),
    .io_cpu_tlb_entry_d_0(dcache_io_cpu_tlb_entry_d_0),
    .io_cpu_tlb_entry_d_1(dcache_io_cpu_tlb_entry_d_1),
    .io_cpu_tlb_entry_v_0(dcache_io_cpu_tlb_entry_v_0),
    .io_cpu_tlb_entry_v_1(dcache_io_cpu_tlb_entry_v_1),
    .io_cpu_fence_tlb(dcache_io_cpu_fence_tlb),
    .io_cpu_data_tlb_refill(dcache_io_cpu_data_tlb_refill),
    .io_cpu_data_tlb_invalid(dcache_io_cpu_data_tlb_invalid),
    .io_cpu_data_tlb_mod(dcache_io_cpu_data_tlb_mod),
    .io_axi_ar_ready(dcache_io_axi_ar_ready),
    .io_axi_ar_valid(dcache_io_axi_ar_valid),
    .io_axi_ar_bits_addr(dcache_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(dcache_io_axi_ar_bits_len),
    .io_axi_ar_bits_size(dcache_io_axi_ar_bits_size),
    .io_axi_r_ready(dcache_io_axi_r_ready),
    .io_axi_r_valid(dcache_io_axi_r_valid),
    .io_axi_r_bits_data(dcache_io_axi_r_bits_data),
    .io_axi_r_bits_last(dcache_io_axi_r_bits_last),
    .io_axi_aw_ready(dcache_io_axi_aw_ready),
    .io_axi_aw_valid(dcache_io_axi_aw_valid),
    .io_axi_aw_bits_addr(dcache_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(dcache_io_axi_aw_bits_len),
    .io_axi_aw_bits_size(dcache_io_axi_aw_bits_size),
    .io_axi_w_ready(dcache_io_axi_w_ready),
    .io_axi_w_valid(dcache_io_axi_w_valid),
    .io_axi_w_bits_data(dcache_io_axi_w_bits_data),
    .io_axi_w_bits_strb(dcache_io_axi_w_bits_strb),
    .io_axi_w_bits_last(dcache_io_axi_w_bits_last),
    .io_axi_b_ready(dcache_io_axi_b_ready),
    .io_axi_b_valid(dcache_io_axi_b_valid)
  );
  CacheAXIInterface axi_interface ( // @[Cache.scala 19:29]
    .clock(axi_interface_clock),
    .reset(axi_interface_reset),
    .io_icache_ar_ready(axi_interface_io_icache_ar_ready),
    .io_icache_ar_valid(axi_interface_io_icache_ar_valid),
    .io_icache_ar_bits_addr(axi_interface_io_icache_ar_bits_addr),
    .io_icache_ar_bits_len(axi_interface_io_icache_ar_bits_len),
    .io_icache_ar_bits_size(axi_interface_io_icache_ar_bits_size),
    .io_icache_r_ready(axi_interface_io_icache_r_ready),
    .io_icache_r_valid(axi_interface_io_icache_r_valid),
    .io_icache_r_bits_data(axi_interface_io_icache_r_bits_data),
    .io_icache_r_bits_last(axi_interface_io_icache_r_bits_last),
    .io_dcache_ar_ready(axi_interface_io_dcache_ar_ready),
    .io_dcache_ar_valid(axi_interface_io_dcache_ar_valid),
    .io_dcache_ar_bits_addr(axi_interface_io_dcache_ar_bits_addr),
    .io_dcache_ar_bits_len(axi_interface_io_dcache_ar_bits_len),
    .io_dcache_ar_bits_size(axi_interface_io_dcache_ar_bits_size),
    .io_dcache_r_ready(axi_interface_io_dcache_r_ready),
    .io_dcache_r_valid(axi_interface_io_dcache_r_valid),
    .io_dcache_r_bits_data(axi_interface_io_dcache_r_bits_data),
    .io_dcache_r_bits_last(axi_interface_io_dcache_r_bits_last),
    .io_dcache_aw_ready(axi_interface_io_dcache_aw_ready),
    .io_dcache_aw_valid(axi_interface_io_dcache_aw_valid),
    .io_dcache_aw_bits_addr(axi_interface_io_dcache_aw_bits_addr),
    .io_dcache_aw_bits_len(axi_interface_io_dcache_aw_bits_len),
    .io_dcache_aw_bits_size(axi_interface_io_dcache_aw_bits_size),
    .io_dcache_w_ready(axi_interface_io_dcache_w_ready),
    .io_dcache_w_valid(axi_interface_io_dcache_w_valid),
    .io_dcache_w_bits_data(axi_interface_io_dcache_w_bits_data),
    .io_dcache_w_bits_strb(axi_interface_io_dcache_w_bits_strb),
    .io_dcache_w_bits_last(axi_interface_io_dcache_w_bits_last),
    .io_dcache_b_valid(axi_interface_io_dcache_b_valid),
    .io_axi_ar_ready(axi_interface_io_axi_ar_ready),
    .io_axi_ar_valid(axi_interface_io_axi_ar_valid),
    .io_axi_ar_bits_id(axi_interface_io_axi_ar_bits_id),
    .io_axi_ar_bits_addr(axi_interface_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(axi_interface_io_axi_ar_bits_len),
    .io_axi_ar_bits_size(axi_interface_io_axi_ar_bits_size),
    .io_axi_r_ready(axi_interface_io_axi_r_ready),
    .io_axi_r_valid(axi_interface_io_axi_r_valid),
    .io_axi_r_bits_id(axi_interface_io_axi_r_bits_id),
    .io_axi_r_bits_data(axi_interface_io_axi_r_bits_data),
    .io_axi_r_bits_last(axi_interface_io_axi_r_bits_last),
    .io_axi_aw_ready(axi_interface_io_axi_aw_ready),
    .io_axi_aw_valid(axi_interface_io_axi_aw_valid),
    .io_axi_aw_bits_addr(axi_interface_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(axi_interface_io_axi_aw_bits_len),
    .io_axi_aw_bits_size(axi_interface_io_axi_aw_bits_size),
    .io_axi_w_ready(axi_interface_io_axi_w_ready),
    .io_axi_w_valid(axi_interface_io_axi_w_valid),
    .io_axi_w_bits_data(axi_interface_io_axi_w_bits_data),
    .io_axi_w_bits_strb(axi_interface_io_axi_w_bits_strb),
    .io_axi_w_bits_last(axi_interface_io_axi_w_bits_last),
    .io_axi_b_valid(axi_interface_io_axi_b_valid)
  );
  assign io_inst_inst_0 = icache_io_cpu_inst_0; // @[Cache.scala 24:11]
  assign io_inst_inst_1 = icache_io_cpu_inst_1; // @[Cache.scala 24:11]
  assign io_inst_inst_valid_0 = icache_io_cpu_inst_valid_0; // @[Cache.scala 24:11]
  assign io_inst_inst_valid_1 = icache_io_cpu_inst_valid_1; // @[Cache.scala 24:11]
  assign io_inst_icache_stall = icache_io_cpu_icache_stall; // @[Cache.scala 24:11]
  assign io_inst_tlb1_invalid = icache_io_cpu_tlb1_invalid; // @[Cache.scala 24:11]
  assign io_inst_tlb2_vpn = icache_io_cpu_tlb2_vpn; // @[Cache.scala 24:11]
  assign io_data_dstall = dcache_io_cpu_dstall; // @[Cache.scala 25:11]
  assign io_data_M_rdata = dcache_io_cpu_M_rdata; // @[Cache.scala 25:11]
  assign io_data_tlb_vpn2 = dcache_io_cpu_tlb_vpn2; // @[Cache.scala 25:11]
  assign io_data_data_tlb_refill = dcache_io_cpu_data_tlb_refill; // @[Cache.scala 25:11]
  assign io_data_data_tlb_invalid = dcache_io_cpu_data_tlb_invalid; // @[Cache.scala 25:11]
  assign io_data_data_tlb_mod = dcache_io_cpu_data_tlb_mod; // @[Cache.scala 25:11]
  assign io_axi_ar_valid = axi_interface_io_axi_ar_valid; // @[Cache.scala 26:10]
  assign io_axi_ar_bits_id = axi_interface_io_axi_ar_bits_id; // @[Cache.scala 26:10]
  assign io_axi_ar_bits_addr = axi_interface_io_axi_ar_bits_addr; // @[Cache.scala 26:10]
  assign io_axi_ar_bits_len = axi_interface_io_axi_ar_bits_len; // @[Cache.scala 26:10]
  assign io_axi_ar_bits_size = axi_interface_io_axi_ar_bits_size; // @[Cache.scala 26:10]
  assign io_axi_r_ready = axi_interface_io_axi_r_ready; // @[Cache.scala 26:10]
  assign io_axi_aw_valid = axi_interface_io_axi_aw_valid; // @[Cache.scala 26:10]
  assign io_axi_aw_bits_addr = axi_interface_io_axi_aw_bits_addr; // @[Cache.scala 26:10]
  assign io_axi_aw_bits_len = axi_interface_io_axi_aw_bits_len; // @[Cache.scala 26:10]
  assign io_axi_aw_bits_size = axi_interface_io_axi_aw_bits_size; // @[Cache.scala 26:10]
  assign io_axi_w_valid = axi_interface_io_axi_w_valid; // @[Cache.scala 26:10]
  assign io_axi_w_bits_data = axi_interface_io_axi_w_bits_data; // @[Cache.scala 26:10]
  assign io_axi_w_bits_strb = axi_interface_io_axi_w_bits_strb; // @[Cache.scala 26:10]
  assign io_axi_w_bits_last = axi_interface_io_axi_w_bits_last; // @[Cache.scala 26:10]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_cpu_req = io_inst_req; // @[Cache.scala 24:11]
  assign icache_io_cpu_addr_0 = io_inst_addr_0; // @[Cache.scala 24:11]
  assign icache_io_cpu_addr_1 = io_inst_addr_1; // @[Cache.scala 24:11]
  assign icache_io_cpu_cpu_stall = io_inst_cpu_stall; // @[Cache.scala 24:11]
  assign icache_io_cpu_tlb2_found = io_inst_tlb2_found; // @[Cache.scala 24:11]
  assign icache_io_cpu_tlb2_entry_pfn_0 = io_inst_tlb2_entry_pfn_0; // @[Cache.scala 24:11]
  assign icache_io_cpu_tlb2_entry_pfn_1 = io_inst_tlb2_entry_pfn_1; // @[Cache.scala 24:11]
  assign icache_io_cpu_tlb2_entry_c_0 = io_inst_tlb2_entry_c_0; // @[Cache.scala 24:11]
  assign icache_io_cpu_tlb2_entry_c_1 = io_inst_tlb2_entry_c_1; // @[Cache.scala 24:11]
  assign icache_io_cpu_tlb2_entry_v_0 = io_inst_tlb2_entry_v_0; // @[Cache.scala 24:11]
  assign icache_io_cpu_tlb2_entry_v_1 = io_inst_tlb2_entry_v_1; // @[Cache.scala 24:11]
  assign icache_io_cpu_fence_value = io_inst_fence_value; // @[Cache.scala 24:11]
  assign icache_io_cpu_fence_addr = io_inst_fence_addr; // @[Cache.scala 24:11]
  assign icache_io_cpu_fence_tlb = io_inst_fence_tlb; // @[Cache.scala 24:11]
  assign icache_io_axi_ar_ready = axi_interface_io_icache_ar_ready; // @[Cache.scala 21:17]
  assign icache_io_axi_r_valid = axi_interface_io_icache_r_valid; // @[Cache.scala 21:17]
  assign icache_io_axi_r_bits_data = axi_interface_io_icache_r_bits_data; // @[Cache.scala 21:17]
  assign icache_io_axi_r_bits_last = axi_interface_io_icache_r_bits_last; // @[Cache.scala 21:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_cpu_stallM = io_data_stallM; // @[Cache.scala 25:11]
  assign dcache_io_cpu_E_mem_va = io_data_E_mem_va; // @[Cache.scala 25:11]
  assign dcache_io_cpu_M_mem_va = io_data_M_mem_va; // @[Cache.scala 25:11]
  assign dcache_io_cpu_M_fence_addr = io_data_M_fence_addr; // @[Cache.scala 25:11]
  assign dcache_io_cpu_M_fence_d = io_data_M_fence_d; // @[Cache.scala 25:11]
  assign dcache_io_cpu_M_mem_en = io_data_M_mem_en; // @[Cache.scala 25:11]
  assign dcache_io_cpu_M_mem_write = io_data_M_mem_write; // @[Cache.scala 25:11]
  assign dcache_io_cpu_M_wmask = io_data_M_wmask; // @[Cache.scala 25:11]
  assign dcache_io_cpu_M_mem_size = io_data_M_mem_size; // @[Cache.scala 25:11]
  assign dcache_io_cpu_M_wdata = io_data_M_wdata; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_found = io_data_tlb_found; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_entry_pfn_0 = io_data_tlb_entry_pfn_0; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_entry_pfn_1 = io_data_tlb_entry_pfn_1; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_entry_c_0 = io_data_tlb_entry_c_0; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_entry_c_1 = io_data_tlb_entry_c_1; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_entry_d_0 = io_data_tlb_entry_d_0; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_entry_d_1 = io_data_tlb_entry_d_1; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_entry_v_0 = io_data_tlb_entry_v_0; // @[Cache.scala 25:11]
  assign dcache_io_cpu_tlb_entry_v_1 = io_data_tlb_entry_v_1; // @[Cache.scala 25:11]
  assign dcache_io_cpu_fence_tlb = io_data_fence_tlb; // @[Cache.scala 25:11]
  assign dcache_io_axi_ar_ready = axi_interface_io_dcache_ar_ready; // @[Cache.scala 22:17]
  assign dcache_io_axi_r_valid = axi_interface_io_dcache_r_valid; // @[Cache.scala 22:17]
  assign dcache_io_axi_r_bits_data = axi_interface_io_dcache_r_bits_data; // @[Cache.scala 22:17]
  assign dcache_io_axi_r_bits_last = axi_interface_io_dcache_r_bits_last; // @[Cache.scala 22:17]
  assign dcache_io_axi_aw_ready = axi_interface_io_dcache_aw_ready; // @[Cache.scala 22:17]
  assign dcache_io_axi_w_ready = axi_interface_io_dcache_w_ready; // @[Cache.scala 22:17]
  assign dcache_io_axi_b_valid = axi_interface_io_dcache_b_valid; // @[Cache.scala 22:17]
  assign axi_interface_clock = clock;
  assign axi_interface_reset = reset;
  assign axi_interface_io_icache_ar_valid = icache_io_axi_ar_valid; // @[Cache.scala 21:17]
  assign axi_interface_io_icache_ar_bits_addr = icache_io_axi_ar_bits_addr; // @[Cache.scala 21:17]
  assign axi_interface_io_icache_ar_bits_len = icache_io_axi_ar_bits_len; // @[Cache.scala 21:17]
  assign axi_interface_io_icache_ar_bits_size = icache_io_axi_ar_bits_size; // @[Cache.scala 21:17]
  assign axi_interface_io_icache_r_ready = icache_io_axi_r_ready; // @[Cache.scala 21:17]
  assign axi_interface_io_dcache_ar_valid = dcache_io_axi_ar_valid; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_ar_bits_addr = dcache_io_axi_ar_bits_addr; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_ar_bits_len = dcache_io_axi_ar_bits_len; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_ar_bits_size = dcache_io_axi_ar_bits_size; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_r_ready = dcache_io_axi_r_ready; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_aw_valid = dcache_io_axi_aw_valid; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_aw_bits_addr = dcache_io_axi_aw_bits_addr; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_aw_bits_len = dcache_io_axi_aw_bits_len; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_aw_bits_size = dcache_io_axi_aw_bits_size; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_w_valid = dcache_io_axi_w_valid; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_w_bits_data = dcache_io_axi_w_bits_data; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_w_bits_strb = dcache_io_axi_w_bits_strb; // @[Cache.scala 22:17]
  assign axi_interface_io_dcache_w_bits_last = dcache_io_axi_w_bits_last; // @[Cache.scala 22:17]
  assign axi_interface_io_axi_ar_ready = io_axi_ar_ready; // @[Cache.scala 26:10]
  assign axi_interface_io_axi_r_valid = io_axi_r_valid; // @[Cache.scala 26:10]
  assign axi_interface_io_axi_r_bits_id = io_axi_r_bits_id; // @[Cache.scala 26:10]
  assign axi_interface_io_axi_r_bits_data = io_axi_r_bits_data; // @[Cache.scala 26:10]
  assign axi_interface_io_axi_r_bits_last = io_axi_r_bits_last; // @[Cache.scala 26:10]
  assign axi_interface_io_axi_aw_ready = io_axi_aw_ready; // @[Cache.scala 26:10]
  assign axi_interface_io_axi_w_ready = io_axi_w_ready; // @[Cache.scala 26:10]
  assign axi_interface_io_axi_b_valid = io_axi_b_valid; // @[Cache.scala 26:10]
endmodule
module PuaMips(
  input         clock,
  input         reset,
  input  [5:0]  io_ext_int,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [3:0]  io_axi_ar_bits_id,
  output [31:0] io_axi_ar_bits_addr,
  output [7:0]  io_axi_ar_bits_len,
  output [2:0]  io_axi_ar_bits_size,
  output [1:0]  io_axi_ar_bits_burst,
  output [1:0]  io_axi_ar_bits_lock,
  output [3:0]  io_axi_ar_bits_cache,
  output [2:0]  io_axi_ar_bits_prot,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [3:0]  io_axi_r_bits_id,
  input  [31:0] io_axi_r_bits_data,
  input  [1:0]  io_axi_r_bits_resp,
  input         io_axi_r_bits_last,
  input         io_axi_aw_ready,
  output        io_axi_aw_valid,
  output [3:0]  io_axi_aw_bits_id,
  output [31:0] io_axi_aw_bits_addr,
  output [7:0]  io_axi_aw_bits_len,
  output [2:0]  io_axi_aw_bits_size,
  output [1:0]  io_axi_aw_bits_burst,
  output [1:0]  io_axi_aw_bits_lock,
  output [3:0]  io_axi_aw_bits_cache,
  output [2:0]  io_axi_aw_bits_prot,
  input         io_axi_w_ready,
  output        io_axi_w_valid,
  output [3:0]  io_axi_w_bits_id,
  output [31:0] io_axi_w_bits_data,
  output [3:0]  io_axi_w_bits_strb,
  output        io_axi_w_bits_last,
  output        io_axi_b_ready,
  input         io_axi_b_valid,
  input  [3:0]  io_axi_b_bits_id,
  input  [1:0]  io_axi_b_bits_resp,
  output [31:0] io_debug_wb_pc,
  output [3:0]  io_debug_wb_rf_wen,
  output [4:0]  io_debug_wb_rf_wnum,
  output [31:0] io_debug_wb_rf_wdata,
  output [31:0] io_debug_cp0_count,
  output [31:0] io_debug_cp0_random,
  output [31:0] io_debug_cp0_cause,
  output        io_debug_int,
  output        io_debug_commit
);
  wire  core_clock; // @[PuaMips.scala 14:21]
  wire  core_reset; // @[PuaMips.scala 14:21]
  wire [5:0] core_io_ext_int; // @[PuaMips.scala 14:21]
  wire  core_io_inst_req; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_inst_addr_0; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_inst_addr_1; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_inst_inst_0; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_inst_inst_1; // @[PuaMips.scala 14:21]
  wire  core_io_inst_inst_valid_0; // @[PuaMips.scala 14:21]
  wire  core_io_inst_inst_valid_1; // @[PuaMips.scala 14:21]
  wire  core_io_inst_cpu_stall; // @[PuaMips.scala 14:21]
  wire  core_io_inst_icache_stall; // @[PuaMips.scala 14:21]
  wire  core_io_inst_tlb1_invalid; // @[PuaMips.scala 14:21]
  wire [18:0] core_io_inst_tlb2_vpn; // @[PuaMips.scala 14:21]
  wire  core_io_inst_tlb2_found; // @[PuaMips.scala 14:21]
  wire [19:0] core_io_inst_tlb2_entry_pfn_0; // @[PuaMips.scala 14:21]
  wire [19:0] core_io_inst_tlb2_entry_pfn_1; // @[PuaMips.scala 14:21]
  wire  core_io_inst_tlb2_entry_c_0; // @[PuaMips.scala 14:21]
  wire  core_io_inst_tlb2_entry_c_1; // @[PuaMips.scala 14:21]
  wire  core_io_inst_tlb2_entry_v_0; // @[PuaMips.scala 14:21]
  wire  core_io_inst_tlb2_entry_v_1; // @[PuaMips.scala 14:21]
  wire  core_io_inst_fence_value; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_inst_fence_addr; // @[PuaMips.scala 14:21]
  wire  core_io_inst_fence_tlb; // @[PuaMips.scala 14:21]
  wire  core_io_data_stallM; // @[PuaMips.scala 14:21]
  wire  core_io_data_dstall; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_data_E_mem_va; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_data_M_mem_va; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_data_M_fence_addr; // @[PuaMips.scala 14:21]
  wire  core_io_data_M_fence_d; // @[PuaMips.scala 14:21]
  wire  core_io_data_M_mem_en; // @[PuaMips.scala 14:21]
  wire  core_io_data_M_mem_write; // @[PuaMips.scala 14:21]
  wire [3:0] core_io_data_M_wmask; // @[PuaMips.scala 14:21]
  wire [1:0] core_io_data_M_mem_size; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_data_M_wdata; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_data_M_rdata; // @[PuaMips.scala 14:21]
  wire [18:0] core_io_data_tlb_vpn2; // @[PuaMips.scala 14:21]
  wire  core_io_data_tlb_found; // @[PuaMips.scala 14:21]
  wire [19:0] core_io_data_tlb_entry_pfn_0; // @[PuaMips.scala 14:21]
  wire [19:0] core_io_data_tlb_entry_pfn_1; // @[PuaMips.scala 14:21]
  wire  core_io_data_tlb_entry_c_0; // @[PuaMips.scala 14:21]
  wire  core_io_data_tlb_entry_c_1; // @[PuaMips.scala 14:21]
  wire  core_io_data_tlb_entry_d_0; // @[PuaMips.scala 14:21]
  wire  core_io_data_tlb_entry_d_1; // @[PuaMips.scala 14:21]
  wire  core_io_data_tlb_entry_v_0; // @[PuaMips.scala 14:21]
  wire  core_io_data_tlb_entry_v_1; // @[PuaMips.scala 14:21]
  wire  core_io_data_fence_tlb; // @[PuaMips.scala 14:21]
  wire  core_io_data_data_tlb_refill; // @[PuaMips.scala 14:21]
  wire  core_io_data_data_tlb_invalid; // @[PuaMips.scala 14:21]
  wire  core_io_data_data_tlb_mod; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_debug_wb_pc; // @[PuaMips.scala 14:21]
  wire [3:0] core_io_debug_wb_rf_wen; // @[PuaMips.scala 14:21]
  wire [4:0] core_io_debug_wb_rf_wnum; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_debug_wb_rf_wdata; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_debug_cp0_count; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_debug_cp0_random; // @[PuaMips.scala 14:21]
  wire [31:0] core_io_debug_cp0_cause; // @[PuaMips.scala 14:21]
  wire  core_io_debug_int; // @[PuaMips.scala 14:21]
  wire  core_io_debug_commit; // @[PuaMips.scala 14:21]
  wire  cache_clock; // @[PuaMips.scala 15:21]
  wire  cache_reset; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_req; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_inst_addr_0; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_inst_addr_1; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_inst_inst_0; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_inst_inst_1; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_inst_valid_0; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_inst_valid_1; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_cpu_stall; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_icache_stall; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_tlb1_invalid; // @[PuaMips.scala 15:21]
  wire [18:0] cache_io_inst_tlb2_vpn; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_tlb2_found; // @[PuaMips.scala 15:21]
  wire [19:0] cache_io_inst_tlb2_entry_pfn_0; // @[PuaMips.scala 15:21]
  wire [19:0] cache_io_inst_tlb2_entry_pfn_1; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_tlb2_entry_c_0; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_tlb2_entry_c_1; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_tlb2_entry_v_0; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_tlb2_entry_v_1; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_fence_value; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_inst_fence_addr; // @[PuaMips.scala 15:21]
  wire  cache_io_inst_fence_tlb; // @[PuaMips.scala 15:21]
  wire  cache_io_data_stallM; // @[PuaMips.scala 15:21]
  wire  cache_io_data_dstall; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_data_E_mem_va; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_data_M_mem_va; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_data_M_fence_addr; // @[PuaMips.scala 15:21]
  wire  cache_io_data_M_fence_d; // @[PuaMips.scala 15:21]
  wire  cache_io_data_M_mem_en; // @[PuaMips.scala 15:21]
  wire  cache_io_data_M_mem_write; // @[PuaMips.scala 15:21]
  wire [3:0] cache_io_data_M_wmask; // @[PuaMips.scala 15:21]
  wire [1:0] cache_io_data_M_mem_size; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_data_M_wdata; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_data_M_rdata; // @[PuaMips.scala 15:21]
  wire [18:0] cache_io_data_tlb_vpn2; // @[PuaMips.scala 15:21]
  wire  cache_io_data_tlb_found; // @[PuaMips.scala 15:21]
  wire [19:0] cache_io_data_tlb_entry_pfn_0; // @[PuaMips.scala 15:21]
  wire [19:0] cache_io_data_tlb_entry_pfn_1; // @[PuaMips.scala 15:21]
  wire  cache_io_data_tlb_entry_c_0; // @[PuaMips.scala 15:21]
  wire  cache_io_data_tlb_entry_c_1; // @[PuaMips.scala 15:21]
  wire  cache_io_data_tlb_entry_d_0; // @[PuaMips.scala 15:21]
  wire  cache_io_data_tlb_entry_d_1; // @[PuaMips.scala 15:21]
  wire  cache_io_data_tlb_entry_v_0; // @[PuaMips.scala 15:21]
  wire  cache_io_data_tlb_entry_v_1; // @[PuaMips.scala 15:21]
  wire  cache_io_data_fence_tlb; // @[PuaMips.scala 15:21]
  wire  cache_io_data_data_tlb_refill; // @[PuaMips.scala 15:21]
  wire  cache_io_data_data_tlb_invalid; // @[PuaMips.scala 15:21]
  wire  cache_io_data_data_tlb_mod; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_ar_ready; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_ar_valid; // @[PuaMips.scala 15:21]
  wire [3:0] cache_io_axi_ar_bits_id; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_axi_ar_bits_addr; // @[PuaMips.scala 15:21]
  wire [7:0] cache_io_axi_ar_bits_len; // @[PuaMips.scala 15:21]
  wire [2:0] cache_io_axi_ar_bits_size; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_r_ready; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_r_valid; // @[PuaMips.scala 15:21]
  wire [3:0] cache_io_axi_r_bits_id; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_axi_r_bits_data; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_r_bits_last; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_aw_ready; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_aw_valid; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_axi_aw_bits_addr; // @[PuaMips.scala 15:21]
  wire [7:0] cache_io_axi_aw_bits_len; // @[PuaMips.scala 15:21]
  wire [2:0] cache_io_axi_aw_bits_size; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_w_ready; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_w_valid; // @[PuaMips.scala 15:21]
  wire [31:0] cache_io_axi_w_bits_data; // @[PuaMips.scala 15:21]
  wire [3:0] cache_io_axi_w_bits_strb; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_w_bits_last; // @[PuaMips.scala 15:21]
  wire  cache_io_axi_b_valid; // @[PuaMips.scala 15:21]
  Core core ( // @[PuaMips.scala 14:21]
    .clock(core_clock),
    .reset(core_reset),
    .io_ext_int(core_io_ext_int),
    .io_inst_req(core_io_inst_req),
    .io_inst_addr_0(core_io_inst_addr_0),
    .io_inst_addr_1(core_io_inst_addr_1),
    .io_inst_inst_0(core_io_inst_inst_0),
    .io_inst_inst_1(core_io_inst_inst_1),
    .io_inst_inst_valid_0(core_io_inst_inst_valid_0),
    .io_inst_inst_valid_1(core_io_inst_inst_valid_1),
    .io_inst_cpu_stall(core_io_inst_cpu_stall),
    .io_inst_icache_stall(core_io_inst_icache_stall),
    .io_inst_tlb1_invalid(core_io_inst_tlb1_invalid),
    .io_inst_tlb2_vpn(core_io_inst_tlb2_vpn),
    .io_inst_tlb2_found(core_io_inst_tlb2_found),
    .io_inst_tlb2_entry_pfn_0(core_io_inst_tlb2_entry_pfn_0),
    .io_inst_tlb2_entry_pfn_1(core_io_inst_tlb2_entry_pfn_1),
    .io_inst_tlb2_entry_c_0(core_io_inst_tlb2_entry_c_0),
    .io_inst_tlb2_entry_c_1(core_io_inst_tlb2_entry_c_1),
    .io_inst_tlb2_entry_v_0(core_io_inst_tlb2_entry_v_0),
    .io_inst_tlb2_entry_v_1(core_io_inst_tlb2_entry_v_1),
    .io_inst_fence_value(core_io_inst_fence_value),
    .io_inst_fence_addr(core_io_inst_fence_addr),
    .io_inst_fence_tlb(core_io_inst_fence_tlb),
    .io_data_stallM(core_io_data_stallM),
    .io_data_dstall(core_io_data_dstall),
    .io_data_E_mem_va(core_io_data_E_mem_va),
    .io_data_M_mem_va(core_io_data_M_mem_va),
    .io_data_M_fence_addr(core_io_data_M_fence_addr),
    .io_data_M_fence_d(core_io_data_M_fence_d),
    .io_data_M_mem_en(core_io_data_M_mem_en),
    .io_data_M_mem_write(core_io_data_M_mem_write),
    .io_data_M_wmask(core_io_data_M_wmask),
    .io_data_M_mem_size(core_io_data_M_mem_size),
    .io_data_M_wdata(core_io_data_M_wdata),
    .io_data_M_rdata(core_io_data_M_rdata),
    .io_data_tlb_vpn2(core_io_data_tlb_vpn2),
    .io_data_tlb_found(core_io_data_tlb_found),
    .io_data_tlb_entry_pfn_0(core_io_data_tlb_entry_pfn_0),
    .io_data_tlb_entry_pfn_1(core_io_data_tlb_entry_pfn_1),
    .io_data_tlb_entry_c_0(core_io_data_tlb_entry_c_0),
    .io_data_tlb_entry_c_1(core_io_data_tlb_entry_c_1),
    .io_data_tlb_entry_d_0(core_io_data_tlb_entry_d_0),
    .io_data_tlb_entry_d_1(core_io_data_tlb_entry_d_1),
    .io_data_tlb_entry_v_0(core_io_data_tlb_entry_v_0),
    .io_data_tlb_entry_v_1(core_io_data_tlb_entry_v_1),
    .io_data_fence_tlb(core_io_data_fence_tlb),
    .io_data_data_tlb_refill(core_io_data_data_tlb_refill),
    .io_data_data_tlb_invalid(core_io_data_data_tlb_invalid),
    .io_data_data_tlb_mod(core_io_data_data_tlb_mod),
    .io_debug_wb_pc(core_io_debug_wb_pc),
    .io_debug_wb_rf_wen(core_io_debug_wb_rf_wen),
    .io_debug_wb_rf_wnum(core_io_debug_wb_rf_wnum),
    .io_debug_wb_rf_wdata(core_io_debug_wb_rf_wdata),
    .io_debug_cp0_count(core_io_debug_cp0_count),
    .io_debug_cp0_random(core_io_debug_cp0_random),
    .io_debug_cp0_cause(core_io_debug_cp0_cause),
    .io_debug_int(core_io_debug_int),
    .io_debug_commit(core_io_debug_commit)
  );
  Cache cache ( // @[PuaMips.scala 15:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_inst_req(cache_io_inst_req),
    .io_inst_addr_0(cache_io_inst_addr_0),
    .io_inst_addr_1(cache_io_inst_addr_1),
    .io_inst_inst_0(cache_io_inst_inst_0),
    .io_inst_inst_1(cache_io_inst_inst_1),
    .io_inst_inst_valid_0(cache_io_inst_inst_valid_0),
    .io_inst_inst_valid_1(cache_io_inst_inst_valid_1),
    .io_inst_cpu_stall(cache_io_inst_cpu_stall),
    .io_inst_icache_stall(cache_io_inst_icache_stall),
    .io_inst_tlb1_invalid(cache_io_inst_tlb1_invalid),
    .io_inst_tlb2_vpn(cache_io_inst_tlb2_vpn),
    .io_inst_tlb2_found(cache_io_inst_tlb2_found),
    .io_inst_tlb2_entry_pfn_0(cache_io_inst_tlb2_entry_pfn_0),
    .io_inst_tlb2_entry_pfn_1(cache_io_inst_tlb2_entry_pfn_1),
    .io_inst_tlb2_entry_c_0(cache_io_inst_tlb2_entry_c_0),
    .io_inst_tlb2_entry_c_1(cache_io_inst_tlb2_entry_c_1),
    .io_inst_tlb2_entry_v_0(cache_io_inst_tlb2_entry_v_0),
    .io_inst_tlb2_entry_v_1(cache_io_inst_tlb2_entry_v_1),
    .io_inst_fence_value(cache_io_inst_fence_value),
    .io_inst_fence_addr(cache_io_inst_fence_addr),
    .io_inst_fence_tlb(cache_io_inst_fence_tlb),
    .io_data_stallM(cache_io_data_stallM),
    .io_data_dstall(cache_io_data_dstall),
    .io_data_E_mem_va(cache_io_data_E_mem_va),
    .io_data_M_mem_va(cache_io_data_M_mem_va),
    .io_data_M_fence_addr(cache_io_data_M_fence_addr),
    .io_data_M_fence_d(cache_io_data_M_fence_d),
    .io_data_M_mem_en(cache_io_data_M_mem_en),
    .io_data_M_mem_write(cache_io_data_M_mem_write),
    .io_data_M_wmask(cache_io_data_M_wmask),
    .io_data_M_mem_size(cache_io_data_M_mem_size),
    .io_data_M_wdata(cache_io_data_M_wdata),
    .io_data_M_rdata(cache_io_data_M_rdata),
    .io_data_tlb_vpn2(cache_io_data_tlb_vpn2),
    .io_data_tlb_found(cache_io_data_tlb_found),
    .io_data_tlb_entry_pfn_0(cache_io_data_tlb_entry_pfn_0),
    .io_data_tlb_entry_pfn_1(cache_io_data_tlb_entry_pfn_1),
    .io_data_tlb_entry_c_0(cache_io_data_tlb_entry_c_0),
    .io_data_tlb_entry_c_1(cache_io_data_tlb_entry_c_1),
    .io_data_tlb_entry_d_0(cache_io_data_tlb_entry_d_0),
    .io_data_tlb_entry_d_1(cache_io_data_tlb_entry_d_1),
    .io_data_tlb_entry_v_0(cache_io_data_tlb_entry_v_0),
    .io_data_tlb_entry_v_1(cache_io_data_tlb_entry_v_1),
    .io_data_fence_tlb(cache_io_data_fence_tlb),
    .io_data_data_tlb_refill(cache_io_data_data_tlb_refill),
    .io_data_data_tlb_invalid(cache_io_data_data_tlb_invalid),
    .io_data_data_tlb_mod(cache_io_data_data_tlb_mod),
    .io_axi_ar_ready(cache_io_axi_ar_ready),
    .io_axi_ar_valid(cache_io_axi_ar_valid),
    .io_axi_ar_bits_id(cache_io_axi_ar_bits_id),
    .io_axi_ar_bits_addr(cache_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(cache_io_axi_ar_bits_len),
    .io_axi_ar_bits_size(cache_io_axi_ar_bits_size),
    .io_axi_r_ready(cache_io_axi_r_ready),
    .io_axi_r_valid(cache_io_axi_r_valid),
    .io_axi_r_bits_id(cache_io_axi_r_bits_id),
    .io_axi_r_bits_data(cache_io_axi_r_bits_data),
    .io_axi_r_bits_last(cache_io_axi_r_bits_last),
    .io_axi_aw_ready(cache_io_axi_aw_ready),
    .io_axi_aw_valid(cache_io_axi_aw_valid),
    .io_axi_aw_bits_addr(cache_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(cache_io_axi_aw_bits_len),
    .io_axi_aw_bits_size(cache_io_axi_aw_bits_size),
    .io_axi_w_ready(cache_io_axi_w_ready),
    .io_axi_w_valid(cache_io_axi_w_valid),
    .io_axi_w_bits_data(cache_io_axi_w_bits_data),
    .io_axi_w_bits_strb(cache_io_axi_w_bits_strb),
    .io_axi_w_bits_last(cache_io_axi_w_bits_last),
    .io_axi_b_valid(cache_io_axi_b_valid)
  );
  assign io_axi_ar_valid = cache_io_axi_ar_valid; // @[PuaMips.scala 22:10]
  assign io_axi_ar_bits_id = cache_io_axi_ar_bits_id; // @[PuaMips.scala 22:10]
  assign io_axi_ar_bits_addr = cache_io_axi_ar_bits_addr; // @[PuaMips.scala 22:10]
  assign io_axi_ar_bits_len = cache_io_axi_ar_bits_len; // @[PuaMips.scala 22:10]
  assign io_axi_ar_bits_size = cache_io_axi_ar_bits_size; // @[PuaMips.scala 22:10]
  assign io_axi_ar_bits_burst = 2'h1; // @[PuaMips.scala 22:10]
  assign io_axi_ar_bits_lock = 2'h0; // @[PuaMips.scala 22:10]
  assign io_axi_ar_bits_cache = 4'h0; // @[PuaMips.scala 22:10]
  assign io_axi_ar_bits_prot = 3'h0; // @[PuaMips.scala 22:10]
  assign io_axi_r_ready = cache_io_axi_r_ready; // @[PuaMips.scala 22:10]
  assign io_axi_aw_valid = cache_io_axi_aw_valid; // @[PuaMips.scala 22:10]
  assign io_axi_aw_bits_id = 4'h0; // @[PuaMips.scala 22:10]
  assign io_axi_aw_bits_addr = cache_io_axi_aw_bits_addr; // @[PuaMips.scala 22:10]
  assign io_axi_aw_bits_len = cache_io_axi_aw_bits_len; // @[PuaMips.scala 22:10]
  assign io_axi_aw_bits_size = cache_io_axi_aw_bits_size; // @[PuaMips.scala 22:10]
  assign io_axi_aw_bits_burst = 2'h1; // @[PuaMips.scala 22:10]
  assign io_axi_aw_bits_lock = 2'h0; // @[PuaMips.scala 22:10]
  assign io_axi_aw_bits_cache = 4'h0; // @[PuaMips.scala 22:10]
  assign io_axi_aw_bits_prot = 3'h0; // @[PuaMips.scala 22:10]
  assign io_axi_w_valid = cache_io_axi_w_valid; // @[PuaMips.scala 22:10]
  assign io_axi_w_bits_id = 4'h0; // @[PuaMips.scala 22:10]
  assign io_axi_w_bits_data = cache_io_axi_w_bits_data; // @[PuaMips.scala 22:10]
  assign io_axi_w_bits_strb = cache_io_axi_w_bits_strb; // @[PuaMips.scala 22:10]
  assign io_axi_w_bits_last = cache_io_axi_w_bits_last; // @[PuaMips.scala 22:10]
  assign io_axi_b_ready = 1'h1; // @[PuaMips.scala 22:10]
  assign io_debug_wb_pc = core_io_debug_wb_pc; // @[PuaMips.scala 21:12]
  assign io_debug_wb_rf_wen = core_io_debug_wb_rf_wen; // @[PuaMips.scala 21:12]
  assign io_debug_wb_rf_wnum = core_io_debug_wb_rf_wnum; // @[PuaMips.scala 21:12]
  assign io_debug_wb_rf_wdata = core_io_debug_wb_rf_wdata; // @[PuaMips.scala 21:12]
  assign io_debug_cp0_count = core_io_debug_cp0_count; // @[PuaMips.scala 21:12]
  assign io_debug_cp0_random = core_io_debug_cp0_random; // @[PuaMips.scala 21:12]
  assign io_debug_cp0_cause = core_io_debug_cp0_cause; // @[PuaMips.scala 21:12]
  assign io_debug_int = core_io_debug_int; // @[PuaMips.scala 21:12]
  assign io_debug_commit = core_io_debug_commit; // @[PuaMips.scala 21:12]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_ext_int = io_ext_int; // @[PuaMips.scala 20:14]
  assign core_io_inst_inst_0 = cache_io_inst_inst_0; // @[PuaMips.scala 17:16]
  assign core_io_inst_inst_1 = cache_io_inst_inst_1; // @[PuaMips.scala 17:16]
  assign core_io_inst_inst_valid_0 = cache_io_inst_inst_valid_0; // @[PuaMips.scala 17:16]
  assign core_io_inst_inst_valid_1 = cache_io_inst_inst_valid_1; // @[PuaMips.scala 17:16]
  assign core_io_inst_icache_stall = cache_io_inst_icache_stall; // @[PuaMips.scala 17:16]
  assign core_io_inst_tlb1_invalid = cache_io_inst_tlb1_invalid; // @[PuaMips.scala 17:16]
  assign core_io_inst_tlb2_vpn = cache_io_inst_tlb2_vpn; // @[PuaMips.scala 17:16]
  assign core_io_data_dstall = cache_io_data_dstall; // @[PuaMips.scala 18:16]
  assign core_io_data_M_rdata = cache_io_data_M_rdata; // @[PuaMips.scala 18:16]
  assign core_io_data_tlb_vpn2 = cache_io_data_tlb_vpn2; // @[PuaMips.scala 18:16]
  assign core_io_data_data_tlb_refill = cache_io_data_data_tlb_refill; // @[PuaMips.scala 18:16]
  assign core_io_data_data_tlb_invalid = cache_io_data_data_tlb_invalid; // @[PuaMips.scala 18:16]
  assign core_io_data_data_tlb_mod = cache_io_data_data_tlb_mod; // @[PuaMips.scala 18:16]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_inst_req = core_io_inst_req; // @[PuaMips.scala 17:16]
  assign cache_io_inst_addr_0 = core_io_inst_addr_0; // @[PuaMips.scala 17:16]
  assign cache_io_inst_addr_1 = core_io_inst_addr_1; // @[PuaMips.scala 17:16]
  assign cache_io_inst_cpu_stall = core_io_inst_cpu_stall; // @[PuaMips.scala 17:16]
  assign cache_io_inst_tlb2_found = core_io_inst_tlb2_found; // @[PuaMips.scala 17:16]
  assign cache_io_inst_tlb2_entry_pfn_0 = core_io_inst_tlb2_entry_pfn_0; // @[PuaMips.scala 17:16]
  assign cache_io_inst_tlb2_entry_pfn_1 = core_io_inst_tlb2_entry_pfn_1; // @[PuaMips.scala 17:16]
  assign cache_io_inst_tlb2_entry_c_0 = core_io_inst_tlb2_entry_c_0; // @[PuaMips.scala 17:16]
  assign cache_io_inst_tlb2_entry_c_1 = core_io_inst_tlb2_entry_c_1; // @[PuaMips.scala 17:16]
  assign cache_io_inst_tlb2_entry_v_0 = core_io_inst_tlb2_entry_v_0; // @[PuaMips.scala 17:16]
  assign cache_io_inst_tlb2_entry_v_1 = core_io_inst_tlb2_entry_v_1; // @[PuaMips.scala 17:16]
  assign cache_io_inst_fence_value = core_io_inst_fence_value; // @[PuaMips.scala 17:16]
  assign cache_io_inst_fence_addr = core_io_inst_fence_addr; // @[PuaMips.scala 17:16]
  assign cache_io_inst_fence_tlb = core_io_inst_fence_tlb; // @[PuaMips.scala 17:16]
  assign cache_io_data_stallM = core_io_data_stallM; // @[PuaMips.scala 18:16]
  assign cache_io_data_E_mem_va = core_io_data_E_mem_va; // @[PuaMips.scala 18:16]
  assign cache_io_data_M_mem_va = core_io_data_M_mem_va; // @[PuaMips.scala 18:16]
  assign cache_io_data_M_fence_addr = core_io_data_M_fence_addr; // @[PuaMips.scala 18:16]
  assign cache_io_data_M_fence_d = core_io_data_M_fence_d; // @[PuaMips.scala 18:16]
  assign cache_io_data_M_mem_en = core_io_data_M_mem_en; // @[PuaMips.scala 18:16]
  assign cache_io_data_M_mem_write = core_io_data_M_mem_write; // @[PuaMips.scala 18:16]
  assign cache_io_data_M_wmask = core_io_data_M_wmask; // @[PuaMips.scala 18:16]
  assign cache_io_data_M_mem_size = core_io_data_M_mem_size; // @[PuaMips.scala 18:16]
  assign cache_io_data_M_wdata = core_io_data_M_wdata; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_found = core_io_data_tlb_found; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_entry_pfn_0 = core_io_data_tlb_entry_pfn_0; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_entry_pfn_1 = core_io_data_tlb_entry_pfn_1; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_entry_c_0 = core_io_data_tlb_entry_c_0; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_entry_c_1 = core_io_data_tlb_entry_c_1; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_entry_d_0 = core_io_data_tlb_entry_d_0; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_entry_d_1 = core_io_data_tlb_entry_d_1; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_entry_v_0 = core_io_data_tlb_entry_v_0; // @[PuaMips.scala 18:16]
  assign cache_io_data_tlb_entry_v_1 = core_io_data_tlb_entry_v_1; // @[PuaMips.scala 18:16]
  assign cache_io_data_fence_tlb = core_io_data_fence_tlb; // @[PuaMips.scala 18:16]
  assign cache_io_axi_ar_ready = io_axi_ar_ready; // @[PuaMips.scala 22:10]
  assign cache_io_axi_r_valid = io_axi_r_valid; // @[PuaMips.scala 22:10]
  assign cache_io_axi_r_bits_id = io_axi_r_bits_id; // @[PuaMips.scala 22:10]
  assign cache_io_axi_r_bits_data = io_axi_r_bits_data; // @[PuaMips.scala 22:10]
  assign cache_io_axi_r_bits_last = io_axi_r_bits_last; // @[PuaMips.scala 22:10]
  assign cache_io_axi_aw_ready = io_axi_aw_ready; // @[PuaMips.scala 22:10]
  assign cache_io_axi_w_ready = io_axi_w_ready; // @[PuaMips.scala 22:10]
  assign cache_io_axi_b_valid = io_axi_b_valid; // @[PuaMips.scala 22:10]
endmodule
